

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701;

  XOR2_X1 U361 ( .A(G122), .B(G104), .Z(n474) );
  AND2_X1 U362 ( .A1(n496), .A2(n571), .ZN(n497) );
  INV_X1 U363 ( .A(G953), .ZN(n687) );
  AND2_X2 U364 ( .A1(n568), .A2(n589), .ZN(n563) );
  NAND2_X2 U365 ( .A1(n497), .A2(n593), .ZN(n512) );
  XNOR2_X2 U366 ( .A(n598), .B(KEYINPUT6), .ZN(n562) );
  NOR2_X1 U367 ( .A1(n622), .A2(G902), .ZN(n439) );
  INV_X1 U368 ( .A(n592), .ZN(n571) );
  NOR2_X1 U369 ( .A1(n625), .A2(n673), .ZN(n354) );
  NOR2_X1 U370 ( .A1(n653), .A2(n673), .ZN(n355) );
  XNOR2_X1 U371 ( .A(n428), .B(n427), .ZN(n592) );
  XNOR2_X1 U372 ( .A(n482), .B(n403), .ZN(n459) );
  INV_X4 U373 ( .A(G143), .ZN(n402) );
  XOR2_X1 U374 ( .A(G146), .B(G125), .Z(n461) );
  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n468) );
  OR2_X1 U376 ( .A1(n547), .A2(n546), .ZN(n372) );
  XNOR2_X1 U377 ( .A(n435), .B(KEYINPUT3), .ZN(n456) );
  XNOR2_X1 U378 ( .A(n495), .B(n494), .ZN(n526) );
  XNOR2_X1 U379 ( .A(n493), .B(G478), .ZN(n494) );
  XNOR2_X1 U380 ( .A(G116), .B(G137), .ZN(n429) );
  NAND2_X1 U381 ( .A1(n360), .A2(n359), .ZN(n358) );
  XNOR2_X1 U382 ( .A(n532), .B(KEYINPUT46), .ZN(n359) );
  AND2_X1 U383 ( .A1(n699), .A2(n525), .ZN(n360) );
  INV_X1 U384 ( .A(KEYINPUT48), .ZN(n357) );
  XOR2_X1 U385 ( .A(G137), .B(G140), .Z(n415) );
  NAND2_X1 U386 ( .A1(n687), .A2(G234), .ZN(n416) );
  XOR2_X1 U387 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n417) );
  XOR2_X1 U388 ( .A(n461), .B(KEYINPUT10), .Z(n472) );
  XOR2_X1 U389 ( .A(G902), .B(KEYINPUT15), .Z(n410) );
  OR2_X1 U390 ( .A1(G237), .A2(G902), .ZN(n464) );
  XNOR2_X1 U391 ( .A(n511), .B(n373), .ZN(n547) );
  INV_X1 U392 ( .A(KEYINPUT19), .ZN(n373) );
  XNOR2_X1 U393 ( .A(n409), .B(n343), .ZN(n517) );
  XNOR2_X1 U394 ( .A(n368), .B(G110), .ZN(n453) );
  INV_X1 U395 ( .A(KEYINPUT82), .ZN(n368) );
  XOR2_X1 U396 ( .A(G116), .B(G107), .Z(n488) );
  XNOR2_X1 U397 ( .A(n419), .B(n418), .ZN(n420) );
  INV_X1 U398 ( .A(KEYINPUT24), .ZN(n418) );
  XOR2_X1 U399 ( .A(G128), .B(KEYINPUT23), .Z(n419) );
  XNOR2_X1 U400 ( .A(G134), .B(G122), .ZN(n481) );
  XOR2_X1 U401 ( .A(G140), .B(G143), .Z(n467) );
  XNOR2_X1 U402 ( .A(G113), .B(G131), .ZN(n466) );
  XOR2_X1 U403 ( .A(KEYINPUT90), .B(KEYINPUT12), .Z(n470) );
  XNOR2_X1 U404 ( .A(n432), .B(n378), .ZN(n655) );
  XNOR2_X1 U405 ( .A(n405), .B(n379), .ZN(n378) );
  XNOR2_X1 U406 ( .A(n408), .B(n453), .ZN(n379) );
  XNOR2_X1 U407 ( .A(n404), .B(G107), .ZN(n405) );
  XNOR2_X1 U408 ( .A(n370), .B(n674), .ZN(n650) );
  XNOR2_X1 U409 ( .A(n463), .B(n352), .ZN(n370) );
  XNOR2_X1 U410 ( .A(n462), .B(n457), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n381), .B(n465), .ZN(n531) );
  XNOR2_X1 U412 ( .A(n363), .B(n362), .ZN(n361) );
  INV_X1 U413 ( .A(KEYINPUT106), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n517), .B(KEYINPUT1), .ZN(n590) );
  NOR2_X1 U415 ( .A1(n659), .A2(G902), .ZN(n480) );
  XNOR2_X1 U416 ( .A(n426), .B(n398), .ZN(n427) );
  XNOR2_X1 U417 ( .A(n353), .B(KEYINPUT22), .ZN(n573) );
  BUF_X1 U418 ( .A(n660), .Z(n669) );
  NOR2_X1 U419 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U420 ( .A(n407), .B(n406), .ZN(n408) );
  INV_X1 U421 ( .A(KEYINPUT4), .ZN(n403) );
  XNOR2_X1 U422 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U423 ( .A(n539), .B(n399), .ZN(n578) );
  NAND2_X1 U424 ( .A1(n365), .A2(n364), .ZN(n363) );
  INV_X1 U425 ( .A(n642), .ZN(n364) );
  INV_X1 U426 ( .A(KEYINPUT99), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n456), .B(n436), .ZN(n437) );
  NAND2_X1 U428 ( .A1(n383), .A2(n344), .ZN(n686) );
  XNOR2_X1 U429 ( .A(n358), .B(n357), .ZN(n383) );
  INV_X1 U430 ( .A(n648), .ZN(n382) );
  XNOR2_X1 U431 ( .A(n395), .B(n394), .ZN(n612) );
  XNOR2_X1 U432 ( .A(KEYINPUT105), .B(KEYINPUT41), .ZN(n394) );
  NOR2_X1 U433 ( .A1(n339), .A2(n582), .ZN(n395) );
  INV_X1 U434 ( .A(n372), .ZN(n549) );
  NAND2_X1 U435 ( .A1(n650), .A2(n620), .ZN(n391) );
  NOR2_X1 U436 ( .A1(n541), .A2(n448), .ZN(n502) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n447) );
  XNOR2_X1 U438 ( .A(KEYINPUT30), .B(KEYINPUT103), .ZN(n384) );
  NOR2_X1 U439 ( .A1(n547), .A2(n528), .ZN(n519) );
  INV_X1 U440 ( .A(KEYINPUT0), .ZN(n371) );
  BUF_X1 U441 ( .A(n598), .Z(n351) );
  XNOR2_X1 U442 ( .A(n369), .B(n456), .ZN(n674) );
  XNOR2_X1 U443 ( .A(n454), .B(n455), .ZN(n369) );
  XNOR2_X1 U444 ( .A(G119), .B(G110), .ZN(n422) );
  XNOR2_X1 U445 ( .A(n492), .B(n491), .ZN(n666) );
  XNOR2_X1 U446 ( .A(n397), .B(n396), .ZN(n659) );
  XNOR2_X1 U447 ( .A(n476), .B(n474), .ZN(n396) );
  XNOR2_X1 U448 ( .A(n475), .B(n473), .ZN(n397) );
  XNOR2_X1 U449 ( .A(n380), .B(KEYINPUT40), .ZN(n701) );
  NOR2_X1 U450 ( .A1(n531), .A2(n642), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n501), .B(KEYINPUT108), .ZN(n699) );
  XNOR2_X1 U452 ( .A(n374), .B(n347), .ZN(n697) );
  INV_X1 U453 ( .A(n567), .ZN(n375) );
  XNOR2_X1 U454 ( .A(n390), .B(n389), .ZN(n367) );
  INV_X1 U455 ( .A(KEYINPUT32), .ZN(n389) );
  NOR2_X1 U456 ( .A1(n573), .A2(n572), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n356), .B(n348), .ZN(n658) );
  NAND2_X1 U458 ( .A1(n669), .A2(G469), .ZN(n356) );
  OR2_X1 U459 ( .A1(n527), .A2(n526), .ZN(n339) );
  XNOR2_X1 U460 ( .A(n684), .B(G146), .ZN(n432) );
  AND2_X1 U461 ( .A1(G210), .A2(n464), .ZN(n340) );
  NOR2_X1 U462 ( .A1(n557), .A2(n339), .ZN(n341) );
  XOR2_X1 U463 ( .A(G131), .B(G134), .Z(n342) );
  NOR2_X1 U464 ( .A1(n655), .A2(G902), .ZN(n343) );
  AND2_X1 U465 ( .A1(n649), .A2(n382), .ZN(n344) );
  AND2_X1 U466 ( .A1(n561), .A2(n628), .ZN(n345) );
  XNOR2_X1 U467 ( .A(KEYINPUT97), .B(KEYINPUT33), .ZN(n346) );
  XOR2_X1 U468 ( .A(KEYINPUT77), .B(KEYINPUT35), .Z(n347) );
  XOR2_X1 U469 ( .A(n657), .B(n656), .Z(n348) );
  XOR2_X1 U470 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n349) );
  XOR2_X1 U471 ( .A(n499), .B(KEYINPUT36), .Z(n350) );
  XNOR2_X2 U472 ( .A(n564), .B(n346), .ZN(n613) );
  NAND2_X1 U473 ( .A1(n565), .A2(n341), .ZN(n353) );
  XNOR2_X1 U474 ( .A(n354), .B(n627), .ZN(G57) );
  XNOR2_X1 U475 ( .A(n355), .B(n654), .ZN(G51) );
  NAND2_X1 U476 ( .A1(n598), .A2(n579), .ZN(n385) );
  XNOR2_X2 U477 ( .A(n439), .B(n440), .ZN(n598) );
  INV_X1 U478 ( .A(n363), .ZN(n533) );
  NAND2_X1 U479 ( .A1(n361), .A2(n393), .ZN(n392) );
  XNOR2_X1 U480 ( .A(n498), .B(n366), .ZN(n365) );
  NAND2_X1 U481 ( .A1(n367), .A2(n635), .ZN(n576) );
  XNOR2_X1 U482 ( .A(n367), .B(G119), .ZN(G21) );
  XNOR2_X2 U483 ( .A(n372), .B(n371), .ZN(n565) );
  NOR2_X2 U484 ( .A1(n697), .A2(n576), .ZN(n388) );
  NAND2_X1 U485 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U486 ( .A(n566), .B(n377), .ZN(n376) );
  INV_X1 U487 ( .A(KEYINPUT34), .ZN(n377) );
  AND2_X2 U488 ( .A1(n590), .A2(n563), .ZN(n564) );
  XNOR2_X1 U489 ( .A(n386), .B(n349), .ZN(n679) );
  NAND2_X1 U490 ( .A1(n502), .A2(n578), .ZN(n381) );
  NAND2_X1 U491 ( .A1(n387), .A2(n345), .ZN(n386) );
  XNOR2_X1 U492 ( .A(n388), .B(KEYINPUT44), .ZN(n387) );
  INV_X1 U493 ( .A(n506), .ZN(n539) );
  NAND2_X1 U494 ( .A1(n506), .A2(n579), .ZN(n511) );
  XNOR2_X2 U495 ( .A(n391), .B(n340), .ZN(n506) );
  XNOR2_X2 U496 ( .A(n459), .B(n342), .ZN(n684) );
  XNOR2_X2 U497 ( .A(n402), .B(G128), .ZN(n482) );
  XNOR2_X1 U498 ( .A(n392), .B(n350), .ZN(n500) );
  INV_X1 U499 ( .A(n511), .ZN(n393) );
  NOR2_X2 U500 ( .A1(n663), .A2(n673), .ZN(n664) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n622) );
  XNOR2_X1 U502 ( .A(n459), .B(n458), .ZN(n463) );
  AND2_X1 U503 ( .A1(n621), .A2(n615), .ZN(n616) );
  XOR2_X1 U504 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n398) );
  XNOR2_X1 U505 ( .A(KEYINPUT72), .B(KEYINPUT38), .ZN(n399) );
  AND2_X1 U506 ( .A1(n613), .A2(n612), .ZN(n400) );
  XNOR2_X1 U507 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n401) );
  NOR2_X1 U508 ( .A1(n696), .A2(n701), .ZN(n532) );
  XNOR2_X1 U509 ( .A(n421), .B(n420), .ZN(n423) );
  INV_X1 U510 ( .A(KEYINPUT96), .ZN(n493) );
  NOR2_X1 U511 ( .A1(n614), .A2(n400), .ZN(n615) );
  XNOR2_X1 U512 ( .A(n490), .B(n489), .ZN(n491) );
  INV_X1 U513 ( .A(KEYINPUT63), .ZN(n626) );
  XNOR2_X1 U514 ( .A(n626), .B(KEYINPUT80), .ZN(n627) );
  NOR2_X1 U515 ( .A1(G952), .A2(n687), .ZN(n673) );
  XOR2_X1 U516 ( .A(KEYINPUT78), .B(KEYINPUT39), .Z(n465) );
  XNOR2_X1 U517 ( .A(KEYINPUT67), .B(G469), .ZN(n409) );
  XOR2_X1 U518 ( .A(n415), .B(G104), .Z(n404) );
  AND2_X1 U519 ( .A1(G227), .A2(n687), .ZN(n407) );
  XNOR2_X1 U520 ( .A(G101), .B(KEYINPUT74), .ZN(n406) );
  XOR2_X1 U521 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n412) );
  XNOR2_X1 U522 ( .A(KEYINPUT81), .B(n410), .ZN(n620) );
  NAND2_X1 U523 ( .A1(G234), .A2(n620), .ZN(n411) );
  XNOR2_X1 U524 ( .A(n412), .B(n411), .ZN(n425) );
  NAND2_X1 U525 ( .A1(n425), .A2(G221), .ZN(n414) );
  XOR2_X1 U526 ( .A(KEYINPUT86), .B(KEYINPUT21), .Z(n413) );
  XNOR2_X1 U527 ( .A(n414), .B(n413), .ZN(n593) );
  XNOR2_X1 U528 ( .A(n593), .B(KEYINPUT87), .ZN(n557) );
  XOR2_X1 U529 ( .A(n415), .B(n472), .Z(n685) );
  XNOR2_X1 U530 ( .A(n417), .B(n416), .ZN(n487) );
  NAND2_X1 U531 ( .A1(G221), .A2(n487), .ZN(n421) );
  XNOR2_X1 U532 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U533 ( .A(n685), .B(n424), .ZN(n668) );
  NOR2_X1 U534 ( .A1(G902), .A2(n668), .ZN(n428) );
  NAND2_X1 U535 ( .A1(n425), .A2(G217), .ZN(n426) );
  NOR2_X1 U536 ( .A1(n557), .A2(n571), .ZN(n589) );
  NAND2_X1 U537 ( .A1(n517), .A2(n589), .ZN(n541) );
  NAND2_X1 U538 ( .A1(G214), .A2(n464), .ZN(n579) );
  XNOR2_X1 U539 ( .A(G472), .B(KEYINPUT69), .ZN(n440) );
  XOR2_X1 U540 ( .A(KEYINPUT88), .B(KEYINPUT5), .Z(n430) );
  XNOR2_X1 U541 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U542 ( .A(n432), .B(n431), .ZN(n438) );
  XOR2_X1 U543 ( .A(KEYINPUT68), .B(G119), .Z(n434) );
  XNOR2_X1 U544 ( .A(G113), .B(G101), .ZN(n433) );
  XNOR2_X1 U545 ( .A(n434), .B(n433), .ZN(n435) );
  AND2_X1 U546 ( .A1(n468), .A2(G210), .ZN(n436) );
  NAND2_X1 U547 ( .A1(G234), .A2(G237), .ZN(n441) );
  XNOR2_X1 U548 ( .A(n441), .B(KEYINPUT14), .ZN(n444) );
  AND2_X1 U549 ( .A1(G953), .A2(n444), .ZN(n442) );
  NAND2_X1 U550 ( .A1(G902), .A2(n442), .ZN(n542) );
  XNOR2_X1 U551 ( .A(KEYINPUT98), .B(n542), .ZN(n443) );
  NOR2_X1 U552 ( .A1(G900), .A2(n443), .ZN(n445) );
  NAND2_X1 U553 ( .A1(G952), .A2(n444), .ZN(n609) );
  NOR2_X1 U554 ( .A1(G953), .A2(n609), .ZN(n544) );
  NOR2_X1 U555 ( .A1(n445), .A2(n544), .ZN(n446) );
  XNOR2_X1 U556 ( .A(n446), .B(KEYINPUT75), .ZN(n496) );
  NAND2_X1 U557 ( .A1(n447), .A2(n496), .ZN(n448) );
  INV_X1 U558 ( .A(n474), .ZN(n449) );
  NAND2_X1 U559 ( .A1(n449), .A2(KEYINPUT16), .ZN(n452) );
  INV_X1 U560 ( .A(KEYINPUT16), .ZN(n450) );
  NAND2_X1 U561 ( .A1(n450), .A2(n474), .ZN(n451) );
  NAND2_X1 U562 ( .A1(n452), .A2(n451), .ZN(n455) );
  XNOR2_X1 U563 ( .A(n488), .B(n453), .ZN(n454) );
  INV_X1 U564 ( .A(KEYINPUT18), .ZN(n457) );
  XNOR2_X1 U565 ( .A(KEYINPUT17), .B(KEYINPUT83), .ZN(n458) );
  AND2_X1 U566 ( .A1(G224), .A2(n687), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n467), .B(n466), .ZN(n476) );
  NAND2_X1 U568 ( .A1(G214), .A2(n468), .ZN(n469) );
  XNOR2_X1 U569 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U570 ( .A(n471), .B(KEYINPUT11), .Z(n475) );
  INV_X1 U571 ( .A(n472), .ZN(n473) );
  XOR2_X1 U572 ( .A(KEYINPUT13), .B(KEYINPUT91), .Z(n478) );
  XNOR2_X1 U573 ( .A(KEYINPUT92), .B(G475), .ZN(n477) );
  XNOR2_X1 U574 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U575 ( .A(n480), .B(n479), .Z(n503) );
  XNOR2_X1 U576 ( .A(n482), .B(n481), .ZN(n486) );
  XOR2_X1 U577 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n484) );
  XNOR2_X1 U578 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n483) );
  XNOR2_X1 U579 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U580 ( .A(n486), .B(n485), .Z(n492) );
  NAND2_X1 U581 ( .A1(G217), .A2(n487), .ZN(n490) );
  XNOR2_X1 U582 ( .A(n488), .B(KEYINPUT95), .ZN(n489) );
  NOR2_X1 U583 ( .A1(n666), .A2(G902), .ZN(n495) );
  NAND2_X1 U584 ( .A1(n503), .A2(n526), .ZN(n646) );
  NOR2_X1 U585 ( .A1(n531), .A2(n646), .ZN(n648) );
  OR2_X1 U586 ( .A1(n526), .A2(n503), .ZN(n642) );
  NOR2_X1 U587 ( .A1(n562), .A2(n512), .ZN(n498) );
  INV_X1 U588 ( .A(KEYINPUT107), .ZN(n499) );
  NAND2_X1 U589 ( .A1(n500), .A2(n590), .ZN(n501) );
  NAND2_X1 U590 ( .A1(n642), .A2(n646), .ZN(n555) );
  INV_X1 U591 ( .A(n555), .ZN(n583) );
  NAND2_X1 U592 ( .A1(KEYINPUT47), .A2(n583), .ZN(n507) );
  INV_X1 U593 ( .A(n502), .ZN(n504) );
  INV_X1 U594 ( .A(n503), .ZN(n527) );
  NAND2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n567) );
  NOR2_X1 U596 ( .A1(n504), .A2(n567), .ZN(n505) );
  NAND2_X1 U597 ( .A1(n506), .A2(n505), .ZN(n638) );
  NAND2_X1 U598 ( .A1(n507), .A2(n638), .ZN(n508) );
  XNOR2_X1 U599 ( .A(KEYINPUT76), .B(n508), .ZN(n523) );
  XNOR2_X1 U600 ( .A(KEYINPUT65), .B(KEYINPUT47), .ZN(n509) );
  NAND2_X1 U601 ( .A1(n509), .A2(n555), .ZN(n510) );
  XNOR2_X1 U602 ( .A(n510), .B(KEYINPUT71), .ZN(n518) );
  XOR2_X1 U603 ( .A(KEYINPUT104), .B(KEYINPUT28), .Z(n515) );
  INV_X1 U604 ( .A(n512), .ZN(n513) );
  NAND2_X1 U605 ( .A1(n513), .A2(n598), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U607 ( .A1(n517), .A2(n516), .ZN(n528) );
  NAND2_X1 U608 ( .A1(n518), .A2(n519), .ZN(n521) );
  INV_X1 U609 ( .A(n519), .ZN(n639) );
  NAND2_X1 U610 ( .A1(n639), .A2(KEYINPUT47), .ZN(n520) );
  NAND2_X1 U611 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U612 ( .A(n524), .B(KEYINPUT70), .ZN(n525) );
  NAND2_X1 U613 ( .A1(n579), .A2(n578), .ZN(n582) );
  INV_X1 U614 ( .A(n528), .ZN(n529) );
  NAND2_X1 U615 ( .A1(n612), .A2(n529), .ZN(n530) );
  XOR2_X1 U616 ( .A(KEYINPUT42), .B(n530), .Z(n696) );
  NAND2_X1 U617 ( .A1(n533), .A2(n579), .ZN(n534) );
  XOR2_X1 U618 ( .A(KEYINPUT100), .B(n534), .Z(n535) );
  INV_X1 U619 ( .A(n590), .ZN(n569) );
  NAND2_X1 U620 ( .A1(n535), .A2(n569), .ZN(n538) );
  XOR2_X1 U621 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n536) );
  XNOR2_X1 U622 ( .A(KEYINPUT43), .B(n536), .ZN(n537) );
  XNOR2_X1 U623 ( .A(n538), .B(n537), .ZN(n540) );
  NAND2_X1 U624 ( .A1(n540), .A2(n539), .ZN(n649) );
  NOR2_X1 U625 ( .A1(n351), .A2(n541), .ZN(n548) );
  NOR2_X1 U626 ( .A1(G898), .A2(n542), .ZN(n543) );
  NOR2_X1 U627 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U628 ( .A(n545), .B(KEYINPUT84), .ZN(n546) );
  NAND2_X1 U629 ( .A1(n548), .A2(n565), .ZN(n631) );
  INV_X1 U630 ( .A(KEYINPUT31), .ZN(n554) );
  XOR2_X1 U631 ( .A(KEYINPUT0), .B(n549), .Z(n551) );
  AND2_X1 U632 ( .A1(n590), .A2(n589), .ZN(n550) );
  NAND2_X1 U633 ( .A1(n351), .A2(n550), .ZN(n602) );
  NOR2_X1 U634 ( .A1(n551), .A2(n602), .ZN(n552) );
  XNOR2_X1 U635 ( .A(n552), .B(KEYINPUT89), .ZN(n553) );
  XNOR2_X1 U636 ( .A(n554), .B(n553), .ZN(n645) );
  NAND2_X1 U637 ( .A1(n631), .A2(n645), .ZN(n556) );
  NAND2_X1 U638 ( .A1(n556), .A2(n555), .ZN(n561) );
  INV_X1 U639 ( .A(n562), .ZN(n568) );
  NOR2_X1 U640 ( .A1(n568), .A2(n573), .ZN(n558) );
  NAND2_X1 U641 ( .A1(n569), .A2(n558), .ZN(n559) );
  XNOR2_X1 U642 ( .A(n559), .B(KEYINPUT79), .ZN(n560) );
  NAND2_X1 U643 ( .A1(n560), .A2(n592), .ZN(n628) );
  NAND2_X1 U644 ( .A1(n613), .A2(n565), .ZN(n566) );
  NOR2_X1 U645 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U646 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U647 ( .A1(n573), .A2(n592), .ZN(n575) );
  NOR2_X1 U648 ( .A1(n351), .A2(n590), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n635) );
  NOR2_X1 U650 ( .A1(n686), .A2(n679), .ZN(n577) );
  XNOR2_X1 U651 ( .A(n577), .B(KEYINPUT2), .ZN(n621) );
  INV_X1 U652 ( .A(n613), .ZN(n587) );
  NOR2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U654 ( .A(n580), .B(KEYINPUT114), .ZN(n581) );
  NOR2_X1 U655 ( .A1(n339), .A2(n581), .ZN(n585) );
  NOR2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U659 ( .A(n588), .B(KEYINPUT115), .ZN(n606) );
  OR2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U661 ( .A(KEYINPUT50), .B(n591), .ZN(n600) );
  NOR2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U663 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U665 ( .A(KEYINPUT112), .B(n596), .ZN(n597) );
  NOR2_X1 U666 ( .A1(n351), .A2(n597), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U669 ( .A(KEYINPUT51), .B(n603), .Z(n604) );
  NAND2_X1 U670 ( .A1(n604), .A2(n612), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n606), .A2(n605), .ZN(n608) );
  XOR2_X1 U672 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n607) );
  XNOR2_X1 U673 ( .A(n608), .B(n607), .ZN(n610) );
  NOR2_X1 U674 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U675 ( .A(KEYINPUT117), .B(n611), .Z(n614) );
  XNOR2_X1 U676 ( .A(KEYINPUT118), .B(n616), .ZN(n617) );
  NAND2_X1 U677 ( .A1(n617), .A2(n687), .ZN(n619) );
  XNOR2_X1 U678 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n618) );
  XNOR2_X1 U679 ( .A(n619), .B(n618), .ZN(G75) );
  NOR2_X2 U680 ( .A1(n621), .A2(n620), .ZN(n660) );
  NAND2_X1 U681 ( .A1(n660), .A2(G472), .ZN(n624) );
  XNOR2_X1 U682 ( .A(n622), .B(KEYINPUT62), .ZN(n623) );
  XNOR2_X1 U683 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U684 ( .A(G101), .B(n628), .ZN(G3) );
  NOR2_X1 U685 ( .A1(n642), .A2(n631), .ZN(n630) );
  XNOR2_X1 U686 ( .A(G104), .B(KEYINPUT109), .ZN(n629) );
  XNOR2_X1 U687 ( .A(n630), .B(n629), .ZN(G6) );
  NOR2_X1 U688 ( .A1(n646), .A2(n631), .ZN(n633) );
  XNOR2_X1 U689 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n632) );
  XNOR2_X1 U690 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U691 ( .A(G107), .B(n634), .ZN(G9) );
  XNOR2_X1 U692 ( .A(G110), .B(n635), .ZN(G12) );
  NOR2_X1 U693 ( .A1(n646), .A2(n639), .ZN(n637) );
  XNOR2_X1 U694 ( .A(G128), .B(KEYINPUT29), .ZN(n636) );
  XNOR2_X1 U695 ( .A(n637), .B(n636), .ZN(G30) );
  XNOR2_X1 U696 ( .A(G143), .B(n638), .ZN(G45) );
  NOR2_X1 U697 ( .A1(n642), .A2(n639), .ZN(n640) );
  XOR2_X1 U698 ( .A(KEYINPUT110), .B(n640), .Z(n641) );
  XNOR2_X1 U699 ( .A(G146), .B(n641), .ZN(G48) );
  NOR2_X1 U700 ( .A1(n642), .A2(n645), .ZN(n644) );
  XNOR2_X1 U701 ( .A(G113), .B(KEYINPUT111), .ZN(n643) );
  XNOR2_X1 U702 ( .A(n644), .B(n643), .ZN(G15) );
  NOR2_X1 U703 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U704 ( .A(G116), .B(n647), .Z(G18) );
  XOR2_X1 U705 ( .A(G134), .B(n648), .Z(G36) );
  XNOR2_X1 U706 ( .A(G140), .B(n649), .ZN(G42) );
  NAND2_X1 U707 ( .A1(n660), .A2(G210), .ZN(n652) );
  XNOR2_X1 U708 ( .A(n650), .B(n401), .ZN(n651) );
  XNOR2_X1 U709 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U710 ( .A(KEYINPUT56), .B(KEYINPUT120), .ZN(n654) );
  XOR2_X1 U711 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n657) );
  XNOR2_X1 U712 ( .A(n655), .B(KEYINPUT121), .ZN(n656) );
  NOR2_X1 U713 ( .A1(n673), .A2(n658), .ZN(G54) );
  XOR2_X1 U714 ( .A(n659), .B(KEYINPUT59), .Z(n662) );
  NAND2_X1 U715 ( .A1(n660), .A2(G475), .ZN(n661) );
  XNOR2_X1 U716 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U717 ( .A(n664), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U718 ( .A1(G478), .A2(n669), .ZN(n665) );
  XNOR2_X1 U719 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U720 ( .A1(n673), .A2(n667), .ZN(G63) );
  XNOR2_X1 U721 ( .A(n668), .B(KEYINPUT122), .ZN(n671) );
  NAND2_X1 U722 ( .A1(G217), .A2(n669), .ZN(n670) );
  XNOR2_X1 U723 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U724 ( .A1(n673), .A2(n672), .ZN(G66) );
  OR2_X1 U725 ( .A1(G898), .A2(n687), .ZN(n675) );
  NAND2_X1 U726 ( .A1(n675), .A2(n674), .ZN(n683) );
  NAND2_X1 U727 ( .A1(G953), .A2(G224), .ZN(n676) );
  XNOR2_X1 U728 ( .A(KEYINPUT61), .B(n676), .ZN(n677) );
  NAND2_X1 U729 ( .A1(n677), .A2(G898), .ZN(n678) );
  XNOR2_X1 U730 ( .A(n678), .B(KEYINPUT123), .ZN(n681) );
  NOR2_X1 U731 ( .A1(G953), .A2(n679), .ZN(n680) );
  NOR2_X1 U732 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U733 ( .A(n683), .B(n682), .ZN(G69) );
  XNOR2_X1 U734 ( .A(n685), .B(n684), .ZN(n689) );
  XNOR2_X1 U735 ( .A(n686), .B(n689), .ZN(n688) );
  NAND2_X1 U736 ( .A1(n688), .A2(n687), .ZN(n693) );
  XNOR2_X1 U737 ( .A(G227), .B(n689), .ZN(n690) );
  NAND2_X1 U738 ( .A1(n690), .A2(G900), .ZN(n691) );
  NAND2_X1 U739 ( .A1(n691), .A2(G953), .ZN(n692) );
  NAND2_X1 U740 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U741 ( .A(KEYINPUT124), .B(n694), .ZN(G72) );
  XOR2_X1 U742 ( .A(G137), .B(KEYINPUT126), .Z(n695) );
  XNOR2_X1 U743 ( .A(n696), .B(n695), .ZN(G39) );
  XNOR2_X1 U744 ( .A(n697), .B(G122), .ZN(n698) );
  XNOR2_X1 U745 ( .A(n698), .B(KEYINPUT125), .ZN(G24) );
  XOR2_X1 U746 ( .A(G125), .B(n699), .Z(n700) );
  XNOR2_X1 U747 ( .A(KEYINPUT37), .B(n700), .ZN(G27) );
  XOR2_X1 U748 ( .A(G131), .B(n701), .Z(G33) );
endmodule

