//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  NAND2_X1  g0009(.A1(new_n203), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n212), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(new_n217), .B2(new_n216), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT67), .B(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n202), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n214), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n220), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n253), .A3(G274), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n253), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n255), .B1(G238), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT13), .ZN(new_n259));
  INV_X1    g0059(.A(G226), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G232), .B2(new_n261), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G97), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n256), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n258), .A2(new_n259), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n259), .B1(new_n258), .B2(new_n272), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT14), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(G169), .ZN(new_n277));
  INV_X1    g0077(.A(G179), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n276), .B1(new_n275), .B2(G169), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n206), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n207), .A2(new_n264), .A3(KEYINPUT68), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G20), .B2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n242), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n207), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n289), .A2(new_n290), .B1(new_n207), .B2(G68), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n282), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT11), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G1), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n202), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT12), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n206), .A3(new_n281), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G68), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n299), .B1(new_n300), .B2(new_n302), .C1(new_n292), .C2(new_n293), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n279), .A2(new_n280), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n275), .A2(G200), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n303), .A2(new_n294), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n275), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n295), .B1(G41), .B2(G45), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n253), .A2(G232), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n254), .A2(new_n313), .A3(KEYINPUT75), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT75), .B1(new_n254), .B2(new_n313), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT70), .B1(new_n266), .B2(G33), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT70), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(new_n264), .A3(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n320), .A3(new_n267), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n260), .A2(G1698), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G223), .B2(G1698), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n317), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n256), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT76), .B1(new_n316), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G223), .A2(G1698), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n260), .B2(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n328), .A2(new_n318), .A3(new_n267), .A4(new_n320), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n253), .B1(new_n329), .B2(new_n317), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NOR4_X1   g0131(.A1(new_n330), .A2(new_n314), .A3(new_n315), .A4(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n311), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n254), .A2(new_n313), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n254), .A2(new_n313), .A3(KEYINPUT75), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n325), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(G179), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(G58), .B(G68), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n286), .A2(G159), .B1(new_n342), .B2(G20), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n321), .A2(new_n344), .A3(new_n207), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G68), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n321), .B2(new_n207), .ZN(new_n347));
  OAI211_X1 g0147(.A(KEYINPUT16), .B(new_n343), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n348), .A2(new_n282), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT3), .B(G33), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(G20), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n268), .A2(new_n207), .A3(new_n352), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n202), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n343), .B1(new_n358), .B2(KEYINPUT72), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  AOI211_X1 g0160(.A(new_n360), .B(new_n202), .C1(new_n356), .C2(new_n357), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n350), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT8), .B(G58), .Z(new_n363));
  INV_X1    g0163(.A(new_n282), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(new_n296), .A4(new_n301), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT8), .B(G58), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n297), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT73), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n301), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n367), .B(new_n370), .C1(new_n373), .C2(new_n300), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n370), .B1(new_n365), .B2(new_n367), .ZN(new_n377));
  INV_X1    g0177(.A(new_n374), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n349), .A2(new_n362), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT18), .B1(new_n341), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n336), .A2(new_n337), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n331), .B1(new_n382), .B2(new_n330), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n316), .A2(KEYINPUT76), .A3(new_n325), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n339), .B1(new_n385), .B2(new_n311), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n375), .A2(new_n379), .ZN(new_n387));
  INV_X1    g0187(.A(new_n343), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n268), .A2(new_n207), .B1(new_n353), .B2(new_n352), .ZN(new_n389));
  AOI211_X1 g0189(.A(G20), .B(new_n351), .C1(new_n265), .C2(new_n267), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(new_n360), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n358), .A2(KEYINPUT72), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT16), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n348), .A2(new_n282), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n386), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n381), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n338), .A2(G190), .ZN(new_n401));
  INV_X1    g0201(.A(G200), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n385), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n400), .B1(new_n403), .B2(new_n396), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n402), .B1(new_n326), .B2(new_n332), .ZN(new_n405));
  INV_X1    g0205(.A(new_n401), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n380), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n399), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G222), .A2(G1698), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n261), .A2(G223), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n355), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(new_n256), .C1(G77), .C2(new_n355), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n257), .A2(G226), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n254), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n307), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(G200), .B2(new_n416), .ZN(new_n418));
  INV_X1    g0218(.A(new_n300), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n242), .B1(new_n295), .B2(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G50), .B2(new_n296), .ZN(new_n422));
  OAI21_X1  g0222(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n423));
  INV_X1    g0223(.A(G150), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n423), .B1(new_n366), .B2(new_n289), .C1(new_n287), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n282), .B2(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n426), .A2(KEYINPUT9), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(KEYINPUT9), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n418), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT10), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n416), .A2(G179), .ZN(new_n431));
  AOI211_X1 g0231(.A(new_n426), .B(new_n431), .C1(new_n311), .C2(new_n416), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n419), .A2(G77), .A3(new_n301), .ZN(new_n435));
  XOR2_X1   g0235(.A(new_n435), .B(KEYINPUT69), .Z(new_n436));
  NAND2_X1  g0236(.A1(G20), .A2(G77), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT15), .B(G87), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n437), .B1(new_n289), .B2(new_n438), .C1(new_n287), .C2(new_n366), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(new_n282), .B1(new_n290), .B2(new_n297), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G244), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n256), .A2(new_n251), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n355), .A2(G232), .A3(new_n261), .ZN(new_n444));
  INV_X1    g0244(.A(G107), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n355), .A2(G1698), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n444), .B1(new_n445), .B2(new_n355), .C1(new_n446), .C2(new_n221), .ZN(new_n447));
  AOI211_X1 g0247(.A(new_n255), .B(new_n443), .C1(new_n447), .C2(new_n256), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n441), .B1(new_n448), .B2(G169), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n278), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n441), .B1(G190), .B2(new_n448), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n402), .B2(new_n448), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n310), .A2(new_n410), .A3(new_n434), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n318), .A2(new_n320), .A3(new_n207), .A4(new_n267), .ZN(new_n459));
  INV_X1    g0259(.A(G87), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT22), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n355), .A2(new_n462), .A3(new_n207), .A4(G87), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n445), .A2(KEYINPUT23), .A3(G20), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT23), .B1(new_n445), .B2(G20), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(KEYINPUT87), .B(new_n458), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n461), .B2(new_n463), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT24), .B1(new_n470), .B2(new_n471), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n469), .B(new_n282), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n295), .A2(G33), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT78), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n300), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT25), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n296), .B2(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n445), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n478), .A2(G107), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n318), .A2(new_n320), .A3(new_n267), .ZN(new_n484));
  INV_X1    g0284(.A(G257), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n261), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(KEYINPUT88), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT88), .ZN(new_n488));
  INV_X1    g0288(.A(new_n486), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n321), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n261), .A2(G250), .ZN(new_n492));
  INV_X1    g0292(.A(G294), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n321), .A2(new_n492), .B1(new_n264), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n256), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n295), .B(G45), .C1(new_n249), .C2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT80), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n498), .A2(new_n499), .B1(KEYINPUT5), .B2(new_n249), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n250), .A2(G1), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(KEYINPUT80), .C1(KEYINPUT5), .C2(new_n249), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(G274), .A3(new_n253), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n256), .B1(new_n500), .B2(new_n502), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G264), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n497), .A2(new_n278), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n494), .B1(new_n487), .B2(new_n490), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n503), .B(new_n505), .C1(new_n507), .C2(new_n253), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n311), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n483), .A2(KEYINPUT89), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT89), .ZN(new_n511));
  INV_X1    g0311(.A(new_n482), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT87), .B1(new_n464), .B2(new_n468), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(KEYINPUT24), .A3(new_n472), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n470), .A2(new_n471), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n364), .B1(new_n515), .B2(new_n458), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n506), .A2(new_n509), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n511), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(G97), .B1(new_n477), .B2(new_n300), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n296), .A2(new_n270), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT79), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT79), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g0328(.A(G97), .B(G107), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n530));
  NOR2_X1   g0330(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(KEYINPUT6), .B2(new_n270), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n533), .A2(new_n207), .B1(new_n290), .B2(new_n287), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n445), .B1(new_n356), .B2(new_n357), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n282), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n504), .A2(G257), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n503), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n442), .A2(G1698), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT4), .B1(new_n484), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n355), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n355), .A2(G250), .A3(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G283), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n256), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n278), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n503), .A3(new_n538), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n311), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n537), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(G200), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n547), .A2(G190), .A3(new_n503), .A4(new_n538), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(new_n528), .A3(new_n536), .A4(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n289), .A2(KEYINPUT19), .A3(new_n270), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n460), .A2(new_n270), .A3(new_n445), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n271), .B2(G20), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n557), .B2(KEYINPUT19), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n459), .A2(new_n202), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n282), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n438), .A2(new_n297), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n477), .A2(new_n300), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(new_n561), .C1(new_n438), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n442), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(G238), .B2(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(G116), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n321), .A2(new_n565), .B1(new_n264), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n256), .ZN(new_n568));
  INV_X1    g0368(.A(G274), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n501), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n570), .B(new_n253), .C1(G250), .C2(new_n501), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n278), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n311), .B1(new_n568), .B2(new_n571), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n563), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT81), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n562), .B2(new_n460), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n478), .A2(KEYINPUT81), .A3(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n560), .A2(new_n561), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n572), .A2(G200), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n568), .A2(G190), .A3(new_n571), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n551), .A2(new_n554), .A3(new_n575), .A4(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n496), .A2(new_n256), .B1(G264), .B2(new_n504), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n585), .A2(G190), .A3(new_n503), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n508), .A2(G200), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n475), .A2(new_n586), .A3(new_n482), .A4(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n504), .A2(G270), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT82), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n504), .A2(KEYINPUT82), .A3(G270), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n485), .A2(new_n261), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(G264), .B2(new_n261), .ZN(new_n595));
  INV_X1    g0395(.A(G303), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n321), .A2(new_n595), .B1(new_n596), .B2(new_n355), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n256), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n592), .A2(new_n503), .A3(new_n593), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G200), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n545), .B(new_n207), .C1(G33), .C2(new_n270), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n566), .A2(G20), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n282), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT20), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT83), .B1(new_n603), .B2(new_n604), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n296), .A2(new_n566), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n478), .B2(new_n566), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n606), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n600), .A2(KEYINPUT85), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n307), .B2(new_n599), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT85), .B1(new_n600), .B2(new_n612), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n593), .A2(new_n503), .A3(new_n598), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT82), .B1(new_n504), .B2(G270), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n311), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT84), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT21), .A4(new_n611), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n599), .A2(G169), .A3(new_n611), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT21), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT84), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n619), .A2(G179), .A3(new_n611), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n622), .A2(new_n625), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n616), .A2(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n457), .A2(new_n521), .A3(new_n589), .A4(new_n629), .ZN(G372));
  NOR2_X1   g0430(.A1(new_n517), .A2(new_n518), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n589), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n575), .ZN(new_n633));
  INV_X1    g0433(.A(new_n551), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(KEYINPUT26), .A3(new_n575), .A4(new_n583), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n583), .A2(new_n575), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n551), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n633), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n457), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n386), .A2(new_n397), .A3(new_n396), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n397), .B1(new_n386), .B2(new_n396), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n381), .A2(KEYINPUT90), .A3(new_n398), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n308), .A2(new_n451), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n304), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n649), .B2(new_n409), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n432), .B1(new_n650), .B2(new_n430), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n641), .A2(new_n651), .ZN(G369));
  NAND3_X1  g0452(.A1(new_n295), .A2(new_n207), .A3(G13), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT91), .Z(new_n655));
  INV_X1    g0455(.A(G213), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n653), .B2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n628), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n588), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n521), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n631), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n661), .A2(new_n612), .ZN(new_n668));
  MUX2_X1   g0468(.A(new_n629), .B(new_n628), .S(new_n668), .Z(new_n669));
  XNOR2_X1  g0469(.A(KEYINPUT92), .B(G330), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n631), .A2(new_n660), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n521), .A2(new_n664), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n517), .A2(new_n661), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n667), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0478(.A(new_n215), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  NOR4_X1   g0480(.A1(new_n680), .A2(new_n295), .A3(G116), .A4(new_n556), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n211), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT28), .Z(new_n683));
  NAND2_X1  g0483(.A1(new_n640), .A2(new_n661), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n589), .B1(new_n520), .B2(new_n628), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT96), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n638), .A2(KEYINPUT95), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT95), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n690), .B(new_n636), .C1(new_n551), .C2(new_n637), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n633), .B1(new_n692), .B2(new_n635), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n589), .B(KEYINPUT96), .C1(new_n520), .C2(new_n628), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n688), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n661), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n685), .B1(new_n696), .B2(KEYINPUT29), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n629), .A2(new_n521), .A3(new_n589), .A4(new_n661), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n585), .A2(new_n547), .A3(new_n540), .A4(new_n573), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n599), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n549), .A2(new_n278), .A3(new_n572), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(KEYINPUT30), .A3(new_n585), .A4(new_n619), .ZN(new_n703));
  AOI21_X1  g0503(.A(G179), .B1(new_n568), .B2(new_n571), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n599), .A2(new_n704), .A3(new_n508), .A4(new_n549), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT31), .B1(new_n706), .B2(new_n660), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT94), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n660), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT94), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n698), .A2(new_n709), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n670), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n697), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n683), .B1(new_n718), .B2(G1), .ZN(G364));
  OAI21_X1  g0519(.A(G20), .B1(KEYINPUT97), .B2(G169), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(KEYINPUT97), .A2(G169), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n206), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n215), .A2(new_n321), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n247), .A2(new_n250), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n728), .B(new_n729), .C1(new_n250), .C2(new_n211), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n215), .A2(new_n355), .ZN(new_n731));
  INV_X1    g0531(.A(G355), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(G116), .B2(new_n215), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n727), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n207), .A2(G13), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n295), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n680), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n207), .A2(new_n278), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G190), .A3(new_n402), .ZN(new_n741));
  INV_X1    g0541(.A(G322), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n207), .A2(G179), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G190), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n355), .B(new_n743), .C1(G329), .C2(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n740), .A2(KEYINPUT98), .A3(new_n745), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT98), .B1(new_n740), .B2(new_n745), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G311), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n744), .A2(new_n307), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n744), .A2(G190), .A3(G200), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n596), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n740), .A2(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n307), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(G326), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n307), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n207), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n758), .A2(G190), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G294), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n748), .A2(new_n753), .A3(new_n760), .A4(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n746), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT32), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(new_n445), .B2(new_n754), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  INV_X1    g0572(.A(new_n759), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(new_n242), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n751), .A2(new_n290), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n355), .B1(new_n756), .B2(new_n460), .C1(new_n201), .C2(new_n741), .ZN(new_n776));
  OR4_X1    g0576(.A1(new_n771), .A2(new_n774), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G97), .A2(new_n763), .B1(new_n764), .B2(G68), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT99), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n767), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT100), .ZN(new_n781));
  INV_X1    g0581(.A(new_n723), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n780), .B2(KEYINPUT100), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n739), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n726), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n669), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n738), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n671), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n669), .A2(new_n670), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(G396));
  AOI22_X1  g0590(.A1(G137), .A2(new_n759), .B1(new_n764), .B2(G150), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT103), .Z(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT104), .B(G143), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n792), .B1(new_n768), .B2(new_n751), .C1(new_n741), .C2(new_n793), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT34), .Z(new_n795));
  INV_X1    g0595(.A(new_n754), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n763), .A2(G58), .B1(new_n796), .B2(G68), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n321), .B1(new_n747), .B2(G132), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n797), .B(new_n798), .C1(new_n242), .C2(new_n756), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n762), .A2(new_n270), .B1(new_n741), .B2(new_n493), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT102), .Z(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n268), .B1(new_n746), .B2(new_n802), .C1(new_n773), .C2(new_n596), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n752), .B2(G116), .ZN(new_n804));
  INV_X1    g0604(.A(new_n756), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n764), .A2(G283), .B1(new_n805), .B2(G107), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n804), .B(new_n806), .C1(new_n460), .C2(new_n754), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n795), .A2(new_n799), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n723), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n782), .A2(new_n725), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT101), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n787), .B1(new_n290), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n441), .A2(new_n660), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n454), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n452), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n451), .A2(new_n661), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n809), .B(new_n813), .C1(new_n819), .C2(new_n725), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n819), .A2(new_n640), .A3(new_n661), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(KEYINPUT105), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n684), .A2(new_n818), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n717), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n787), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n824), .A2(new_n717), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n820), .B1(new_n826), .B2(new_n827), .ZN(G384));
  INV_X1    g0628(.A(KEYINPUT35), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n209), .B(G116), .C1(new_n533), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n829), .B2(new_n533), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT36), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n211), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n295), .B(G13), .C1(new_n833), .C2(new_n243), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n707), .A2(new_n708), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n698), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n306), .A2(new_n661), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n309), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n304), .B(new_n308), .C1(new_n306), .C2(new_n661), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n818), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(KEYINPUT108), .A2(KEYINPUT40), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n837), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n407), .A2(new_n380), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n845), .A2(new_n350), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n374), .B(new_n369), .C1(new_n846), .C2(new_n395), .ZN(new_n847));
  INV_X1    g0647(.A(new_n658), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n386), .A2(new_n847), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT37), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n396), .A2(new_n848), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n844), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n341), .A2(new_n380), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n852), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n848), .B(new_n847), .C1(new_n399), .C2(new_n409), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT40), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n843), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n837), .A2(new_n841), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT108), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n404), .A2(new_n408), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n645), .A2(new_n871), .A3(new_n646), .ZN(new_n872));
  INV_X1    g0672(.A(new_n853), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n844), .A2(KEYINPUT90), .A3(new_n853), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n855), .B2(new_n854), .ZN(new_n877));
  INV_X1    g0677(.A(new_n854), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(new_n642), .A3(KEYINPUT37), .A4(new_n856), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT106), .B(new_n862), .C1(new_n874), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n864), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n878), .A2(new_n856), .B1(new_n875), .B2(KEYINPUT37), .ZN(new_n883));
  NOR4_X1   g0683(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT90), .A4(new_n857), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n872), .A2(new_n873), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n870), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n868), .B1(KEYINPUT40), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT109), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n456), .B1(new_n698), .B2(new_n836), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n893), .A2(new_n670), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT107), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n882), .B2(new_n888), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n304), .A2(new_n660), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n865), .A2(new_n897), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n898), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n647), .A2(new_n848), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n839), .A2(new_n840), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n821), .B2(new_n817), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n904), .B1(new_n907), .B2(new_n865), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n896), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n903), .A2(new_n896), .A3(new_n908), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n651), .B1(new_n697), .B2(new_n456), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n912), .B(new_n913), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n895), .A2(new_n914), .B1(new_n295), .B2(new_n735), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n895), .A2(new_n914), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n835), .B1(new_n915), .B2(new_n916), .ZN(G367));
  INV_X1    g0717(.A(new_n718), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n676), .A2(new_n663), .ZN(new_n919));
  INV_X1    g0719(.A(new_n665), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n672), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n671), .B(new_n665), .C1(new_n676), .C2(new_n663), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n718), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT113), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n634), .A2(new_n660), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n537), .A2(new_n660), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n551), .A2(new_n554), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n665), .B2(new_n666), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT44), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n665), .A2(new_n666), .A3(new_n929), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT45), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n672), .A2(new_n676), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n931), .B2(new_n934), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT113), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n718), .A2(new_n923), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n925), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT114), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n925), .A2(new_n938), .A3(KEYINPUT114), .A4(new_n940), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n918), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n680), .B(KEYINPUT41), .Z(new_n946));
  OAI21_X1  g0746(.A(new_n736), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n920), .A2(new_n929), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT42), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n551), .B1(new_n521), .B2(new_n928), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n661), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n661), .B1(new_n580), .B2(new_n579), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n633), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT110), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n952), .A2(new_n637), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT111), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n961));
  NAND3_X1  g0761(.A1(new_n951), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  MUX2_X1   g0762(.A(new_n961), .B(KEYINPUT43), .S(new_n959), .Z(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n951), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n672), .A2(new_n676), .A3(new_n929), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n947), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n960), .A2(new_n726), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n728), .A2(new_n237), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n727), .B1(new_n215), .B2(new_n438), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n738), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n773), .A2(new_n802), .B1(new_n445), .B2(new_n762), .ZN(new_n972));
  INV_X1    g0772(.A(new_n764), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n973), .A2(new_n493), .B1(new_n270), .B2(new_n754), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n752), .A2(G283), .ZN(new_n976));
  INV_X1    g0776(.A(G317), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n741), .A2(new_n596), .B1(new_n746), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n484), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT115), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n805), .B(G116), .C1(new_n981), .C2(KEYINPUT46), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT46), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n763), .A2(G68), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n201), .B2(new_n756), .C1(new_n773), .C2(new_n793), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n355), .B1(new_n741), .B2(new_n424), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G137), .B2(new_n747), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n764), .A2(G159), .B1(new_n796), .B2(G77), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(new_n242), .C2(new_n751), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n980), .A2(new_n984), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT47), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n971), .B1(new_n992), .B2(new_n723), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n968), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n967), .A2(new_n994), .ZN(G387));
  NAND2_X1  g0795(.A1(new_n925), .A2(new_n940), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n996), .B(new_n680), .C1(new_n718), .C2(new_n923), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n676), .A2(new_n785), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n234), .A2(new_n250), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n556), .A2(G116), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n999), .A2(new_n728), .B1(new_n1000), .B2(new_n731), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n366), .B2(G50), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n363), .A2(new_n1002), .A3(new_n242), .ZN(new_n1005));
  AOI21_X1  g0805(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n1000), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1001), .A2(new_n1007), .B1(new_n445), .B2(new_n679), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n727), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n738), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n973), .A2(new_n366), .B1(new_n290), .B2(new_n756), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G159), .B2(new_n759), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n752), .A2(G68), .ZN(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT117), .B(G150), .Z(new_n1014));
  OAI22_X1  g0814(.A1(new_n741), .A2(new_n242), .B1(new_n1014), .B2(new_n746), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(new_n321), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n438), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n763), .A2(new_n1017), .B1(new_n796), .B2(G97), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1012), .A2(new_n1013), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n751), .A2(new_n596), .B1(new_n977), .B2(new_n741), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT118), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(KEYINPUT118), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G311), .A2(new_n764), .B1(new_n759), .B2(G322), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n762), .A2(new_n755), .B1(new_n756), .B2(new_n493), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n484), .B1(G326), .B2(new_n747), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n566), .C2(new_n754), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT49), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1019), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1010), .B1(new_n1033), .B2(new_n723), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n923), .A2(new_n737), .B1(new_n998), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n997), .A2(new_n1035), .ZN(G393));
  NOR2_X1   g0836(.A1(new_n728), .A2(new_n241), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n727), .B1(new_n215), .B2(new_n270), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n738), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n741), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G317), .A2(new_n759), .B1(new_n1040), .B2(G311), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT119), .B(KEYINPUT52), .Z(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n973), .A2(new_n596), .B1(new_n566), .B2(new_n762), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G283), .B2(new_n805), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n268), .B1(new_n746), .B2(new_n742), .C1(new_n445), .C2(new_n754), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n752), .B2(G294), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n762), .A2(new_n290), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n973), .A2(new_n242), .B1(new_n756), .B2(new_n202), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G87), .C2(new_n796), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n793), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n321), .B1(new_n747), .B2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n366), .C2(new_n751), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G150), .A2(new_n759), .B1(new_n1040), .B2(G159), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT51), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1048), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1039), .B1(new_n1057), .B2(new_n723), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n929), .B2(new_n785), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n938), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n736), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n943), .A2(new_n944), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n680), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n996), .B2(new_n1060), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(G390));
  NAND3_X1  g0866(.A1(new_n837), .A2(new_n841), .A3(G330), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n907), .A2(new_n900), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n898), .B2(new_n902), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n899), .B1(new_n882), .B2(new_n888), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n695), .A2(new_n661), .A3(new_n816), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n906), .B1(new_n1072), .B2(new_n817), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1068), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n864), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n887), .B2(KEYINPUT106), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n862), .B1(new_n874), .B2(new_n880), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT106), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1072), .A2(new_n817), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1081), .B(new_n899), .C1(new_n1082), .C2(new_n906), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n716), .A2(new_n905), .A3(new_n670), .A4(new_n819), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n901), .B1(new_n1081), .B2(new_n897), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1084), .C1(new_n1085), .C2(new_n1069), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n837), .A2(G330), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n457), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n651), .C1(new_n697), .C2(new_n456), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n821), .A2(new_n817), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n716), .A2(new_n670), .A3(new_n819), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1092), .A2(new_n906), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1093), .B2(new_n1068), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n906), .B1(new_n1087), .B2(new_n818), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1082), .A2(new_n1084), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1075), .A2(new_n1086), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1097), .B(KEYINPUT120), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1075), .A2(new_n1086), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n680), .B(new_n1098), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n737), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n738), .B1(new_n811), .B2(new_n363), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1049), .B1(G283), .B2(new_n759), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n445), .B2(new_n973), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n751), .A2(new_n270), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n268), .B1(new_n746), .B2(new_n493), .C1(new_n741), .C2(new_n566), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n754), .A2(new_n202), .B1(new_n756), .B2(new_n460), .ZN(new_n1109));
  OR4_X1    g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1014), .A2(new_n756), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT53), .Z(new_n1112));
  AND2_X1   g0912(.A1(new_n747), .A2(G125), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n268), .B(new_n1113), .C1(G132), .C2(new_n1040), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G159), .A2(new_n763), .B1(new_n759), .B2(G128), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n764), .A2(G137), .B1(new_n796), .B2(G50), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  NAND2_X1  g0917(.A1(new_n752), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1110), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1104), .B1(new_n1120), .B2(new_n723), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n1085), .B2(new_n725), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1102), .A2(new_n1103), .A3(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(G330), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n426), .A2(new_n658), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n434), .B(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1126), .B(new_n1127), .Z(new_n1128));
  NOR3_X1   g0928(.A1(new_n890), .A2(new_n1124), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1128), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1077), .A2(new_n1080), .B1(KEYINPUT108), .B2(new_n869), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n865), .A2(KEYINPUT40), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1131), .A2(new_n867), .B1(new_n1132), .B2(new_n843), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1133), .B2(G330), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n903), .A2(new_n896), .A3(new_n908), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1129), .A2(new_n1134), .B1(new_n1135), .B2(new_n909), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1128), .B1(new_n890), .B2(new_n1124), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(G330), .A3(new_n1130), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n910), .A2(new_n1137), .A3(new_n911), .A4(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT124), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1090), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1098), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(KEYINPUT57), .A4(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1143), .A2(new_n1136), .A3(new_n1139), .A4(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT124), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1144), .A2(KEYINPUT125), .A3(new_n1146), .A4(new_n680), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT57), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  AND4_X1   g0951(.A1(KEYINPUT57), .A2(new_n1143), .A3(new_n1139), .A4(new_n1136), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1063), .B1(new_n1152), .B2(new_n1141), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT125), .B1(new_n1153), .B2(new_n1146), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n787), .B1(new_n242), .B2(new_n812), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n321), .A2(new_n249), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n985), .B1(new_n755), .B2(new_n746), .C1(new_n445), .C2(new_n741), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n1017), .C2(new_n752), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n754), .A2(new_n201), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G77), .B2(new_n805), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G97), .A2(new_n764), .B1(new_n759), .B2(G116), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT58), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1157), .B(new_n242), .C1(G33), .C2(G41), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n752), .A2(G137), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n763), .A2(G150), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G125), .A2(new_n759), .B1(new_n764), .B2(G132), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G128), .A2(new_n1040), .B1(new_n805), .B2(new_n1117), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n768), .B2(new_n754), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT121), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1164), .B(new_n1165), .C1(new_n1171), .C2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(KEYINPUT122), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT122), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n723), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1156), .B1(new_n1178), .B2(new_n1180), .C1(new_n1130), .C2(new_n725), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT123), .Z(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1140), .B2(new_n737), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1155), .A2(new_n1183), .ZN(G375));
  AOI21_X1  g0984(.A(new_n736), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n906), .A2(new_n724), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n738), .B1(new_n811), .B2(G68), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n973), .A2(new_n566), .B1(new_n756), .B2(new_n270), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G294), .B2(new_n759), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n752), .A2(G107), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n268), .B1(new_n746), .B2(new_n596), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G283), .B2(new_n1040), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n763), .A2(new_n1017), .B1(new_n796), .B2(G77), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n752), .A2(G150), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1040), .A2(G137), .B1(new_n747), .B2(G128), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1160), .B1(G132), .B2(new_n759), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1195), .A2(new_n484), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n764), .A2(new_n1117), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n242), .B2(new_n762), .C1(new_n768), .C2(new_n756), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1194), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1187), .B1(new_n1201), .B2(new_n723), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1185), .B1(new_n1186), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1094), .A2(new_n1090), .A3(new_n1096), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n946), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1203), .B1(new_n1099), .B2(new_n1206), .ZN(G381));
  OR4_X1    g1007(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(G387), .A2(new_n1208), .A3(G390), .A4(G378), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(new_n1155), .A3(new_n1183), .ZN(G407));
  INV_X1    g1010(.A(G378), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n656), .A2(G343), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(G407), .B(G213), .C1(G375), .C2(new_n1213), .ZN(G409));
  OAI211_X1 g1014(.A(G378), .B(new_n1183), .C1(new_n1151), .C2(new_n1154), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1148), .A2(new_n946), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1140), .A2(new_n737), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1181), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1211), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1212), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT60), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1097), .A2(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(new_n1204), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1204), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n680), .A3(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1226), .A2(G384), .A3(new_n1203), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G384), .B1(new_n1226), .B2(new_n1203), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1220), .A2(new_n1221), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT62), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1212), .A2(G2897), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT126), .Z(new_n1234));
  XNOR2_X1  g1034(.A(new_n1229), .B(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT61), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1212), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT62), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n1229), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1231), .A2(new_n1236), .A3(new_n1237), .A4(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G390), .B1(new_n967), .B2(new_n994), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  XOR2_X1   g1043(.A(G393), .B(G396), .Z(new_n1244));
  NAND3_X1  g1044(.A1(new_n967), .A2(new_n994), .A3(G390), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1244), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n967), .A2(new_n994), .A3(G390), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1248), .B2(new_n1242), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1241), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1235), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1250), .B(new_n1237), .C1(new_n1238), .C2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT127), .B1(new_n1230), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1230), .A2(new_n1256), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1238), .A2(new_n1259), .A3(KEYINPUT63), .A4(new_n1229), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1255), .A2(new_n1257), .A3(new_n1258), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1252), .A2(new_n1261), .ZN(G405));
  NAND2_X1  g1062(.A1(G375), .A2(new_n1211), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1229), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1215), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1263), .B2(new_n1215), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1251), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1267), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(new_n1250), .A3(new_n1265), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(G402));
endmodule


