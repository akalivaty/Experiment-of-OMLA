

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n571), .A2(n570), .ZN(n684) );
  AND2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n914) );
  AND2_X1 U559 ( .A1(n547), .A2(n546), .ZN(n543) );
  AND2_X1 U560 ( .A1(n544), .A2(KEYINPUT64), .ZN(n542) );
  XNOR2_X1 U561 ( .A(n536), .B(KEYINPUT28), .ZN(n535) );
  AND2_X1 U562 ( .A1(n530), .A2(n534), .ZN(n529) );
  BUF_X1 U563 ( .A(n748), .Z(n758) );
  AND2_X1 U564 ( .A1(n602), .A2(n601), .ZN(n719) );
  BUF_X1 U565 ( .A(n615), .Z(n606) );
  NAND2_X1 U566 ( .A1(n603), .A2(n557), .ZN(n556) );
  OR2_X2 U567 ( .A1(n781), .A2(KEYINPUT33), .ZN(n522) );
  INV_X4 U568 ( .A(G2105), .ZN(n603) );
  NAND2_X2 U569 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X2 U570 ( .A(n558), .B(n556), .ZN(n615) );
  NAND2_X1 U571 ( .A1(G299), .A2(KEYINPUT92), .ZN(n534) );
  NAND2_X1 U572 ( .A1(n528), .A2(n533), .ZN(n527) );
  INV_X1 U573 ( .A(n1013), .ZN(n551) );
  AND2_X1 U574 ( .A1(n1013), .A2(KEYINPUT97), .ZN(n553) );
  INV_X1 U575 ( .A(n792), .ZN(n555) );
  XOR2_X1 U576 ( .A(KEYINPUT31), .B(n755), .Z(n756) );
  INV_X1 U577 ( .A(G2104), .ZN(n557) );
  XOR2_X1 U578 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U579 ( .A1(n529), .A2(n527), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n551), .A2(n780), .ZN(n550) );
  INV_X1 U581 ( .A(n807), .ZN(n721) );
  NAND2_X1 U582 ( .A1(n549), .A2(n554), .ZN(n547) );
  NAND2_X1 U583 ( .A1(G1976), .A2(G288), .ZN(n1013) );
  NAND2_X1 U584 ( .A1(n914), .A2(G113), .ZN(n597) );
  NAND2_X1 U585 ( .A1(n911), .A2(G101), .ZN(n605) );
  XNOR2_X1 U586 ( .A(n581), .B(n580), .ZN(G168) );
  INV_X1 U587 ( .A(KEYINPUT7), .ZN(n579) );
  AND2_X1 U588 ( .A1(n524), .A2(n995), .ZN(n521) );
  AND2_X1 U589 ( .A1(n794), .A2(n793), .ZN(n523) );
  OR2_X1 U590 ( .A1(n792), .A2(n783), .ZN(n524) );
  AND2_X1 U591 ( .A1(n555), .A2(n550), .ZN(n525) );
  AND2_X1 U592 ( .A1(n780), .A2(n554), .ZN(n526) );
  INV_X1 U593 ( .A(KEYINPUT64), .ZN(n554) );
  INV_X1 U594 ( .A(n741), .ZN(n528) );
  NAND2_X1 U595 ( .A1(n741), .A2(KEYINPUT92), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n531), .A2(n535), .ZN(n743) );
  NAND2_X1 U597 ( .A1(n740), .A2(n532), .ZN(n531) );
  NOR2_X1 U598 ( .A1(G299), .A2(KEYINPUT92), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n741), .A2(G299), .ZN(n536) );
  NAND2_X1 U600 ( .A1(n537), .A2(n830), .ZN(n844) );
  XNOR2_X1 U601 ( .A(n539), .B(n538), .ZN(n537) );
  INV_X1 U602 ( .A(KEYINPUT99), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n540), .A2(n523), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n522), .A2(n521), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n543), .A2(n541), .ZN(n781) );
  NAND2_X1 U606 ( .A1(n545), .A2(n542), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n548), .A2(n780), .ZN(n544) );
  INV_X1 U608 ( .A(n549), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n548), .A2(n526), .ZN(n546) );
  INV_X1 U610 ( .A(n779), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n552), .A2(n525), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n779), .A2(n553), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n615), .A2(G137), .ZN(n598) );
  XNOR2_X2 U614 ( .A(KEYINPUT66), .B(KEYINPUT17), .ZN(n558) );
  XOR2_X1 U615 ( .A(KEYINPUT93), .B(KEYINPUT30), .Z(n559) );
  INV_X1 U616 ( .A(KEYINPUT26), .ZN(n722) );
  NOR2_X1 U617 ( .A1(n1004), .A2(n726), .ZN(n731) );
  XNOR2_X1 U618 ( .A(n750), .B(n559), .ZN(n751) );
  INV_X1 U619 ( .A(KEYINPUT29), .ZN(n742) );
  INV_X1 U620 ( .A(KEYINPUT95), .ZN(n764) );
  AND2_X1 U621 ( .A1(G40), .A2(n717), .ZN(n718) );
  NAND2_X1 U622 ( .A1(n688), .A2(G54), .ZN(n640) );
  INV_X1 U623 ( .A(KEYINPUT77), .ZN(n645) );
  XNOR2_X1 U624 ( .A(n645), .B(KEYINPUT15), .ZN(n646) );
  INV_X1 U625 ( .A(KEYINPUT5), .ZN(n575) );
  NOR2_X2 U626 ( .A1(n571), .A2(G651), .ZN(n688) );
  INV_X1 U627 ( .A(KEYINPUT23), .ZN(n604) );
  XNOR2_X1 U628 ( .A(n579), .B(KEYINPUT78), .ZN(n580) );
  XNOR2_X1 U629 ( .A(n605), .B(n604), .ZN(n717) );
  NOR2_X1 U630 ( .A1(n596), .A2(n595), .ZN(G171) );
  INV_X1 U631 ( .A(G651), .ZN(n570) );
  NOR2_X1 U632 ( .A1(G543), .A2(n570), .ZN(n560) );
  XOR2_X2 U633 ( .A(KEYINPUT1), .B(n560), .Z(n681) );
  XOR2_X1 U634 ( .A(G543), .B(KEYINPUT0), .Z(n571) );
  NAND2_X1 U635 ( .A1(G49), .A2(n688), .ZN(n562) );
  NAND2_X1 U636 ( .A1(G74), .A2(G651), .ZN(n561) );
  NAND2_X1 U637 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U638 ( .A1(n681), .A2(n563), .ZN(n564) );
  XNOR2_X1 U639 ( .A(n564), .B(KEYINPUT80), .ZN(n566) );
  NAND2_X1 U640 ( .A1(G87), .A2(n571), .ZN(n565) );
  NAND2_X1 U641 ( .A1(n566), .A2(n565), .ZN(G288) );
  NAND2_X1 U642 ( .A1(G63), .A2(n681), .ZN(n568) );
  NAND2_X1 U643 ( .A1(G51), .A2(n688), .ZN(n567) );
  NAND2_X1 U644 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U645 ( .A(n569), .B(KEYINPUT6), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G76), .A2(n684), .ZN(n574) );
  NOR2_X1 U647 ( .A1(G651), .A2(G543), .ZN(n680) );
  NAND2_X1 U648 ( .A1(n680), .A2(G89), .ZN(n572) );
  XNOR2_X1 U649 ( .A(n572), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U651 ( .A(n576), .B(n575), .ZN(n577) );
  NOR2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U653 ( .A1(G91), .A2(n680), .ZN(n583) );
  NAND2_X1 U654 ( .A1(G65), .A2(n681), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G78), .A2(n684), .ZN(n584) );
  XNOR2_X1 U657 ( .A(KEYINPUT71), .B(n584), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n688), .A2(G53), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(G299) );
  NAND2_X1 U661 ( .A1(G64), .A2(n681), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G52), .A2(n688), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n680), .A2(G90), .ZN(n591) );
  XOR2_X1 U665 ( .A(KEYINPUT69), .B(n591), .Z(n593) );
  NAND2_X1 U666 ( .A1(n684), .A2(G77), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U668 ( .A(KEYINPUT9), .B(n594), .Z(n595) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n599), .B(KEYINPUT67), .ZN(n602) );
  NOR2_X4 U671 ( .A1(G2104), .A2(n603), .ZN(n915) );
  NAND2_X1 U672 ( .A1(G125), .A2(n915), .ZN(n600) );
  XOR2_X1 U673 ( .A(KEYINPUT65), .B(n600), .Z(n601) );
  AND2_X2 U674 ( .A1(n603), .A2(G2104), .ZN(n911) );
  AND2_X1 U675 ( .A1(n719), .A2(n717), .ZN(G160) );
  NAND2_X1 U676 ( .A1(G111), .A2(n914), .ZN(n608) );
  NAND2_X1 U677 ( .A1(G135), .A2(n606), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U679 ( .A1(n915), .A2(G123), .ZN(n609) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n609), .Z(n610) );
  NOR2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n911), .A2(G99), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n973) );
  XNOR2_X1 U684 ( .A(G2096), .B(n973), .ZN(n614) );
  OR2_X1 U685 ( .A1(G2100), .A2(n614), .ZN(G156) );
  INV_X1 U686 ( .A(G132), .ZN(G219) );
  INV_X1 U687 ( .A(G82), .ZN(G220) );
  NAND2_X1 U688 ( .A1(G102), .A2(n911), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G138), .A2(n615), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT84), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G114), .A2(n914), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G126), .A2(n915), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n720) );
  BUF_X1 U696 ( .A(n720), .Z(G164) );
  NAND2_X1 U697 ( .A1(G94), .A2(G452), .ZN(n623) );
  XOR2_X1 U698 ( .A(KEYINPUT70), .B(n623), .Z(G173) );
  NAND2_X1 U699 ( .A1(G7), .A2(G661), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n624), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U701 ( .A(G223), .ZN(n856) );
  NAND2_X1 U702 ( .A1(n856), .A2(G567), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT11), .ZN(n626) );
  XNOR2_X1 U704 ( .A(KEYINPUT73), .B(n626), .ZN(G234) );
  NAND2_X1 U705 ( .A1(G56), .A2(n681), .ZN(n627) );
  XOR2_X1 U706 ( .A(KEYINPUT14), .B(n627), .Z(n633) );
  NAND2_X1 U707 ( .A1(n680), .A2(G81), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n628), .B(KEYINPUT12), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G68), .A2(n684), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U711 ( .A(KEYINPUT13), .B(n631), .Z(n632) );
  NOR2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n688), .A2(G43), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n1004) );
  INV_X1 U715 ( .A(G860), .ZN(n652) );
  NOR2_X1 U716 ( .A1(n1004), .A2(n652), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT74), .B(n636), .Z(G153) );
  INV_X1 U718 ( .A(G868), .ZN(n698) );
  NOR2_X1 U719 ( .A1(n698), .A2(G171), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n637), .B(KEYINPUT75), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n681), .A2(G66), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G92), .A2(n680), .ZN(n639) );
  NAND2_X1 U723 ( .A1(G79), .A2(n684), .ZN(n638) );
  NAND2_X1 U724 ( .A1(n639), .A2(n638), .ZN(n642) );
  XOR2_X1 U725 ( .A(KEYINPUT76), .B(n640), .Z(n641) );
  NOR2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n647) );
  XNOR2_X2 U728 ( .A(n647), .B(n646), .ZN(n998) );
  OR2_X1 U729 ( .A1(G868), .A2(n998), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(G284) );
  NAND2_X1 U731 ( .A1(G868), .A2(G286), .ZN(n651) );
  NAND2_X1 U732 ( .A1(G299), .A2(n698), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(G297) );
  NAND2_X1 U734 ( .A1(n652), .A2(G559), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n653), .A2(n998), .ZN(n654) );
  XNOR2_X1 U736 ( .A(n654), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U737 ( .A1(G868), .A2(n1004), .ZN(n655) );
  XOR2_X1 U738 ( .A(KEYINPUT79), .B(n655), .Z(n658) );
  NAND2_X1 U739 ( .A1(G868), .A2(n998), .ZN(n656) );
  NOR2_X1 U740 ( .A1(G559), .A2(n656), .ZN(n657) );
  NOR2_X1 U741 ( .A1(n658), .A2(n657), .ZN(G282) );
  NAND2_X1 U742 ( .A1(G559), .A2(n998), .ZN(n659) );
  XNOR2_X1 U743 ( .A(n659), .B(n1004), .ZN(n696) );
  NOR2_X1 U744 ( .A1(n696), .A2(G860), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G67), .A2(n681), .ZN(n661) );
  NAND2_X1 U746 ( .A1(G55), .A2(n688), .ZN(n660) );
  NAND2_X1 U747 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U748 ( .A1(G93), .A2(n680), .ZN(n663) );
  NAND2_X1 U749 ( .A1(G80), .A2(n684), .ZN(n662) );
  NAND2_X1 U750 ( .A1(n663), .A2(n662), .ZN(n664) );
  OR2_X1 U751 ( .A1(n665), .A2(n664), .ZN(n699) );
  XOR2_X1 U752 ( .A(n666), .B(n699), .Z(G145) );
  NAND2_X1 U753 ( .A1(G88), .A2(n680), .ZN(n668) );
  NAND2_X1 U754 ( .A1(G75), .A2(n684), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n668), .A2(n667), .ZN(n672) );
  NAND2_X1 U756 ( .A1(G62), .A2(n681), .ZN(n670) );
  NAND2_X1 U757 ( .A1(G50), .A2(n688), .ZN(n669) );
  NAND2_X1 U758 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U759 ( .A1(n672), .A2(n671), .ZN(G166) );
  NAND2_X1 U760 ( .A1(G85), .A2(n680), .ZN(n674) );
  NAND2_X1 U761 ( .A1(G72), .A2(n684), .ZN(n673) );
  NAND2_X1 U762 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U763 ( .A1(G47), .A2(n688), .ZN(n675) );
  XOR2_X1 U764 ( .A(KEYINPUT68), .B(n675), .Z(n676) );
  NOR2_X1 U765 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U766 ( .A1(n681), .A2(G60), .ZN(n678) );
  NAND2_X1 U767 ( .A1(n679), .A2(n678), .ZN(G290) );
  NAND2_X1 U768 ( .A1(G86), .A2(n680), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G61), .A2(n681), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U771 ( .A1(n684), .A2(G73), .ZN(n685) );
  XOR2_X1 U772 ( .A(KEYINPUT2), .B(n685), .Z(n686) );
  NOR2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n688), .A2(G48), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(G305) );
  XNOR2_X1 U776 ( .A(G166), .B(KEYINPUT19), .ZN(n695) );
  XOR2_X1 U777 ( .A(G290), .B(G299), .Z(n691) );
  XNOR2_X1 U778 ( .A(G288), .B(n691), .ZN(n692) );
  XOR2_X1 U779 ( .A(n699), .B(n692), .Z(n693) );
  XNOR2_X1 U780 ( .A(n693), .B(G305), .ZN(n694) );
  XNOR2_X1 U781 ( .A(n695), .B(n694), .ZN(n865) );
  XNOR2_X1 U782 ( .A(n696), .B(n865), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n697), .A2(G868), .ZN(n701) );
  NAND2_X1 U784 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U785 ( .A1(n701), .A2(n700), .ZN(G295) );
  NAND2_X1 U786 ( .A1(G2078), .A2(G2084), .ZN(n702) );
  XOR2_X1 U787 ( .A(KEYINPUT20), .B(n702), .Z(n703) );
  NAND2_X1 U788 ( .A1(G2090), .A2(n703), .ZN(n704) );
  XNOR2_X1 U789 ( .A(KEYINPUT21), .B(n704), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n705), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U791 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U792 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  NOR2_X1 U793 ( .A1(G220), .A2(G219), .ZN(n706) );
  XNOR2_X1 U794 ( .A(KEYINPUT22), .B(n706), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n707), .A2(G96), .ZN(n708) );
  NOR2_X1 U796 ( .A1(n708), .A2(G218), .ZN(n709) );
  XNOR2_X1 U797 ( .A(n709), .B(KEYINPUT81), .ZN(n863) );
  NAND2_X1 U798 ( .A1(G2106), .A2(n863), .ZN(n710) );
  XNOR2_X1 U799 ( .A(KEYINPUT82), .B(n710), .ZN(n714) );
  NAND2_X1 U800 ( .A1(G108), .A2(G120), .ZN(n711) );
  NOR2_X1 U801 ( .A1(G237), .A2(n711), .ZN(n712) );
  NAND2_X1 U802 ( .A1(G69), .A2(n712), .ZN(n864) );
  NAND2_X1 U803 ( .A1(G567), .A2(n864), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n935) );
  NAND2_X1 U805 ( .A1(G483), .A2(G661), .ZN(n715) );
  NOR2_X1 U806 ( .A1(n935), .A2(n715), .ZN(n716) );
  XOR2_X1 U807 ( .A(KEYINPUT83), .B(n716), .Z(n862) );
  NAND2_X1 U808 ( .A1(n862), .A2(G36), .ZN(G176) );
  INV_X1 U809 ( .A(G166), .ZN(G303) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n807) );
  NOR2_X2 U811 ( .A1(n720), .A2(G1384), .ZN(n808) );
  NAND2_X2 U812 ( .A1(n721), .A2(n808), .ZN(n748) );
  INV_X1 U813 ( .A(G1996), .ZN(n1026) );
  NOR2_X1 U814 ( .A1(n748), .A2(n1026), .ZN(n723) );
  XNOR2_X1 U815 ( .A(n723), .B(n722), .ZN(n725) );
  NAND2_X1 U816 ( .A1(n758), .A2(G1341), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n731), .A2(n998), .ZN(n730) );
  XNOR2_X2 U819 ( .A(n748), .B(KEYINPUT91), .ZN(n734) );
  NAND2_X1 U820 ( .A1(G2067), .A2(n734), .ZN(n728) );
  NAND2_X1 U821 ( .A1(G1348), .A2(n758), .ZN(n727) );
  NAND2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n733) );
  OR2_X1 U824 ( .A1(n998), .A2(n731), .ZN(n732) );
  NAND2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n740) );
  NAND2_X1 U826 ( .A1(n734), .A2(G2072), .ZN(n736) );
  INV_X1 U827 ( .A(KEYINPUT27), .ZN(n735) );
  XNOR2_X1 U828 ( .A(n736), .B(n735), .ZN(n739) );
  INV_X1 U829 ( .A(n734), .ZN(n737) );
  NAND2_X1 U830 ( .A1(G1956), .A2(n737), .ZN(n738) );
  XNOR2_X1 U831 ( .A(n743), .B(n742), .ZN(n747) );
  INV_X1 U832 ( .A(G1961), .ZN(n999) );
  NAND2_X1 U833 ( .A1(n999), .A2(n758), .ZN(n745) );
  XNOR2_X1 U834 ( .A(G2078), .B(KEYINPUT25), .ZN(n1025) );
  NAND2_X1 U835 ( .A1(n734), .A2(n1025), .ZN(n744) );
  NAND2_X1 U836 ( .A1(n745), .A2(n744), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n752), .A2(G171), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n757) );
  NAND2_X1 U839 ( .A1(G8), .A2(n748), .ZN(n792) );
  NOR2_X1 U840 ( .A1(G1966), .A2(n792), .ZN(n770) );
  NOR2_X1 U841 ( .A1(G2084), .A2(n758), .ZN(n771) );
  NOR2_X1 U842 ( .A1(n770), .A2(n771), .ZN(n749) );
  NAND2_X1 U843 ( .A1(n749), .A2(G8), .ZN(n750) );
  NOR2_X1 U844 ( .A1(G168), .A2(n751), .ZN(n754) );
  NOR2_X1 U845 ( .A1(G171), .A2(n752), .ZN(n753) );
  NOR2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n768) );
  NAND2_X1 U848 ( .A1(n768), .A2(G286), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G1971), .A2(n792), .ZN(n760) );
  NOR2_X1 U850 ( .A1(G2090), .A2(n758), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n761), .A2(G303), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U854 ( .A(n765), .B(n764), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n766), .A2(G8), .ZN(n767) );
  XNOR2_X1 U856 ( .A(n767), .B(KEYINPUT32), .ZN(n776) );
  INV_X1 U857 ( .A(n768), .ZN(n769) );
  NOR2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U861 ( .A(KEYINPUT94), .B(n774), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U863 ( .A(n777), .B(KEYINPUT96), .ZN(n784) );
  NOR2_X1 U864 ( .A1(G1976), .A2(G288), .ZN(n782) );
  NOR2_X1 U865 ( .A1(G1971), .A2(G303), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n782), .A2(n778), .ZN(n1014) );
  NAND2_X1 U867 ( .A1(n784), .A2(n1014), .ZN(n779) );
  INV_X1 U868 ( .A(KEYINPUT97), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n782), .A2(KEYINPUT33), .ZN(n783) );
  XOR2_X1 U870 ( .A(G1981), .B(G305), .Z(n995) );
  NOR2_X1 U871 ( .A1(G2090), .A2(G303), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G8), .A2(n785), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n784), .A2(n786), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(KEYINPUT98), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n788), .A2(n792), .ZN(n794) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U877 ( .A(n789), .B(KEYINPUT90), .Z(n790) );
  XNOR2_X1 U878 ( .A(KEYINPUT24), .B(n790), .ZN(n791) );
  OR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U880 ( .A(KEYINPUT37), .B(G2067), .ZN(n839) );
  NAND2_X1 U881 ( .A1(G116), .A2(n914), .ZN(n796) );
  NAND2_X1 U882 ( .A1(G128), .A2(n915), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n798) );
  XOR2_X1 U884 ( .A(KEYINPUT87), .B(KEYINPUT35), .Z(n797) );
  XNOR2_X1 U885 ( .A(n798), .B(n797), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G140), .A2(n606), .ZN(n799) );
  XNOR2_X1 U887 ( .A(n799), .B(KEYINPUT86), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G104), .A2(n911), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U890 ( .A(KEYINPUT34), .B(n802), .Z(n803) );
  NAND2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U892 ( .A(KEYINPUT36), .B(n805), .Z(n922) );
  OR2_X1 U893 ( .A1(n839), .A2(n922), .ZN(n806) );
  XNOR2_X1 U894 ( .A(KEYINPUT88), .B(n806), .ZN(n978) );
  XOR2_X1 U895 ( .A(G1986), .B(G290), .Z(n1015) );
  NAND2_X1 U896 ( .A1(n978), .A2(n1015), .ZN(n810) );
  NOR2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U898 ( .A(KEYINPUT85), .B(n809), .Z(n841) );
  NAND2_X1 U899 ( .A1(n810), .A2(n841), .ZN(n829) );
  NAND2_X1 U900 ( .A1(G95), .A2(n911), .ZN(n812) );
  NAND2_X1 U901 ( .A1(G131), .A2(n606), .ZN(n811) );
  NAND2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G107), .A2(n914), .ZN(n814) );
  NAND2_X1 U904 ( .A1(G119), .A2(n915), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U907 ( .A(n817), .B(KEYINPUT89), .Z(n899) );
  INV_X1 U908 ( .A(G1991), .ZN(n1021) );
  NOR2_X1 U909 ( .A1(n899), .A2(n1021), .ZN(n826) );
  NAND2_X1 U910 ( .A1(n915), .A2(G129), .ZN(n819) );
  NAND2_X1 U911 ( .A1(G141), .A2(n606), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n822) );
  NAND2_X1 U913 ( .A1(G105), .A2(n911), .ZN(n820) );
  XOR2_X1 U914 ( .A(KEYINPUT38), .B(n820), .Z(n821) );
  NOR2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n914), .A2(G117), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n900) );
  AND2_X1 U918 ( .A1(n900), .A2(G1996), .ZN(n825) );
  NOR2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n972) );
  INV_X1 U920 ( .A(n841), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n972), .A2(n827), .ZN(n834) );
  INV_X1 U922 ( .A(n834), .ZN(n828) );
  AND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n837) );
  NOR2_X1 U925 ( .A1(G1996), .A2(n900), .ZN(n969) );
  AND2_X1 U926 ( .A1(n899), .A2(n1021), .ZN(n831) );
  XNOR2_X1 U927 ( .A(n831), .B(KEYINPUT100), .ZN(n976) );
  NOR2_X1 U928 ( .A1(G1986), .A2(G290), .ZN(n832) );
  NOR2_X1 U929 ( .A1(n976), .A2(n832), .ZN(n833) );
  NOR2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n969), .A2(n835), .ZN(n836) );
  XNOR2_X1 U932 ( .A(n837), .B(n836), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n838), .A2(n978), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n839), .A2(n922), .ZN(n982) );
  NAND2_X1 U935 ( .A1(n840), .A2(n982), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U938 ( .A(n845), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U939 ( .A(G2454), .B(G2451), .ZN(n854) );
  XNOR2_X1 U940 ( .A(G2430), .B(G2446), .ZN(n852) );
  XOR2_X1 U941 ( .A(G2435), .B(G2427), .Z(n847) );
  XNOR2_X1 U942 ( .A(KEYINPUT102), .B(G2438), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U944 ( .A(n848), .B(G2443), .Z(n850) );
  XNOR2_X1 U945 ( .A(G1341), .B(G1348), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U947 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U948 ( .A(n854), .B(n853), .ZN(n855) );
  NAND2_X1 U949 ( .A1(n855), .A2(G14), .ZN(n938) );
  XNOR2_X1 U950 ( .A(KEYINPUT103), .B(n938), .ZN(G401) );
  NAND2_X1 U951 ( .A1(G2106), .A2(n856), .ZN(G217) );
  INV_X1 U952 ( .A(G661), .ZN(n858) );
  NAND2_X1 U953 ( .A1(G2), .A2(G15), .ZN(n857) );
  NOR2_X1 U954 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U955 ( .A(KEYINPUT104), .B(n859), .Z(G259) );
  NAND2_X1 U956 ( .A1(G3), .A2(G1), .ZN(n860) );
  XOR2_X1 U957 ( .A(KEYINPUT105), .B(n860), .Z(n861) );
  NAND2_X1 U958 ( .A1(n862), .A2(n861), .ZN(G188) );
  INV_X1 U960 ( .A(G120), .ZN(G236) );
  INV_X1 U961 ( .A(G108), .ZN(G238) );
  INV_X1 U962 ( .A(G96), .ZN(G221) );
  INV_X1 U963 ( .A(G69), .ZN(G235) );
  NOR2_X1 U964 ( .A1(n864), .A2(n863), .ZN(G325) );
  INV_X1 U965 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U966 ( .A(n998), .B(G286), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n868) );
  XOR2_X1 U968 ( .A(n1004), .B(G171), .Z(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n869) );
  NOR2_X1 U970 ( .A1(G37), .A2(n869), .ZN(G397) );
  XOR2_X1 U971 ( .A(G1981), .B(G1966), .Z(n871) );
  XNOR2_X1 U972 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n881) );
  XOR2_X1 U974 ( .A(KEYINPUT109), .B(G2474), .Z(n873) );
  XNOR2_X1 U975 ( .A(G1956), .B(KEYINPUT107), .ZN(n872) );
  XNOR2_X1 U976 ( .A(n873), .B(n872), .ZN(n877) );
  XOR2_X1 U977 ( .A(G1976), .B(G1971), .Z(n875) );
  XNOR2_X1 U978 ( .A(G1986), .B(G1961), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U980 ( .A(n877), .B(n876), .Z(n879) );
  XNOR2_X1 U981 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n878) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U983 ( .A(n881), .B(n880), .Z(G229) );
  XOR2_X1 U984 ( .A(G2096), .B(KEYINPUT106), .Z(n883) );
  XNOR2_X1 U985 ( .A(G2090), .B(KEYINPUT43), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(n884), .B(KEYINPUT42), .Z(n886) );
  XNOR2_X1 U988 ( .A(G2067), .B(G2072), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U990 ( .A(G2678), .B(G2100), .Z(n888) );
  XNOR2_X1 U991 ( .A(G2078), .B(G2084), .ZN(n887) );
  XNOR2_X1 U992 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(G227) );
  NAND2_X1 U994 ( .A1(G124), .A2(n915), .ZN(n891) );
  XNOR2_X1 U995 ( .A(n891), .B(KEYINPUT44), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n606), .A2(G136), .ZN(n892) );
  XNOR2_X1 U997 ( .A(n892), .B(KEYINPUT110), .ZN(n893) );
  NAND2_X1 U998 ( .A1(n894), .A2(n893), .ZN(n898) );
  NAND2_X1 U999 ( .A1(G100), .A2(n911), .ZN(n896) );
  NAND2_X1 U1000 ( .A1(G112), .A2(n914), .ZN(n895) );
  NAND2_X1 U1001 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U1002 ( .A1(n898), .A2(n897), .ZN(G162) );
  XOR2_X1 U1003 ( .A(n900), .B(n899), .Z(n901) );
  XNOR2_X1 U1004 ( .A(n901), .B(G162), .ZN(n926) );
  XNOR2_X1 U1005 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n606), .ZN(n904) );
  NAND2_X1 U1007 ( .A1(n911), .A2(G106), .ZN(n902) );
  XOR2_X1 U1008 ( .A(KEYINPUT111), .B(n902), .Z(n903) );
  NAND2_X1 U1009 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1010 ( .A(n906), .B(n905), .Z(n910) );
  NAND2_X1 U1011 ( .A1(G118), .A2(n914), .ZN(n908) );
  NAND2_X1 U1012 ( .A1(G130), .A2(n915), .ZN(n907) );
  NAND2_X1 U1013 ( .A1(n908), .A2(n907), .ZN(n909) );
  NOR2_X1 U1014 ( .A1(n910), .A2(n909), .ZN(n924) );
  NAND2_X1 U1015 ( .A1(G103), .A2(n911), .ZN(n913) );
  NAND2_X1 U1016 ( .A1(G139), .A2(n606), .ZN(n912) );
  NAND2_X1 U1017 ( .A1(n913), .A2(n912), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(G115), .A2(n914), .ZN(n917) );
  NAND2_X1 U1019 ( .A1(G127), .A2(n915), .ZN(n916) );
  NAND2_X1 U1020 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1021 ( .A(KEYINPUT47), .B(n918), .Z(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1023 ( .A(KEYINPUT114), .B(n921), .Z(n984) );
  XOR2_X1 U1024 ( .A(n984), .B(n922), .Z(n923) );
  XNOR2_X1 U1025 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n926), .B(n925), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n928) );
  XNOR2_X1 U1028 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(n928), .B(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n973), .B(n929), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n931), .B(n930), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(G164), .B(G160), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(n933), .B(n932), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(G37), .A2(n934), .ZN(G395) );
  INV_X1 U1035 ( .A(n935), .ZN(G319) );
  NOR2_X1 U1036 ( .A1(G229), .A2(G227), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(KEYINPUT49), .B(n936), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(G397), .A2(n937), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(G319), .A2(n938), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(KEYINPUT116), .B(n939), .ZN(n940) );
  NOR2_X1 U1041 ( .A1(G395), .A2(n940), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(G225) );
  INV_X1 U1043 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1044 ( .A(n999), .B(G5), .ZN(n964) );
  XOR2_X1 U1045 ( .A(G1966), .B(G21), .Z(n950) );
  XNOR2_X1 U1046 ( .A(G1986), .B(G24), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n944) );
  XNOR2_X1 U1048 ( .A(G23), .B(G1976), .ZN(n943) );
  NOR2_X1 U1049 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1050 ( .A(KEYINPUT125), .B(n945), .ZN(n946) );
  NOR2_X1 U1051 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n948), .ZN(n949) );
  NAND2_X1 U1053 ( .A1(n950), .A2(n949), .ZN(n962) );
  XOR2_X1 U1054 ( .A(G1956), .B(G20), .Z(n953) );
  XOR2_X1 U1055 ( .A(G6), .B(KEYINPUT124), .Z(n951) );
  XNOR2_X1 U1056 ( .A(G1981), .B(n951), .ZN(n952) );
  NAND2_X1 U1057 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1058 ( .A(KEYINPUT59), .B(G1348), .Z(n954) );
  XNOR2_X1 U1059 ( .A(G4), .B(n954), .ZN(n955) );
  NOR2_X1 U1060 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1061 ( .A(G1341), .B(KEYINPUT123), .ZN(n957) );
  XNOR2_X1 U1062 ( .A(n957), .B(G19), .ZN(n958) );
  NAND2_X1 U1063 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1064 ( .A(KEYINPUT60), .B(n960), .ZN(n961) );
  NOR2_X1 U1065 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1066 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1067 ( .A(n965), .B(KEYINPUT61), .ZN(n966) );
  XNOR2_X1 U1068 ( .A(n966), .B(KEYINPUT126), .ZN(n967) );
  NOR2_X1 U1069 ( .A1(G16), .A2(n967), .ZN(n1049) );
  XOR2_X1 U1070 ( .A(G2090), .B(G162), .Z(n968) );
  NOR2_X1 U1071 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1072 ( .A(KEYINPUT51), .B(n970), .Z(n971) );
  NAND2_X1 U1073 ( .A1(n972), .A2(n971), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(G160), .B(G2084), .ZN(n974) );
  NAND2_X1 U1075 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1076 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1078 ( .A(KEYINPUT117), .B(n979), .Z(n980) );
  NOR2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n989) );
  XOR2_X1 U1081 ( .A(G164), .B(G2078), .Z(n986) );
  XNOR2_X1 U1082 ( .A(G2072), .B(n984), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1084 ( .A(KEYINPUT50), .B(n987), .Z(n988) );
  NOR2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1086 ( .A(KEYINPUT52), .B(n990), .ZN(n992) );
  INV_X1 U1087 ( .A(KEYINPUT55), .ZN(n991) );
  NAND2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1089 ( .A1(n993), .A2(G29), .ZN(n994) );
  XNOR2_X1 U1090 ( .A(KEYINPUT118), .B(n994), .ZN(n1047) );
  XOR2_X1 U1091 ( .A(KEYINPUT56), .B(G16), .Z(n1020) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G168), .ZN(n996) );
  NAND2_X1 U1093 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1094 ( .A(KEYINPUT57), .B(n997), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(n998), .B(G1348), .ZN(n1002) );
  XNOR2_X1 U1096 ( .A(G171), .B(KEYINPUT121), .ZN(n1000) );
  XNOR2_X1 U1097 ( .A(n1000), .B(n999), .ZN(n1001) );
  NAND2_X1 U1098 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1099 ( .A(n1003), .B(KEYINPUT122), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1004), .B(G1341), .ZN(n1006) );
  XNOR2_X1 U1101 ( .A(G299), .B(G1956), .ZN(n1005) );
  NOR2_X1 U1102 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  NAND2_X1 U1103 ( .A1(G1971), .A2(G303), .ZN(n1007) );
  NAND2_X1 U1104 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1105 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1106 ( .A1(n1012), .A2(n1011), .ZN(n1018) );
  AND2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  NAND2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1045) );
  XOR2_X1 U1111 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n1040) );
  XNOR2_X1 U1112 ( .A(G2090), .B(G35), .ZN(n1035) );
  XNOR2_X1 U1113 ( .A(G25), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1114 ( .A1(n1022), .A2(G28), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(G2067), .B(G26), .ZN(n1024) );
  XNOR2_X1 U1116 ( .A(G33), .B(G2072), .ZN(n1023) );
  NOR2_X1 U1117 ( .A1(n1024), .A2(n1023), .ZN(n1030) );
  XOR2_X1 U1118 ( .A(n1025), .B(G27), .Z(n1028) );
  XOR2_X1 U1119 ( .A(n1026), .B(G32), .Z(n1027) );
  NOR2_X1 U1120 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1121 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1122 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1123 ( .A(KEYINPUT53), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1124 ( .A1(n1035), .A2(n1034), .ZN(n1038) );
  XOR2_X1 U1125 ( .A(G2084), .B(G34), .Z(n1036) );
  XNOR2_X1 U1126 ( .A(KEYINPUT54), .B(n1036), .ZN(n1037) );
  NAND2_X1 U1127 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1128 ( .A(n1040), .B(n1039), .ZN(n1041) );
  OR2_X1 U1129 ( .A1(G29), .A2(n1041), .ZN(n1042) );
  NAND2_X1 U1130 ( .A1(G11), .A2(n1042), .ZN(n1043) );
  XNOR2_X1 U1131 ( .A(KEYINPUT120), .B(n1043), .ZN(n1044) );
  NOR2_X1 U1132 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NAND2_X1 U1133 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NOR2_X1 U1134 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XOR2_X1 U1135 ( .A(KEYINPUT62), .B(n1050), .Z(n1051) );
  XNOR2_X1 U1136 ( .A(KEYINPUT127), .B(n1051), .ZN(G311) );
  INV_X1 U1137 ( .A(G311), .ZN(G150) );
  INV_X1 U1138 ( .A(G171), .ZN(G301) );
endmodule

