//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT65), .A2(G116), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT65), .A2(G116), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G119), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  INV_X1    g006(.A(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT2), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n190), .A2(new_n192), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n190), .B2(new_n192), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  AND4_X1   g019(.A1(new_n201), .A2(new_n203), .A3(new_n205), .A4(G128), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n207), .A2(G128), .B1(new_n203), .B2(new_n205), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n211), .A2(G137), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G134), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n209), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G131), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n203), .A2(new_n205), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G128), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n224), .A2(new_n217), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT30), .B1(new_n222), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n224), .A2(new_n217), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT30), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n217), .B(new_n220), .C1(new_n206), .C2(new_n208), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n200), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n236), .A2(new_n200), .A3(new_n238), .ZN(new_n241));
  NOR2_X1   g055(.A1(G237), .A2(G953), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G210), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT27), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(G101), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR4_X1   g061(.A1(new_n240), .A2(KEYINPUT31), .A3(new_n241), .A4(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n249));
  INV_X1    g063(.A(new_n199), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n190), .A2(new_n192), .A3(new_n197), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n222), .B2(new_n232), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n236), .A2(new_n200), .A3(new_n238), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n249), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n254), .A2(new_n249), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n247), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT31), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n240), .A2(new_n241), .A3(new_n247), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n248), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G472), .A2(G902), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n187), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n233), .A2(new_n239), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n241), .B1(new_n266), .B2(new_n252), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n257), .A2(new_n258), .B1(new_n267), .B2(new_n246), .ZN(new_n268));
  OAI211_X1 g082(.A(KEYINPUT32), .B(new_n263), .C1(new_n268), .C2(new_n248), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n247), .B1(new_n240), .B2(new_n241), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n200), .B1(new_n236), .B2(new_n238), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT28), .B1(new_n241), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n254), .A2(new_n249), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n246), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n270), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n274), .B2(new_n275), .ZN(new_n278));
  OAI21_X1  g092(.A(G472), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n265), .A2(new_n269), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n265), .A2(new_n282), .A3(new_n269), .A4(new_n279), .ZN(new_n283));
  INV_X1    g097(.A(G234), .ZN(new_n284));
  OAI21_X1  g098(.A(G217), .B1(new_n284), .B2(G902), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT67), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n288));
  XNOR2_X1  g102(.A(G119), .B(G128), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT24), .B(G110), .Z(new_n292));
  NAND2_X1  g106(.A1(new_n191), .A2(G128), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT23), .A2(G119), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n191), .A2(G128), .ZN(new_n295));
  OAI221_X1 g109(.A(new_n293), .B1(G128), .B2(new_n294), .C1(new_n295), .C2(KEYINPUT23), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n291), .A2(new_n292), .B1(G110), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G125), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G140), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(KEYINPUT69), .A3(G125), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(KEYINPUT16), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT16), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n305), .A2(new_n202), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n202), .B1(new_n305), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n297), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n291), .A2(new_n292), .B1(G110), .B2(new_n296), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n307), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G146), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n299), .A2(new_n301), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n202), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT22), .B(G137), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(G221), .A3(G234), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n318), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n310), .A2(new_n316), .A3(new_n321), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n288), .B1(new_n325), .B2(G902), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n323), .A2(KEYINPUT25), .A3(new_n277), .A4(new_n324), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n287), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n325), .A2(G902), .A3(new_n286), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n281), .A2(new_n283), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G104), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G107), .ZN(new_n333));
  INV_X1    g147(.A(G107), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G104), .ZN(new_n335));
  OAI21_X1  g149(.A(G101), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(new_n332), .B2(G107), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n334), .A3(G104), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(G107), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT72), .B(G101), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n336), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n226), .A2(G128), .A3(new_n207), .ZN(new_n344));
  INV_X1    g158(.A(new_n208), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(KEYINPUT72), .A2(G101), .ZN(new_n347));
  NOR2_X1   g161(.A1(KEYINPUT72), .A2(G101), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n349), .A2(new_n340), .A3(new_n337), .A4(new_n339), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n336), .C1(new_n206), .C2(new_n208), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT12), .A3(new_n234), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n352), .A2(KEYINPUT74), .A3(KEYINPUT12), .A4(new_n234), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n234), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT12), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n355), .A2(new_n359), .A3(new_n362), .A4(new_n356), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n341), .A2(G101), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(new_n350), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT4), .B1(new_n341), .B2(G101), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n235), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n234), .A2(KEYINPUT73), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT73), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n224), .A2(new_n370), .A3(new_n217), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n343), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n345), .A2(new_n344), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT10), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n351), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n368), .A2(new_n372), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n319), .A2(G227), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT71), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n361), .A2(new_n363), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n368), .A2(new_n375), .A3(new_n377), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n234), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n382), .B1(new_n387), .B2(new_n378), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G469), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n277), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n277), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n382), .B1(new_n360), .B2(new_n378), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n387), .A2(new_n378), .A3(new_n382), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n392), .B(new_n394), .C1(new_n398), .C2(new_n391), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT9), .B(G234), .ZN(new_n400));
  OAI21_X1  g214(.A(G221), .B1(new_n400), .B2(G902), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT70), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G214), .B1(G237), .B2(G902), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G122), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n252), .B1(new_n366), .B2(new_n367), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n190), .A2(KEYINPUT5), .A3(new_n192), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n191), .A3(G116), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n193), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n408), .B(new_n412), .C1(new_n411), .C2(new_n410), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n373), .A3(new_n251), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n406), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n414), .A3(new_n406), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n319), .A2(G224), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n419), .B(KEYINPUT79), .Z(new_n420));
  NAND3_X1  g234(.A1(new_n227), .A2(new_n231), .A3(G125), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n374), .B2(G125), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT78), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT78), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n420), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n209), .A2(new_n300), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n427), .B2(new_n421), .ZN(new_n428));
  INV_X1    g242(.A(new_n425), .ZN(new_n429));
  INV_X1    g243(.A(new_n420), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n415), .A2(KEYINPUT77), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT77), .B1(new_n415), .B2(new_n433), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n418), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n423), .A2(KEYINPUT7), .A3(new_n425), .A4(new_n419), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n406), .B(KEYINPUT8), .ZN(new_n438));
  INV_X1    g252(.A(new_n414), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n373), .B1(new_n413), .B2(new_n251), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n419), .A2(KEYINPUT7), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n422), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n437), .A2(new_n441), .A3(new_n417), .A4(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n444), .A2(new_n277), .ZN(new_n445));
  OAI21_X1  g259(.A(G210), .B1(G237), .B2(G902), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n436), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n436), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n405), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n404), .A2(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n242), .A2(G143), .A3(G214), .ZN(new_n451));
  AOI21_X1  g265(.A(G143), .B1(new_n242), .B2(G214), .ZN(new_n452));
  OAI21_X1  g266(.A(G131), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n454));
  INV_X1    g268(.A(G237), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n319), .A3(G214), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n204), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n242), .A2(G143), .A3(G214), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n215), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT81), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n453), .A2(new_n459), .A3(new_n462), .A4(new_n454), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT80), .B1(new_n308), .B2(new_n309), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n305), .A2(new_n202), .A3(new_n307), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n313), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n457), .A2(new_n458), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT17), .A3(G131), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n464), .A2(new_n465), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G113), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n332), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT18), .A2(G131), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n469), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n303), .A2(new_n304), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n315), .B1(new_n476), .B2(new_n202), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n453), .A2(new_n459), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n314), .A2(KEYINPUT19), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n476), .B2(KEYINPUT19), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n313), .B(new_n480), .C1(new_n482), .C2(G146), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n478), .ZN(new_n484));
  INV_X1    g298(.A(new_n473), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT20), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT82), .B1(G475), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NOR3_X1   g306(.A1(KEYINPUT82), .A2(G475), .A3(G902), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT20), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT83), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n487), .A2(KEYINPUT83), .A3(new_n494), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n471), .A2(new_n478), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n473), .ZN(new_n501));
  OAI21_X1  g315(.A(G475), .B1(new_n501), .B2(G902), .ZN(new_n502));
  XOR2_X1   g316(.A(G128), .B(G143), .Z(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(G134), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n188), .A2(G122), .A3(new_n189), .ZN(new_n505));
  INV_X1    g319(.A(G122), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G116), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n334), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n505), .A2(new_n509), .A3(new_n507), .ZN(new_n510));
  OAI21_X1  g324(.A(G107), .B1(new_n505), .B2(new_n509), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n504), .B(new_n508), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n513), .A2(KEYINPUT13), .B1(new_n204), .B2(G128), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n513), .A2(KEYINPUT13), .ZN(new_n515));
  OAI21_X1  g329(.A(G134), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n516), .A2(new_n503), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n503), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n334), .B1(new_n505), .B2(new_n507), .ZN(new_n519));
  INV_X1    g333(.A(new_n508), .ZN(new_n520));
  OAI22_X1  g334(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G217), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n400), .A2(new_n523), .A3(G953), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n512), .A2(new_n521), .A3(new_n524), .ZN(new_n527));
  AOI21_X1  g341(.A(G902), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G478), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n528), .B(new_n530), .Z(new_n531));
  INV_X1    g345(.A(G952), .ZN(new_n532));
  AOI211_X1 g346(.A(G953), .B(new_n532), .C1(G234), .C2(G237), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT21), .B(G898), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(G902), .B(G953), .C1(new_n284), .C2(new_n455), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n499), .A2(new_n502), .A3(new_n531), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT85), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n331), .A2(new_n450), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(new_n342), .ZN(G3));
  NAND2_X1  g356(.A1(new_n499), .A2(new_n502), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT87), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n529), .A2(G902), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT33), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n526), .A2(new_n546), .A3(new_n527), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n526), .B2(new_n527), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n544), .B(new_n545), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n545), .ZN(new_n551));
  INV_X1    g365(.A(new_n549), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(new_n547), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT87), .B1(new_n528), .B2(G478), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n543), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n538), .B(new_n405), .C1(new_n447), .C2(new_n448), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n557), .A2(KEYINPUT88), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n560));
  INV_X1    g374(.A(new_n558), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n555), .B1(new_n499), .B2(new_n502), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n277), .B1(new_n268), .B2(new_n248), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT86), .A2(G472), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  AND4_X1   g381(.A1(new_n330), .A2(new_n399), .A3(new_n403), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(G104), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(G6));
  NOR2_X1   g386(.A1(new_n489), .A2(KEYINPUT20), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT20), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n487), .B2(new_n488), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n531), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n502), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n558), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n568), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G107), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(G9));
  NAND2_X1  g397(.A1(new_n326), .A2(new_n327), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n286), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n286), .A2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n317), .A2(KEYINPUT91), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n322), .A2(KEYINPUT36), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n310), .A2(new_n316), .A3(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n588), .B1(new_n587), .B2(new_n590), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT92), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(new_n586), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n585), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n567), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n450), .A2(new_n540), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT37), .B(G110), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G12));
  NAND3_X1  g417(.A1(new_n281), .A2(new_n283), .A3(new_n597), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n604), .A2(new_n449), .A3(new_n404), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT95), .B(G900), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n606), .A2(new_n537), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n534), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n573), .B2(new_n575), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n578), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G128), .ZN(G30));
  INV_X1    g426(.A(new_n404), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n608), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n616), .A2(KEYINPUT40), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(KEYINPUT40), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n265), .A2(new_n269), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n267), .A2(new_n247), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n247), .A2(new_n253), .A3(new_n254), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n277), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n597), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n405), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n436), .A2(new_n445), .ZN(new_n627));
  INV_X1    g441(.A(new_n446), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n436), .A2(new_n445), .A3(new_n446), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n543), .A2(new_n577), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n626), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n617), .A2(new_n618), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G143), .ZN(G45));
  INV_X1    g451(.A(new_n608), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n638), .B(new_n555), .C1(new_n499), .C2(new_n502), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n605), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G146), .ZN(G48));
  NAND3_X1  g455(.A1(new_n281), .A2(new_n283), .A3(new_n330), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n383), .B1(new_n360), .B2(KEYINPUT75), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n388), .B1(new_n643), .B2(new_n363), .ZN(new_n644));
  OAI21_X1  g458(.A(G469), .B1(new_n644), .B2(G902), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n392), .A2(new_n645), .A3(new_n403), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n564), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT41), .B(G113), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G15));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n579), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G116), .ZN(G18));
  INV_X1    g466(.A(new_n604), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n391), .B1(new_n390), .B2(new_n277), .ZN(new_n654));
  AOI211_X1 g468(.A(G469), .B(G902), .C1(new_n385), .C2(new_n389), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n405), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n629), .B2(new_n630), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n656), .A2(KEYINPUT98), .A3(new_n658), .A4(new_n403), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n660), .B1(new_n646), .B2(new_n449), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n653), .A2(new_n662), .A3(new_n540), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  INV_X1    g479(.A(new_n329), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n585), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT100), .B1(new_n328), .B2(new_n329), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n264), .B1(new_n268), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n260), .A2(new_n258), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n272), .A2(new_n273), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT31), .B1(new_n673), .B2(new_n247), .ZN(new_n674));
  OAI211_X1 g488(.A(KEYINPUT99), .B(new_n672), .C1(new_n674), .C2(new_n260), .ZN(new_n675));
  AOI22_X1  g489(.A1(G472), .A2(new_n565), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n677), .A2(new_n634), .A3(new_n558), .A4(new_n646), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n506), .ZN(G24));
  NAND4_X1  g493(.A1(new_n562), .A2(new_n597), .A3(new_n676), .A4(new_n608), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n392), .A2(new_n645), .A3(new_n403), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT98), .B1(new_n682), .B2(new_n658), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n646), .A2(new_n449), .A3(new_n660), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n662), .A2(KEYINPUT101), .A3(new_n681), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G125), .ZN(G27));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n395), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n395), .A2(new_n691), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(G469), .A3(new_n396), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n392), .A3(new_n394), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n695), .A2(new_n403), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n447), .A2(new_n448), .A3(new_n657), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n639), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n669), .A2(new_n280), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT42), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n403), .A3(new_n697), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n562), .A2(new_n702), .A3(new_n608), .ZN(new_n703));
  OR3_X1    g517(.A1(new_n642), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n704), .A3(KEYINPUT103), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n562), .A2(new_n608), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n699), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n702), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n642), .A2(new_n701), .A3(new_n703), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n706), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n215), .ZN(G33));
  NOR2_X1   g528(.A1(new_n642), .A2(new_n701), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n610), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT104), .B(G134), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G36));
  AND2_X1   g532(.A1(new_n499), .A2(new_n502), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n556), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT105), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n719), .A2(KEYINPUT106), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n543), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n724), .A2(KEYINPUT43), .A3(new_n556), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n720), .A2(new_n728), .A3(new_n721), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n723), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT107), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT107), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n625), .A2(new_n567), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n731), .A2(KEYINPUT44), .A3(new_n732), .A4(new_n733), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n391), .B1(new_n398), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n692), .A2(KEYINPUT45), .A3(new_n396), .A4(new_n693), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n393), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n392), .B1(new_n741), .B2(KEYINPUT46), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n403), .A3(new_n615), .ZN(new_n745));
  INV_X1    g559(.A(new_n697), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n736), .A2(new_n737), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT108), .B(G137), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G39));
  AND2_X1   g564(.A1(new_n281), .A2(new_n283), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n751), .A2(new_n330), .A3(new_n707), .A4(new_n746), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n744), .A2(new_n403), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n744), .A2(KEYINPUT47), .A3(new_n403), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n298), .ZN(G42));
  XOR2_X1   g573(.A(new_n656), .B(KEYINPUT109), .Z(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT49), .Z(new_n761));
  NAND3_X1  g575(.A1(new_n724), .A2(new_n556), .A3(new_n726), .ZN(new_n762));
  INV_X1    g576(.A(new_n624), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n402), .A2(new_n657), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n633), .A2(new_n763), .A3(new_n669), .A4(new_n764), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n761), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n653), .B(new_n450), .C1(new_n610), .C2(new_n639), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n634), .A2(new_n449), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n597), .A2(new_n638), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n696), .A2(new_n769), .A3(new_n624), .A4(new_n770), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n686), .B(new_n680), .C1(new_n661), .C2(new_n659), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT101), .B1(new_n662), .B2(new_n681), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n768), .B(new_n771), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT112), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n689), .A2(new_n776), .A3(new_n768), .A4(new_n771), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n450), .B(new_n540), .C1(new_n331), .C2(new_n598), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n543), .A2(KEYINPUT110), .A3(new_n531), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT110), .B1(new_n543), .B2(new_n531), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n557), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n561), .A3(new_n568), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n651), .A2(new_n663), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n678), .B1(new_n564), .B2(new_n647), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n502), .A2(new_n531), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n609), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n399), .A2(new_n791), .A3(new_n403), .A4(new_n697), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n604), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n604), .B2(new_n792), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n676), .A2(new_n597), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n715), .A2(new_n610), .B1(new_n708), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n789), .A2(new_n713), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n780), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n705), .A2(new_n712), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n677), .A2(new_n634), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n561), .A3(new_n682), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n648), .A2(new_n651), .A3(new_n663), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n781), .A2(new_n785), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n796), .A2(new_n799), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n804), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n778), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n775), .A2(new_n777), .A3(KEYINPUT52), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(KEYINPUT53), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n802), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n814), .A2(new_n803), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n767), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n746), .A2(new_n646), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT116), .B1(new_n730), .B2(new_n533), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n730), .A2(KEYINPUT116), .A3(new_n533), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n709), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT48), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(KEYINPUT48), .A3(new_n709), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n677), .B1(new_n821), .B2(new_n822), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n662), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n330), .A2(new_n763), .A3(new_n818), .A4(new_n533), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n532), .B(G953), .C1(new_n830), .C2(new_n562), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n826), .A2(new_n827), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n719), .A3(new_n555), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT120), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n823), .B2(new_n798), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n760), .A2(KEYINPUT117), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n760), .A2(KEYINPUT117), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n402), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n756), .A3(new_n757), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n828), .A2(new_n839), .A3(new_n697), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n835), .A2(KEYINPUT51), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n633), .A2(new_n657), .A3(new_n682), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n828), .A2(KEYINPUT50), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n677), .ZN(new_n844));
  INV_X1    g658(.A(new_n822), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n844), .B(new_n842), .C1(new_n845), .C2(new_n820), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n832), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n840), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n828), .A2(new_n839), .A3(KEYINPUT118), .A4(new_n697), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n835), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n843), .A2(KEYINPUT119), .A3(new_n848), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT119), .B1(new_n843), .B2(new_n848), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n850), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT53), .B1(new_n812), .B2(new_n813), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n807), .B(KEYINPUT114), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n710), .A2(new_n711), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n810), .A2(new_n786), .A3(new_n863), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n778), .A2(new_n861), .A3(new_n864), .A4(new_n779), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n860), .A2(new_n865), .A3(KEYINPUT54), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n817), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n766), .B1(new_n867), .B2(new_n868), .ZN(G75));
  NOR2_X1   g683(.A1(new_n319), .A2(G952), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n775), .A2(new_n777), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n813), .A3(new_n801), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n861), .A2(new_n864), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n875), .A2(new_n862), .B1(new_n780), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n277), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n878), .B2(G210), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n418), .B1(new_n434), .B2(new_n435), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n432), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n871), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n879), .B2(new_n882), .ZN(G51));
  XNOR2_X1  g698(.A(new_n877), .B(KEYINPUT54), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n393), .B(KEYINPUT57), .Z(new_n886));
  OAI21_X1  g700(.A(new_n390), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n739), .A2(new_n740), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT121), .Z(new_n889));
  NAND2_X1  g703(.A1(new_n878), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n870), .B1(new_n887), .B2(new_n890), .ZN(G54));
  NAND3_X1  g705(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n892));
  INV_X1    g706(.A(new_n487), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n870), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n548), .B2(new_n549), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n871), .B1(new_n885), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n817), .B2(new_n866), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n548), .A2(new_n549), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(G63));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n905));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT122), .B1(new_n877), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n909));
  INV_X1    g723(.A(new_n907), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n909), .B(new_n910), .C1(new_n860), .C2(new_n865), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n325), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n871), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n591), .A2(new_n592), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n908), .B2(new_n911), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n905), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n908), .A2(new_n911), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n914), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n919), .A2(KEYINPUT61), .A3(new_n871), .A4(new_n912), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(G66));
  INV_X1    g735(.A(G224), .ZN(new_n922));
  OAI21_X1  g736(.A(G953), .B1(new_n535), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n809), .B2(G953), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n880), .B1(G898), .B2(new_n319), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(G69));
  AOI21_X1  g740(.A(new_n319), .B1(G227), .B2(G900), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n482), .B(KEYINPUT123), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n266), .B(new_n928), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT124), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n642), .A2(new_n746), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n784), .A2(new_n613), .A3(new_n615), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n758), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n748), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n636), .A2(new_n689), .A3(new_n768), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT62), .Z(new_n937));
  AND2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(KEYINPUT125), .B(new_n931), .C1(new_n938), .C2(G953), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  AOI21_X1  g754(.A(G953), .B1(new_n935), .B2(new_n937), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n930), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n929), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n689), .A2(new_n768), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n709), .A2(new_n769), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n716), .B1(new_n745), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n758), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n748), .A2(new_n804), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n319), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n319), .A2(G900), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT126), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n944), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n927), .B1(new_n943), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n927), .ZN(new_n956));
  AOI211_X1 g770(.A(new_n953), .B(new_n956), .C1(new_n939), .C2(new_n942), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n949), .B2(new_n789), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n267), .A2(new_n247), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n960), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n938), .B2(new_n809), .ZN(new_n966));
  INV_X1    g780(.A(new_n620), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n964), .B(new_n871), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n815), .A2(new_n816), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n963), .A2(new_n620), .A3(new_n965), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT127), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n969), .B2(new_n971), .ZN(G57));
endmodule


