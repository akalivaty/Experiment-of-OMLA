//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(G122), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G110), .ZN(new_n188));
  INV_X1    g002(.A(G110), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G122), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT87), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n188), .B2(new_n190), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT2), .B(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT67), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G116), .ZN(new_n203));
  INV_X1    g017(.A(G116), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n199), .A2(new_n201), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n206), .A2(new_n200), .A3(new_n208), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT2), .B(G113), .Z(new_n210));
  XNOR2_X1  g024(.A(G116), .B(G119), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT68), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n207), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  OAI211_X1 g030(.A(G104), .B(new_n215), .C1(new_n216), .C2(KEYINPUT80), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT81), .A3(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n215), .B2(G104), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(KEYINPUT80), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n224), .A2(new_n225), .B1(G104), .B2(new_n215), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n214), .B(G101), .C1(new_n222), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n218), .A2(G107), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n218), .A2(G107), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n229), .A2(new_n224), .B1(new_n230), .B2(new_n220), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n215), .A2(G104), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n216), .A2(KEYINPUT80), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n231), .A2(new_n235), .A3(new_n236), .A4(new_n219), .ZN(new_n237));
  OAI21_X1  g051(.A(G101), .B1(new_n222), .B2(new_n226), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT4), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT82), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n237), .A2(new_n238), .A3(new_n241), .A4(KEYINPUT4), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n228), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT84), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n230), .B1(new_n229), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n232), .A2(KEYINPUT84), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n237), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n210), .A2(KEYINPUT68), .A3(new_n211), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n208), .B1(new_n206), .B2(new_n200), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT5), .ZN(new_n251));
  INV_X1    g065(.A(new_n203), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT5), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n196), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n249), .A2(new_n250), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n194), .B1(new_n243), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n213), .A2(new_n227), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n222), .A2(new_n226), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n214), .B1(new_n260), .B2(new_n236), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n241), .B1(new_n261), .B2(new_n238), .ZN(new_n262));
  INV_X1    g076(.A(new_n242), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n194), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n256), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n258), .A2(new_n266), .A3(KEYINPUT6), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n268), .B(new_n194), .C1(new_n243), .C2(new_n257), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT88), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G143), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n272), .A2(new_n274), .A3(new_n275), .A4(G128), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT1), .B1(new_n273), .B2(G146), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(G128), .B1(new_n272), .B2(new_n274), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G125), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n270), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(G128), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n272), .A2(new_n274), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(new_n270), .A3(new_n281), .A4(new_n276), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OR2_X1    g103(.A1(KEYINPUT0), .A2(G128), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n272), .A2(new_n274), .A3(new_n287), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n289), .A2(G125), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n282), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G224), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G953), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n294), .B(new_n296), .Z(new_n297));
  NAND3_X1  g111(.A1(new_n267), .A2(new_n269), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n249), .A2(new_n250), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n251), .A2(KEYINPUT90), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n211), .A2(new_n301), .A3(KEYINPUT5), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n302), .A3(new_n254), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n299), .A2(new_n303), .A3(KEYINPUT91), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n248), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT89), .B1(new_n192), .B2(new_n193), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n189), .A2(G122), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n187), .A2(G110), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT87), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT89), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT8), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT8), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n309), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n237), .A2(new_n247), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n317), .A2(new_n319), .B1(new_n320), .B2(new_n255), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT7), .B1(new_n295), .B2(G953), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n282), .B2(new_n293), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n285), .A2(new_n276), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT88), .B1(new_n325), .B2(G125), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n326), .A2(new_n292), .A3(new_n286), .A4(new_n322), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n308), .A2(new_n321), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n266), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G902), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT92), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n332));
  AOI211_X1 g146(.A(new_n332), .B(G902), .C1(new_n266), .C2(new_n328), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n298), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G210), .B1(G237), .B2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n335), .B(new_n298), .C1(new_n331), .C2(new_n333), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(KEYINPUT93), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(G214), .B1(G237), .B2(G902), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n338), .A2(KEYINPUT93), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(KEYINPUT98), .A2(G122), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT98), .A2(G122), .ZN(new_n344));
  OAI21_X1  g158(.A(G116), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n204), .A2(G122), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(KEYINPUT14), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(G107), .ZN(new_n349));
  INV_X1    g163(.A(G134), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n273), .A2(G128), .ZN(new_n351));
  INV_X1    g165(.A(G128), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G143), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT100), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n353), .A3(new_n350), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n357), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT100), .B1(new_n359), .B2(new_n354), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n345), .B(new_n346), .C1(KEYINPUT14), .C2(new_n215), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n349), .A2(new_n358), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT13), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n352), .B2(G143), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n273), .A2(KEYINPUT13), .A3(G128), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n353), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G134), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT99), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n347), .A2(G107), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n215), .B1(new_n345), .B2(new_n346), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n357), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n362), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(new_n375), .A3(G953), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n362), .B(new_n376), .C1(new_n369), .C2(new_n372), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(KEYINPUT101), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT101), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n373), .A2(new_n381), .A3(new_n377), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n330), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT102), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT102), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(new_n385), .A3(new_n330), .A4(new_n382), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT15), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n384), .A2(new_n386), .B1(new_n387), .B2(G478), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n386), .A2(new_n387), .A3(G478), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G952), .ZN(new_n391));
  AOI211_X1 g205(.A(G953), .B(new_n391), .C1(G234), .C2(G237), .ZN(new_n392));
  INV_X1    g206(.A(G953), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n330), .B(new_n393), .C1(G234), .C2(G237), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(G475), .A2(G902), .ZN(new_n398));
  INV_X1    g212(.A(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G125), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n400), .A2(KEYINPUT16), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n281), .A2(G140), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n402), .A3(KEYINPUT16), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(G146), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(G146), .B1(new_n401), .B2(new_n403), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G237), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n393), .A3(G214), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n273), .ZN(new_n411));
  NOR2_X1   g225(.A1(G237), .A2(G953), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n412), .B(G214), .C1(KEYINPUT94), .C2(G143), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT17), .A3(G131), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(G131), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n407), .B(new_n415), .C1(new_n416), .C2(KEYINPUT17), .ZN(new_n417));
  XOR2_X1   g231(.A(G113), .B(G122), .Z(new_n418));
  XOR2_X1   g232(.A(KEYINPUT97), .B(G104), .Z(new_n419));
  XOR2_X1   g233(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT18), .A2(G131), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n414), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n400), .A2(new_n402), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT95), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n400), .A2(new_n402), .A3(KEYINPUT95), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(G146), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT96), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n423), .A2(G146), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n428), .B1(new_n427), .B2(new_n430), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n422), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n417), .A2(new_n420), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n425), .A2(KEYINPUT19), .A3(new_n426), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(new_n271), .C1(KEYINPUT19), .C2(new_n423), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n416), .A2(new_n436), .A3(new_n404), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n420), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n398), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT20), .ZN(new_n440));
  INV_X1    g254(.A(new_n438), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n417), .A2(new_n420), .A3(new_n433), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n398), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n420), .B1(new_n417), .B2(new_n433), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n330), .B1(new_n434), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n440), .A2(new_n445), .B1(G475), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n390), .A2(new_n397), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n342), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n412), .A2(G210), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT27), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT26), .B(G101), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT71), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n299), .A2(new_n207), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n350), .B2(G137), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT11), .ZN(new_n460));
  INV_X1    g274(.A(G131), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT11), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n458), .B(new_n462), .C1(new_n350), .C2(G137), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n350), .A2(G137), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n461), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G137), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(KEYINPUT65), .A3(G134), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n464), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT65), .B1(new_n466), .B2(G134), .ZN(new_n469));
  OAI21_X1  g283(.A(G131), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(KEYINPUT66), .A3(new_n470), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n325), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT64), .B1(new_n466), .B2(G134), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n464), .B1(new_n476), .B2(new_n462), .ZN(new_n477));
  INV_X1    g291(.A(new_n463), .ZN(new_n478));
  OAI21_X1  g292(.A(G131), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n465), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n457), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n291), .A2(new_n290), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n287), .B1(new_n272), .B2(new_n274), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n289), .A2(KEYINPUT69), .A3(new_n290), .A4(new_n291), .ZN(new_n488));
  INV_X1    g302(.A(new_n465), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n459), .A2(KEYINPUT11), .B1(new_n350), .B2(G137), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n461), .B1(new_n490), .B2(new_n463), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n325), .A2(new_n465), .A3(new_n470), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n492), .A2(new_n457), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n456), .B(KEYINPUT28), .C1(new_n483), .C2(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n494), .A2(KEYINPUT28), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n457), .A3(new_n493), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n280), .B1(new_n471), .B2(new_n472), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n499), .A2(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n500), .B2(new_n457), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n456), .B1(new_n501), .B2(KEYINPUT28), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n455), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT72), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT28), .B1(new_n483), .B2(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n496), .A3(new_n495), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT72), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n455), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n492), .B2(new_n493), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n511), .B2(new_n500), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n454), .B(new_n498), .C1(new_n513), .C2(new_n457), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT31), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n492), .A2(new_n493), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT30), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n475), .A2(new_n511), .A3(new_n482), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n457), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n519), .A2(new_n455), .A3(new_n494), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT70), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n523), .A3(KEYINPUT31), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n515), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n510), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G472), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n330), .A3(KEYINPUT73), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT73), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(G472), .B2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n531), .A2(KEYINPUT32), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n494), .A2(KEYINPUT28), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n516), .A2(new_n213), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n498), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(KEYINPUT28), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT29), .A3(new_n454), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n519), .A2(new_n454), .A3(new_n494), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n507), .B2(new_n454), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n330), .B(new_n538), .C1(new_n540), .C2(KEYINPUT29), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G472), .ZN(new_n542));
  INV_X1    g356(.A(new_n531), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n510), .B2(new_n525), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n533), .B(new_n542), .C1(KEYINPUT32), .C2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT24), .B(G110), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT75), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n202), .A2(G128), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n352), .A2(G119), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI22_X1  g366(.A1(new_n547), .A2(new_n552), .B1(new_n405), .B2(new_n406), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n202), .A2(G128), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT23), .B1(new_n555), .B2(KEYINPUT76), .ZN(new_n556));
  NOR2_X1   g370(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n548), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n556), .A2(KEYINPUT77), .A3(new_n548), .A4(new_n558), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(G110), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT78), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n189), .B1(new_n559), .B2(new_n560), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT78), .B1(new_n566), .B2(new_n562), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n554), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n559), .A2(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n547), .A2(new_n552), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n404), .A3(new_n430), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n393), .A2(G221), .A3(G234), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n573), .B(new_n574), .Z(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n563), .A2(new_n564), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n566), .A2(KEYINPUT78), .A3(new_n562), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n553), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n405), .B(new_n429), .C1(new_n569), .C2(new_n570), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n576), .A2(new_n582), .A3(new_n330), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n576), .A2(new_n582), .A3(KEYINPUT25), .A4(new_n330), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n375), .B1(G234), .B2(new_n330), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(G902), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n576), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G221), .ZN(new_n594));
  INV_X1    g408(.A(new_n374), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n330), .ZN(new_n596));
  INV_X1    g410(.A(G469), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n393), .A2(G227), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT79), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G140), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT85), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n248), .B(new_n325), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(KEYINPUT85), .B(KEYINPUT10), .C1(new_n320), .C2(new_n280), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n605), .A2(new_n606), .B1(new_n603), .B2(new_n604), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n240), .A2(new_n242), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n487), .A2(new_n227), .A3(new_n488), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT83), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT83), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n612), .B(new_n609), .C1(new_n240), .C2(new_n242), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n607), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n480), .ZN(new_n615));
  INV_X1    g429(.A(new_n480), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n616), .B(new_n607), .C1(new_n611), .C2(new_n613), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n602), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n248), .A2(new_n325), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n320), .A2(new_n280), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n480), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT12), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g437(.A(KEYINPUT12), .B(new_n480), .C1(new_n619), .C2(new_n620), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n617), .A2(new_n602), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n597), .B(new_n330), .C1(new_n618), .C2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n597), .A2(new_n330), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n617), .A2(new_n602), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT86), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n617), .A2(KEYINPUT86), .A3(new_n602), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n634), .A3(new_n615), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n617), .A2(new_n625), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n601), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(G469), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n596), .B1(new_n630), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n450), .A2(new_n545), .A3(new_n593), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G101), .ZN(G3));
  AOI21_X1  g455(.A(new_n527), .B1(new_n526), .B2(new_n330), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n544), .B1(new_n642), .B2(KEYINPUT103), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n510), .B2(new_n525), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n527), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n596), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n635), .A2(G469), .A3(new_n637), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n627), .A2(new_n629), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n647), .A2(new_n592), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n337), .A2(new_n338), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT104), .B1(new_n653), .B2(new_n340), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n655));
  INV_X1    g469(.A(new_n340), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n655), .B(new_n656), .C1(new_n337), .C2(new_n338), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n440), .A2(new_n445), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n447), .A2(G475), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(G478), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n383), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n378), .A2(KEYINPUT33), .A3(new_n379), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n380), .A2(new_n382), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n665), .B1(new_n666), .B2(KEYINPUT33), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n330), .A2(G478), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n396), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n658), .A2(new_n659), .A3(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n243), .A2(new_n194), .A3(new_n257), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n308), .A2(new_n321), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n324), .A2(new_n327), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n330), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n332), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n329), .A2(KEYINPUT92), .A3(new_n330), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n335), .B1(new_n680), .B2(new_n298), .ZN(new_n681));
  INV_X1    g495(.A(new_n338), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n340), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n655), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n653), .A2(KEYINPUT104), .A3(new_n340), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n671), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT105), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n672), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n652), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G104), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT106), .B(KEYINPUT34), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G6));
  OR2_X1    g506(.A1(new_n388), .A2(new_n389), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n397), .A3(new_n448), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n652), .A2(new_n658), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT35), .B(G107), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NAND2_X1  g512(.A1(new_n450), .A2(new_n639), .ZN(new_n699));
  OAI22_X1  g513(.A1(new_n580), .A2(new_n581), .B1(KEYINPUT36), .B2(new_n577), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n568), .A2(new_n572), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n590), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n589), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n643), .A2(new_n646), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n699), .B1(new_n706), .B2(KEYINPUT107), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n643), .A2(new_n708), .A3(new_n646), .A4(new_n705), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT37), .B(G110), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT108), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n710), .B(new_n712), .ZN(G12));
  NAND2_X1  g527(.A1(new_n545), .A2(new_n639), .ZN(new_n714));
  INV_X1    g528(.A(new_n705), .ZN(new_n715));
  INV_X1    g529(.A(G900), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n392), .B1(new_n394), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n448), .B(new_n718), .C1(new_n388), .C2(new_n389), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n684), .A2(new_n685), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT109), .B1(new_n714), .B2(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n544), .A2(KEYINPUT32), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n526), .A2(new_n532), .B1(new_n541), .B2(G472), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n651), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n693), .A2(new_n705), .A3(new_n448), .A4(new_n718), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n654), .A2(new_n657), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n722), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT110), .B(G128), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G30));
  XOR2_X1   g546(.A(new_n717), .B(KEYINPUT39), .Z(new_n733));
  NAND2_X1  g547(.A1(new_n639), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT40), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n339), .A2(new_n341), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT38), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n738), .A2(new_n656), .A3(new_n705), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n390), .A2(new_n448), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n519), .A2(new_n494), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n455), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n330), .B1(new_n536), .B2(new_n454), .ZN(new_n743));
  OAI21_X1  g557(.A(G472), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n533), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n723), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n736), .A2(new_n739), .A3(new_n740), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G143), .ZN(G45));
  INV_X1    g562(.A(new_n588), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n585), .B2(new_n586), .ZN(new_n750));
  INV_X1    g564(.A(new_n704), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n718), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n670), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n684), .A2(new_n685), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n714), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n271), .ZN(G48));
  OAI21_X1  g570(.A(new_n330), .B1(new_n618), .B2(new_n626), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(G469), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n648), .A3(new_n627), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n592), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n545), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n672), .B2(new_n687), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT41), .B(G113), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G15));
  NAND4_X1  g578(.A1(new_n658), .A2(new_n545), .A3(new_n695), .A4(new_n760), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G116), .ZN(G18));
  AND3_X1   g580(.A1(new_n758), .A2(new_n648), .A3(new_n627), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n449), .A2(new_n715), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n658), .A2(new_n545), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G119), .ZN(G21));
  NOR3_X1   g584(.A1(new_n759), .A2(new_n592), .A3(new_n396), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n537), .A2(new_n454), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n515), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n521), .B2(new_n520), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n531), .B(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n642), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n771), .A2(new_n658), .A3(new_n740), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G122), .ZN(G24));
  NAND3_X1  g594(.A1(new_n684), .A2(new_n767), .A3(new_n685), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n753), .B(new_n776), .C1(new_n645), .C2(new_n527), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n281), .ZN(G27));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n656), .B1(new_n339), .B2(new_n341), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n545), .A2(new_n593), .A3(new_n639), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n670), .A2(new_n717), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n786), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n651), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n592), .B1(new_n723), .B2(new_n724), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n793), .A3(KEYINPUT42), .A4(new_n788), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G131), .ZN(G33));
  NOR2_X1   g610(.A1(new_n787), .A2(new_n719), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n350), .ZN(G36));
  AOI21_X1  g612(.A(KEYINPUT43), .B1(new_n448), .B2(KEYINPUT113), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n669), .A2(new_n448), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n705), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n647), .A2(KEYINPUT44), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n791), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT115), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n635), .A2(new_n637), .ZN(new_n808));
  OAI21_X1  g622(.A(G469), .B1(new_n808), .B2(KEYINPUT45), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n635), .A2(KEYINPUT45), .A3(new_n637), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n629), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT46), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n627), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n648), .B(new_n733), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT112), .ZN(new_n817));
  INV_X1    g631(.A(new_n815), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n627), .A3(new_n813), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n648), .A4(new_n733), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n805), .B(new_n823), .C1(new_n804), .C2(new_n803), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n647), .A2(new_n802), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT44), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n807), .A2(new_n822), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G137), .ZN(G39));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(KEYINPUT47), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(KEYINPUT47), .ZN(new_n831));
  OAI221_X1 g645(.A(new_n648), .B1(new_n830), .B2(new_n831), .C1(new_n814), .C2(new_n815), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n791), .A2(new_n545), .A3(new_n593), .A4(new_n789), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n813), .A2(new_n627), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n596), .B1(new_n834), .B2(new_n818), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n832), .B(new_n833), .C1(new_n835), .C2(new_n831), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  INV_X1    g651(.A(new_n746), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n758), .A2(new_n627), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT49), .Z(new_n840));
  NOR4_X1   g654(.A1(new_n592), .A2(new_n800), .A3(new_n596), .A4(new_n656), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n840), .A3(new_n738), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n778), .A2(new_n801), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n593), .A2(new_n392), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n786), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n835), .A2(new_n831), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n832), .ZN(new_n849));
  INV_X1    g663(.A(new_n839), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n596), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n746), .A2(new_n759), .A3(new_n791), .A4(new_n845), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n662), .A2(new_n669), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n786), .A2(new_n767), .A3(new_n392), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n705), .A3(new_n778), .A4(new_n801), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n656), .A2(new_n846), .A3(new_n738), .A4(new_n767), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT50), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT50), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n843), .B1(new_n852), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n848), .A2(new_n832), .B1(new_n596), .B2(new_n850), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n863), .B(KEYINPUT51), .C1(new_n866), .C2(new_n847), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n846), .A2(new_n658), .A3(new_n767), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT118), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n857), .A2(new_n793), .A3(new_n801), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT48), .ZN(new_n871));
  INV_X1    g685(.A(new_n670), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n391), .B(G953), .C1(new_n853), .C2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n869), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n865), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n448), .B1(new_n388), .B2(new_n389), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n670), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n397), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n342), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n638), .A2(new_n629), .A3(new_n627), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n880), .A2(new_n593), .A3(new_n648), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n643), .A2(new_n879), .A3(new_n881), .A4(new_n646), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n640), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n707), .B2(new_n709), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n779), .A2(new_n765), .A3(new_n769), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n762), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n797), .B1(new_n790), .B2(new_n794), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n693), .A2(new_n752), .A3(new_n662), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n545), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n782), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n792), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n884), .A2(new_n886), .A3(new_n887), .A4(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n684), .A2(new_n685), .A3(new_n753), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n654), .A2(new_n657), .A3(new_n759), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n725), .A2(new_n893), .B1(new_n894), .B2(new_n890), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n717), .B(KEYINPUT117), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n651), .A2(new_n705), .A3(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n746), .A3(new_n658), .A4(new_n740), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n714), .A2(new_n721), .A3(KEYINPUT109), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n728), .B1(new_n725), .B2(new_n727), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n895), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT52), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n730), .A2(new_n903), .A3(new_n895), .A4(new_n898), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n892), .A2(KEYINPUT53), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n902), .A2(new_n904), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n884), .A2(new_n886), .A3(new_n887), .A4(new_n891), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT54), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n875), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n842), .B1(new_n914), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n393), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n330), .B1(new_n905), .B2(new_n909), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n267), .A2(new_n269), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n297), .ZN(new_n922));
  XOR2_X1   g736(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n918), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n910), .B2(G902), .ZN(new_n927));
  AOI211_X1 g741(.A(KEYINPUT120), .B(new_n330), .C1(new_n905), .C2(new_n909), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n336), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n925), .B1(new_n930), .B2(new_n932), .ZN(G51));
  NOR2_X1   g747(.A1(new_n809), .A2(new_n810), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n628), .B(KEYINPUT57), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n912), .A2(new_n913), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n618), .A2(new_n626), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT121), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n917), .B1(new_n935), .B2(new_n940), .ZN(G54));
  AND2_X1   g755(.A1(KEYINPUT58), .A2(G475), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n443), .B1(new_n929), .B2(new_n942), .ZN(new_n943));
  OAI22_X1  g757(.A1(new_n714), .A2(new_n754), .B1(new_n781), .B2(new_n782), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n729), .B2(new_n722), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n903), .B1(new_n945), .B2(new_n898), .ZN(new_n946));
  AND4_X1   g760(.A1(new_n903), .A2(new_n730), .A3(new_n895), .A4(new_n898), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT53), .B1(new_n948), .B2(new_n892), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n907), .A2(new_n908), .A3(new_n906), .ZN(new_n950));
  OAI21_X1  g764(.A(G902), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT120), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n919), .A2(new_n926), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n443), .A2(new_n942), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n918), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n943), .A2(new_n956), .ZN(G60));
  XNOR2_X1  g771(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n663), .A2(new_n330), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n912), .A2(new_n913), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n667), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n918), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n667), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT60), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n910), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n576), .A2(new_n582), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT123), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT124), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n967), .B1(new_n905), .B2(new_n909), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n917), .B1(new_n974), .B2(new_n703), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n969), .A2(new_n976), .A3(new_n971), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n973), .A2(KEYINPUT61), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n972), .A2(new_n975), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(G66));
  NOR3_X1   g796(.A1(new_n395), .A2(new_n295), .A3(new_n393), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n884), .A2(new_n886), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n393), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n921), .B1(G898), .B2(new_n393), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G69));
  AND3_X1   g801(.A1(new_n836), .A2(new_n887), .A3(new_n945), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n822), .A2(new_n793), .A3(new_n658), .A4(new_n740), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n988), .A2(new_n827), .A3(new_n393), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n425), .A2(new_n426), .ZN(new_n991));
  MUX2_X1   g805(.A(new_n423), .B(new_n991), .S(KEYINPUT19), .Z(new_n992));
  XOR2_X1   g806(.A(new_n513), .B(new_n992), .Z(new_n993));
  OAI211_X1 g807(.A(new_n990), .B(new_n993), .C1(new_n716), .C2(new_n393), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n747), .A2(new_n945), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT62), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n545), .A2(new_n593), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n877), .B(new_n999), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n998), .A2(new_n734), .A3(new_n1000), .A4(new_n791), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n836), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n997), .A2(new_n827), .A3(new_n1004), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n1005), .A2(new_n393), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n994), .B1(new_n1006), .B2(new_n993), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n393), .B1(G227), .B2(G900), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1008), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n994), .B(new_n1010), .C1(new_n1006), .C2(new_n993), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(G72));
  NAND4_X1  g826(.A1(new_n997), .A2(new_n827), .A3(new_n1004), .A4(new_n984), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n917), .B1(new_n1016), .B2(new_n742), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n988), .A2(new_n827), .A3(new_n984), .A4(new_n989), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n1015), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n539), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1021));
  INV_X1    g835(.A(new_n539), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n1015), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1023), .A2(new_n742), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1021), .B1(new_n910), .B2(new_n1024), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n910), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1017), .B(new_n1020), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(G57));
endmodule


