//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT88), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G8gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(G1gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n204), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT14), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT15), .A3(new_n209), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n210), .A2(new_n214), .A3(new_n218), .A4(new_n215), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(KEYINPUT17), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n219), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n208), .B(new_n220), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n204), .B(new_n207), .Z(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n221), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT18), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n222), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n227), .B(KEYINPUT13), .Z(new_n232));
  AOI22_X1  g031(.A1(new_n228), .A2(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n224), .A2(new_n226), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n227), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G113gat), .B(G141gat), .Z(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT11), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G169gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G197gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT12), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n233), .A3(new_n235), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(KEYINPUT89), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT89), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n236), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT29), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  NAND2_X1  g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(KEYINPUT23), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n254), .A2(G169gat), .A3(G176gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT24), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n257), .A2(G183gat), .A3(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(G183gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G190gat), .ZN(new_n260));
  INV_X1    g059(.A(G190gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G183gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n263), .B2(KEYINPUT24), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n252), .A2(KEYINPUT23), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n254), .B1(G169gat), .B2(G176gat), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n265), .A2(KEYINPUT65), .A3(new_n266), .A4(new_n251), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n269));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n255), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n257), .B1(new_n260), .B2(new_n262), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n271), .A2(new_n272), .A3(new_n258), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n268), .A2(new_n269), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT27), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT27), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G183gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n277), .A3(new_n261), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT28), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT27), .B(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(new_n261), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n251), .ZN(new_n285));
  NOR3_X1   g084(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n286));
  OAI22_X1  g085(.A1(new_n285), .A2(new_n286), .B1(new_n259), .B2(new_n261), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n289));
  OAI221_X1 g088(.A(new_n289), .B1(new_n259), .B2(new_n261), .C1(new_n285), .C2(new_n286), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n283), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n249), .B1(new_n274), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G226gat), .ZN(new_n293));
  INV_X1    g092(.A(G233gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n295), .B1(new_n274), .B2(new_n291), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  INV_X1    g098(.A(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n299), .B1(KEYINPUT22), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n304), .B(new_n299), .C1(KEYINPUT22), .C2(new_n302), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n297), .A2(new_n298), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G64gat), .B(G92gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(G36gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT70), .B(G8gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n316), .B(new_n295), .C1(new_n274), .C2(new_n291), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n315), .A2(new_n317), .B1(new_n296), .B2(new_n292), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n309), .B(new_n314), .C1(new_n318), .C2(new_n308), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT30), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT76), .B(KEYINPUT0), .Z(new_n323));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G57gat), .B(G85gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n329));
  INV_X1    g128(.A(G113gat), .ZN(new_n330));
  INV_X1    g129(.A(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  NAND2_X1  g132(.A1(G113gat), .A2(G120gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n336));
  INV_X1    g135(.A(G127gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G134gat), .ZN(new_n338));
  INV_X1    g137(.A(G134gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G127gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n336), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT67), .B1(new_n337), .B2(G134gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G141gat), .B(G148gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(G155gat), .B2(G162gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n346), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G148gat), .ZN(new_n352));
  INV_X1    g151(.A(G148gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G141gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G155gat), .B(G162gat), .ZN(new_n356));
  INV_X1    g155(.A(G155gat), .ZN(new_n357));
  INV_X1    g156(.A(G162gat), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT2), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G127gat), .B(G134gat), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n361), .A2(new_n333), .A3(new_n334), .A4(new_n332), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n343), .A2(new_n350), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n329), .B1(new_n363), .B2(KEYINPUT4), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n338), .A2(new_n340), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n335), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n342), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n361), .B2(new_n336), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n335), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n350), .A2(new_n360), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT74), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n363), .A2(KEYINPUT4), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n364), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n350), .A2(new_n360), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT73), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n350), .A2(new_n360), .A3(KEYINPUT73), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(KEYINPUT3), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n342), .B1(new_n365), .B2(KEYINPUT67), .ZN(new_n382));
  INV_X1    g181(.A(new_n335), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n362), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n350), .A2(new_n360), .A3(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n376), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n374), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT5), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n363), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n392), .B2(new_n376), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n389), .A2(new_n393), .A3(KEYINPUT75), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT75), .B1(new_n389), .B2(new_n393), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI211_X1 g195(.A(KEYINPUT5), .B(new_n376), .C1(new_n381), .C2(new_n387), .ZN(new_n397));
  OR3_X1    g196(.A1(new_n363), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n369), .A2(new_n371), .A3(new_n370), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n373), .A2(new_n399), .A3(KEYINPUT77), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n397), .A2(KEYINPUT78), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n398), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n350), .A2(new_n360), .A3(KEYINPUT73), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT73), .B1(new_n350), .B2(new_n360), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n404), .A2(new_n405), .A3(new_n385), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n386), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n390), .B(new_n375), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n328), .B1(new_n396), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n401), .A2(new_n409), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(new_n327), .C1(new_n395), .C2(new_n394), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n395), .B2(new_n394), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n328), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n322), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT72), .ZN(new_n419));
  INV_X1    g218(.A(new_n319), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n315), .A2(new_n317), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n308), .B1(new_n421), .B2(new_n297), .ZN(new_n422));
  INV_X1    g221(.A(new_n309), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n313), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  AOI22_X1  g224(.A1(KEYINPUT30), .A2(new_n420), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT71), .B(new_n313), .C1(new_n422), .C2(new_n423), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n419), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n425), .ZN(new_n429));
  INV_X1    g228(.A(new_n422), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n430), .A2(KEYINPUT30), .A3(new_n309), .A4(new_n314), .ZN(new_n431));
  AND4_X1   g230(.A1(new_n419), .A2(new_n429), .A3(new_n427), .A4(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n418), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT79), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n426), .A2(new_n419), .A3(new_n427), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n427), .A3(new_n431), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT72), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n418), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT31), .B(G50gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT29), .B1(new_n306), .B2(new_n307), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n377), .B1(new_n443), .B2(KEYINPUT3), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n308), .B1(new_n249), .B2(new_n386), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n386), .A2(new_n249), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n306), .A3(new_n307), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n442), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n453), .B(new_n442), .C1(new_n446), .C2(new_n450), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n445), .A2(new_n442), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n379), .B(new_n380), .C1(new_n443), .C2(KEYINPUT3), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n441), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G78gat), .B(G106gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(G22gat), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n459), .B1(new_n452), .B2(new_n454), .ZN(new_n463));
  INV_X1    g262(.A(new_n441), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n462), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n463), .A2(new_n464), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n441), .B(new_n459), .C1(new_n452), .C2(new_n454), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT68), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n268), .A2(new_n269), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n273), .A2(new_n270), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n288), .A2(new_n290), .ZN(new_n476));
  INV_X1    g275(.A(new_n283), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n369), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n384), .B1(new_n274), .B2(new_n291), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G227gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n294), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n472), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n483), .ZN(new_n485));
  AOI211_X1 g284(.A(KEYINPUT68), .B(new_n485), .C1(new_n479), .C2(new_n480), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT32), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT33), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n484), .B2(new_n486), .ZN(new_n489));
  XOR2_X1   g288(.A(G15gat), .B(G43gat), .Z(new_n490));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n487), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n479), .A2(new_n480), .A3(new_n485), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(KEYINPUT34), .Z(new_n495));
  INV_X1    g294(.A(new_n492), .ZN(new_n496));
  OAI221_X1 g295(.A(KEYINPUT32), .B1(new_n488), .B2(new_n496), .C1(new_n484), .C2(new_n486), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n497), .ZN(new_n499));
  INV_X1    g298(.A(new_n495), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n471), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n498), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n495), .B1(new_n493), .B2(new_n497), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(KEYINPUT86), .A3(new_n471), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n434), .A2(new_n440), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n511), .A3(new_n471), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n417), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n416), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n328), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n415), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n429), .A2(new_n431), .A3(new_n427), .A4(new_n321), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT85), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n512), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n434), .A2(new_n440), .ZN(new_n526));
  INV_X1    g325(.A(new_n471), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT37), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n430), .B2(new_n309), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n529), .B(new_n309), .C1(new_n318), .C2(new_n308), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n313), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT38), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT38), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n318), .B1(new_n306), .B2(new_n307), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n297), .A2(new_n298), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT37), .B1(new_n536), .B2(new_n308), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n534), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n533), .B(new_n319), .C1(new_n532), .C2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n471), .B1(new_n539), .B2(new_n516), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n389), .A2(new_n393), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n389), .A2(new_n393), .A3(KEYINPUT75), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n543), .A2(new_n544), .B1(new_n409), .B2(new_n401), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n381), .A2(new_n387), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n400), .A2(new_n398), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT39), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n376), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n547), .A2(new_n376), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT39), .B1(new_n392), .B2(new_n376), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n327), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT40), .ZN(new_n553));
  OAI22_X1  g352(.A1(new_n545), .A2(new_n327), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT82), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT82), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(new_n557), .A3(new_n553), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT83), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n559), .A2(new_n560), .A3(new_n517), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n560), .B1(new_n559), .B2(new_n517), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n540), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n505), .B2(new_n506), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n501), .A2(KEYINPUT36), .A3(new_n498), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n528), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n248), .B1(new_n525), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n572));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT7), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G99gat), .B(G106gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n220), .B(new_n585), .C1(new_n222), .C2(new_n223), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n221), .A2(new_n584), .B1(KEYINPUT41), .B2(new_n571), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n586), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n575), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n592), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(new_n574), .A3(new_n590), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(KEYINPUT90), .A2(G57gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(G64gat), .Z(new_n598));
  AND2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(KEYINPUT9), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(G57gat), .B2(G64gat), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n604), .A2(new_n599), .A3(new_n600), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n208), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G183gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n609), .B(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n614));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G211gat), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n617), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n596), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n584), .A2(new_n606), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n584), .A2(new_n606), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(KEYINPUT92), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G204gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT93), .B(G176gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n621), .A2(new_n633), .A3(new_n622), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT91), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n584), .A2(new_n635), .A3(KEYINPUT10), .A4(new_n606), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT91), .B1(new_n622), .B2(new_n633), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n624), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n626), .A2(KEYINPUT92), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n626), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n631), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n620), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n570), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n415), .A2(new_n417), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(KEYINPUT94), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n649), .A2(KEYINPUT94), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n648), .A2(new_n517), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT16), .B(G8gat), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n658), .A2(new_n659), .B1(G8gat), .B2(new_n656), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n656), .A2(new_n659), .A3(new_n657), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n505), .A2(new_n565), .A3(new_n506), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT36), .B1(new_n501), .B2(new_n498), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT96), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n647), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n507), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(G15gat), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n647), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT98), .ZN(G1326gat));
  OR3_X1    g477(.A1(new_n647), .A2(KEYINPUT99), .A3(new_n471), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT99), .B1(new_n647), .B2(new_n471), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT43), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n679), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G22gat), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n618), .A2(new_n619), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n644), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n596), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n570), .A2(new_n211), .A3(new_n653), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT45), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n471), .B1(new_n434), .B2(new_n440), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(new_n563), .A3(new_n671), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n523), .B1(new_n509), .B2(KEYINPUT35), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n596), .B(new_n693), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n596), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n525), .B2(new_n569), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n245), .A2(new_n247), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n688), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT100), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n653), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n707), .ZN(G1328gat));
  OAI21_X1  g507(.A(G36gat), .B1(new_n705), .B2(new_n518), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n570), .A2(new_n212), .A3(new_n517), .A4(new_n690), .ZN(new_n710));
  AND2_X1   g509(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n709), .B(new_n713), .C1(new_n711), .C2(new_n710), .ZN(G1329gat));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  AND4_X1   g514(.A1(new_n715), .A2(new_n570), .A3(new_n507), .A4(new_n690), .ZN(new_n716));
  INV_X1    g515(.A(new_n705), .ZN(new_n717));
  INV_X1    g516(.A(new_n673), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(G43gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n715), .B1(new_n717), .B2(new_n671), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n720), .A2(KEYINPUT47), .B1(new_n721), .B2(new_n723), .ZN(G1330gat));
  XNOR2_X1  g523(.A(KEYINPUT103), .B(KEYINPUT48), .ZN(new_n725));
  OAI21_X1  g524(.A(G50gat), .B1(new_n705), .B2(new_n471), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n471), .A2(G50gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n570), .A2(new_n690), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n726), .A2(new_n727), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n725), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n726), .A2(KEYINPUT48), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1331gat));
  NAND2_X1  g534(.A1(new_n620), .A2(new_n248), .ZN(new_n736));
  INV_X1    g535(.A(new_n671), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n528), .A2(new_n564), .A3(new_n737), .ZN(new_n738));
  AOI211_X1 g537(.A(new_n645), .B(new_n736), .C1(new_n525), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n653), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT105), .B(G57gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1332gat));
  XOR2_X1   g541(.A(new_n517), .B(KEYINPUT106), .Z(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT107), .Z(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  NAND2_X1  g547(.A1(new_n739), .A2(new_n718), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n675), .A2(G71gat), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n749), .A2(G71gat), .B1(new_n739), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n739), .A2(new_n527), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n702), .A2(new_n687), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n644), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n701), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n706), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n698), .B1(new_n525), .B2(new_n738), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n755), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n596), .B(new_n755), .C1(new_n695), .C2(new_n696), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n644), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n653), .A2(new_n579), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n759), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n743), .A2(G92gat), .A3(new_n645), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n760), .B2(new_n755), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n762), .A2(new_n763), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n701), .A2(new_n517), .A3(new_n757), .ZN(new_n775));
  AOI22_X1  g574(.A1(KEYINPUT109), .A2(new_n774), .B1(new_n775), .B2(G92gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n762), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n761), .B1(new_n777), .B2(new_n771), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n779), .A3(new_n770), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n769), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(G92gat), .B1(new_n758), .B2(new_n743), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n770), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT111), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n775), .A2(G92gat), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(new_n780), .A3(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n788), .B(new_n785), .C1(new_n791), .C2(new_n769), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(new_n792), .ZN(G1337gat));
  INV_X1    g592(.A(G99gat), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n758), .A2(new_n794), .A3(new_n673), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n765), .A2(new_n507), .A3(new_n644), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(G1338gat));
  OAI21_X1  g596(.A(G106gat), .B1(new_n758), .B2(new_n471), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n471), .A2(G106gat), .A3(new_n645), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n765), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n778), .A2(new_n799), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n803), .A2(KEYINPUT112), .A3(KEYINPUT53), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT112), .B1(new_n803), .B2(KEYINPUT53), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(G1339gat));
  NOR2_X1   g605(.A1(new_n234), .A2(new_n227), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n231), .A2(new_n232), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n240), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n644), .A2(new_n244), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n634), .A2(new_n636), .A3(new_n625), .A4(new_n637), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n639), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n638), .A2(new_n624), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n631), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n631), .A4(new_n814), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n641), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n810), .B1(new_n248), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n698), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n596), .A2(new_n244), .A3(new_n809), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT114), .B1(new_n823), .B2(new_n819), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n632), .A2(new_n639), .A3(new_n640), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n815), .B2(new_n816), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n822), .A2(new_n826), .A3(new_n827), .A4(new_n818), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n687), .B1(new_n821), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n736), .A2(new_n644), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT115), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833));
  INV_X1    g632(.A(new_n831), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n820), .A2(new_n698), .B1(new_n824), .B2(new_n828), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n687), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n706), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n504), .A2(new_n508), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(new_n743), .ZN(new_n840));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n702), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n837), .A2(new_n527), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(new_n653), .A3(new_n507), .A4(new_n743), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n330), .A3(new_n248), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n841), .A2(new_n844), .ZN(G1340gat));
  AOI21_X1  g644(.A(G120gat), .B1(new_n840), .B2(new_n644), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n843), .A2(new_n331), .A3(new_n645), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(G1341gat));
  NAND3_X1  g647(.A1(new_n840), .A2(new_n337), .A3(new_n687), .ZN(new_n849));
  INV_X1    g648(.A(new_n687), .ZN(new_n850));
  OAI21_X1  g649(.A(G127gat), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(G1342gat));
  NOR2_X1   g651(.A1(new_n517), .A2(new_n698), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n339), .A3(new_n839), .A4(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n843), .B2(new_n698), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  NAND3_X1  g657(.A1(new_n832), .A2(new_n527), .A3(new_n836), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n826), .A2(new_n864), .A3(new_n818), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n702), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n596), .B1(new_n866), .B2(new_n810), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n824), .A2(new_n828), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n850), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n834), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n471), .A2(new_n860), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT118), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  INV_X1    g672(.A(new_n871), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n873), .B(new_n874), .C1(new_n869), .C2(new_n834), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n877), .A3(new_n860), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n743), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n706), .A2(new_n671), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n702), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n718), .A2(new_n471), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n838), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n887), .A2(new_n351), .A3(new_n702), .A4(new_n743), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n885), .A2(new_n889), .A3(KEYINPUT58), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n883), .B(new_n888), .C1(new_n884), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1344gat));
  NAND2_X1  g692(.A1(new_n879), .A2(new_n881), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n645), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(KEYINPUT59), .A3(new_n353), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  INV_X1    g696(.A(new_n819), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n867), .B1(new_n898), .B2(new_n822), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n834), .B1(new_n899), .B2(new_n687), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n471), .A2(KEYINPUT57), .ZN(new_n901));
  AOI22_X1  g700(.A1(KEYINPUT57), .A2(new_n859), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n644), .A3(new_n881), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n897), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  AND4_X1   g703(.A1(new_n353), .A2(new_n887), .A3(new_n644), .A4(new_n743), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n896), .A2(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1345gat));
  OAI21_X1  g707(.A(G155gat), .B1(new_n894), .B2(new_n850), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n887), .A2(new_n357), .A3(new_n687), .A4(new_n743), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(KEYINPUT121), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n894), .B2(new_n698), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n887), .A2(new_n358), .A3(new_n853), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1347gat));
  NAND4_X1  g717(.A1(new_n842), .A2(new_n706), .A3(new_n507), .A4(new_n517), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n248), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT123), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n837), .A2(new_n653), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n839), .A2(new_n880), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT122), .Z(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n248), .A2(G169gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(G1348gat));
  OAI21_X1  g726(.A(G176gat), .B1(new_n919), .B2(new_n645), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n645), .A2(G176gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n925), .B2(new_n929), .ZN(G1349gat));
  OAI21_X1  g729(.A(G183gat), .B1(new_n919), .B2(new_n850), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n687), .A2(new_n280), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g733(.A(G190gat), .B1(new_n919), .B2(new_n698), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(KEYINPUT124), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n596), .A2(new_n261), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n939));
  OAI221_X1 g738(.A(new_n937), .B1(new_n925), .B2(new_n938), .C1(new_n935), .C2(new_n939), .ZN(G1351gat));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n886), .A3(new_n880), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n702), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n718), .A2(new_n653), .A3(new_n518), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n902), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n702), .A2(G197gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  XNOR2_X1  g747(.A(KEYINPUT125), .B(G204gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n941), .A2(new_n645), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n902), .A2(new_n644), .A3(new_n944), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n949), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n950), .A2(new_n951), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(G1353gat));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n300), .B1(KEYINPUT126), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n945), .B2(new_n850), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n957), .A2(KEYINPUT126), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n942), .A2(new_n300), .A3(new_n687), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(G1354gat));
  NOR3_X1   g763(.A1(new_n945), .A2(new_n301), .A3(new_n698), .ZN(new_n965));
  AOI21_X1  g764(.A(G218gat), .B1(new_n942), .B2(new_n596), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G1355gat));
endmodule


