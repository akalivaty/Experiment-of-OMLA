//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n566, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  MUX2_X1   g039(.A(new_n463), .B(new_n464), .S(G2105), .Z(G160));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G136), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n466), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n469), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT66), .ZN(G162));
  OAI211_X1 g053(.A(G138), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT67), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n462), .A2(new_n482), .A3(G138), .A4(new_n466), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n481), .A2(KEYINPUT4), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(G126), .B1(new_n470), .B2(new_n471), .ZN(new_n485));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n466), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G102), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  OAI211_X1 g068(.A(KEYINPUT67), .B(new_n493), .C1(new_n479), .C2(new_n480), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n484), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G543), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n497), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n500), .A2(new_n506), .ZN(G303));
  INV_X1    g082(.A(G303), .ZN(G166));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n497), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G89), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n497), .A2(G63), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT71), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n518), .A2(new_n520), .A3(G543), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT70), .B(G51), .ZN(new_n522));
  AOI211_X1 g097(.A(new_n514), .B(new_n517), .C1(new_n521), .C2(new_n522), .ZN(G168));
  NAND2_X1  g098(.A1(new_n521), .A2(G52), .ZN(new_n524));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n497), .ZN(new_n526));
  INV_X1    g101(.A(G64), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n528), .A2(G651), .B1(new_n511), .B2(G90), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  AOI22_X1  g106(.A1(new_n497), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n499), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT72), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n510), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n518), .A2(new_n520), .A3(G543), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n533), .A2(KEYINPUT72), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  NAND2_X1  g121(.A1(G78), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n526), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n499), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n551), .B1(new_n550), .B2(new_n549), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n511), .A2(G91), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n521), .A2(KEYINPUT9), .A3(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n537), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n555), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n559), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(KEYINPUT73), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G299));
  XNOR2_X1  g140(.A(G168), .B(KEYINPUT75), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G286));
  AND2_X1   g142(.A1(new_n521), .A2(G49), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n510), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G288));
  AND2_X1   g148(.A1(G48), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n509), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n510), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n497), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n499), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT76), .Z(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n499), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n585), .A2(new_n586), .B1(G85), .B2(new_n511), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n521), .A2(G47), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n587), .B(new_n588), .C1(new_n586), .C2(new_n585), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n526), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n499), .B1(new_n594), .B2(KEYINPUT79), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(KEYINPUT79), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n521), .A2(G54), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n497), .A2(new_n509), .A3(G92), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G284));
  XNOR2_X1  g178(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NOR2_X1   g179(.A1(G299), .A2(G868), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n566), .ZN(G297));
  AOI21_X1  g181(.A(new_n605), .B1(G868), .B2(new_n566), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n602), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n602), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n468), .A2(G135), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT83), .Z(new_n615));
  OR2_X1    g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(G111), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n488), .B1(new_n617), .B2(G2105), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n473), .A2(G123), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n462), .A2(new_n489), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT82), .B(G2100), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n620), .A2(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n627), .C1(new_n621), .C2(new_n620), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT84), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT85), .ZN(new_n631));
  AND2_X1   g206(.A1(new_n631), .A2(G2438), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(G2438), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT86), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n632), .B2(new_n633), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT14), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n643), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(KEYINPUT87), .B1(new_n646), .B2(new_n647), .ZN(new_n649));
  OAI211_X1 g224(.A(KEYINPUT87), .B(new_n647), .C1(new_n644), .C2(new_n645), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(G14), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(KEYINPUT17), .ZN(new_n660));
  INV_X1    g235(.A(new_n654), .ZN(new_n661));
  INV_X1    g236(.A(new_n655), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n657), .A3(new_n662), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(new_n656), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n659), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT88), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT89), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n680), .C1(new_n671), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  INV_X1    g257(.A(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT90), .B(G1986), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n691), .A3(new_n689), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G6), .A2(G16), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n582), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT32), .B(G1981), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G23), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n572), .B2(new_n700), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT33), .Z(new_n703));
  AOI21_X1  g278(.A(new_n699), .B1(G1976), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n700), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT95), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n704), .B(new_n708), .C1(G1976), .C2(new_n703), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT34), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(new_n466), .B2(G107), .ZN(new_n713));
  INV_X1    g288(.A(G95), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n466), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT92), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G119), .B2(new_n473), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n468), .A2(G131), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n712), .B1(new_n721), .B2(new_n711), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G24), .B(G290), .S(G16), .Z(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT93), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n725), .B1(new_n728), .B2(KEYINPUT94), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(KEYINPUT94), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n710), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT36), .Z(new_n732));
  INV_X1    g307(.A(KEYINPUT99), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n473), .A2(G129), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(KEYINPUT98), .B1(new_n489), .B2(G105), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n489), .A2(KEYINPUT98), .A3(G105), .ZN(new_n737));
  INV_X1    g312(.A(G141), .ZN(new_n738));
  OAI22_X1  g313(.A1(new_n736), .A2(new_n737), .B1(new_n467), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT26), .ZN(new_n741));
  OR4_X1    g316(.A1(new_n733), .A2(new_n735), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n735), .A2(new_n741), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n733), .B1(new_n743), .B2(new_n739), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(KEYINPUT100), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n744), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT100), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n711), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT101), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G29), .B2(G32), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n700), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n700), .A2(G5), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G171), .B2(new_n700), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1961), .ZN(new_n762));
  NOR2_X1   g337(.A1(G168), .A2(new_n700), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n700), .B2(G21), .ZN(new_n764));
  INV_X1    g339(.A(G1966), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n711), .A2(G33), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n767));
  NAND2_X1  g342(.A1(G103), .A2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(G2105), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n468), .A2(G139), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n462), .A2(G127), .ZN(new_n773));
  NAND2_X1  g348(.A1(G115), .A2(G2104), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n466), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n771), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n772), .B2(new_n775), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n766), .B1(new_n777), .B2(new_n711), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n764), .A2(new_n765), .B1(G2072), .B2(new_n778), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n762), .B(new_n779), .C1(G2072), .C2(new_n778), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n700), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n541), .B2(new_n700), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n764), .A2(new_n765), .B1(G1341), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n780), .B(new_n783), .C1(G1341), .C2(new_n782), .ZN(new_n784));
  NOR2_X1   g359(.A1(G4), .A2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  INV_X1    g361(.A(new_n602), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n700), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1348), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n711), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n711), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G2078), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n793), .A2(G28), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n711), .B1(new_n793), .B2(G28), .ZN(new_n795));
  AND2_X1   g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  NOR2_X1   g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n620), .B2(G29), .ZN(new_n799));
  AND2_X1   g374(.A1(KEYINPUT24), .A2(G34), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n711), .B1(KEYINPUT24), .B2(G34), .ZN(new_n801));
  OAI22_X1  g376(.A1(G160), .A2(new_n711), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G2084), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(G2084), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n799), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n791), .A2(G2078), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n711), .A2(G26), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT28), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n468), .A2(G140), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n473), .A2(G128), .ZN(new_n810));
  NOR2_X1   g385(.A1(G104), .A2(G2105), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n808), .B1(new_n813), .B2(G29), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G2067), .Z(new_n815));
  NOR3_X1   g390(.A1(new_n805), .A2(new_n806), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n789), .A2(new_n792), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(G29), .A2(G35), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G162), .B2(G29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT29), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2090), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n784), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n732), .A2(new_n755), .A3(new_n759), .A4(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n526), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n827), .A2(KEYINPUT102), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(KEYINPUT102), .ZN(new_n829));
  OR3_X1    g404(.A1(new_n828), .A2(new_n829), .A3(new_n499), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n511), .A2(G93), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT103), .B(G55), .Z(new_n832));
  OAI211_X1 g407(.A(new_n830), .B(new_n831), .C1(new_n537), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n540), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n602), .A2(G559), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n833), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n620), .B(G160), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n747), .B(KEYINPUT107), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n487), .B2(new_n491), .ZN(new_n850));
  INV_X1    g425(.A(new_n486), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n462), .B2(G126), .ZN(new_n852));
  OAI211_X1 g427(.A(KEYINPUT105), .B(new_n490), .C1(new_n852), .C2(new_n466), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n484), .A2(new_n850), .A3(new_n853), .A4(new_n494), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n813), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n777), .B1(new_n848), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n848), .ZN(new_n857));
  INV_X1    g432(.A(new_n855), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n750), .B(new_n858), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n859), .A2(KEYINPUT106), .A3(new_n777), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT106), .B1(new_n859), .B2(new_n777), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n468), .A2(G142), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n473), .A2(G130), .ZN(new_n864));
  OR2_X1    g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n720), .B(new_n623), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n867), .B(new_n857), .C1(new_n860), .C2(new_n861), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n847), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n869), .A2(new_n871), .ZN(new_n876));
  INV_X1    g451(.A(new_n870), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n846), .A3(new_n872), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  NOR3_X1   g457(.A1(new_n563), .A2(new_n554), .A3(new_n560), .ZN(new_n883));
  INV_X1    g458(.A(new_n600), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT41), .ZN(new_n886));
  INV_X1    g461(.A(new_n610), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n834), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n885), .B2(new_n888), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n582), .B(G290), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n572), .B(G166), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n891), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(G868), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n833), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(G868), .B2(new_n899), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  XNOR2_X1  g476(.A(G331), .B(new_n901), .ZN(G295));
  INV_X1    g477(.A(new_n886), .ZN(new_n903));
  NOR2_X1   g478(.A1(G168), .A2(G171), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(new_n566), .B2(G171), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n834), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n885), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n910), .B2(new_n894), .ZN(new_n911));
  INV_X1    g486(.A(new_n894), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n907), .B2(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(new_n909), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n907), .B2(KEYINPUT109), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n907), .A2(KEYINPUT109), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n911), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n922), .A2(KEYINPUT110), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT110), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n919), .B2(new_n911), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT44), .B1(new_n914), .B2(KEYINPUT43), .ZN(new_n927));
  OAI22_X1  g502(.A1(new_n924), .A2(new_n925), .B1(new_n926), .B2(new_n927), .ZN(G397));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT45), .B1(new_n854), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G160), .A2(G40), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G1996), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT111), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(KEYINPUT46), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT124), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n813), .B(G2067), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n747), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n936), .A2(KEYINPUT46), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT47), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n939), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT112), .Z(new_n945));
  NOR2_X1   g520(.A1(new_n745), .A2(new_n934), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n933), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n720), .B(new_n724), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n933), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n936), .A2(new_n749), .A3(new_n746), .ZN(new_n950));
  NOR2_X1   g525(.A1(G290), .A2(G1986), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n933), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT48), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n947), .A2(new_n949), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  AND4_X1   g529(.A1(new_n723), .A2(new_n947), .A3(new_n721), .A4(new_n950), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n813), .A2(G2067), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n933), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n943), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n854), .A2(new_n929), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT114), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n854), .A2(new_n962), .A3(new_n929), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G2090), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n495), .A2(new_n929), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n931), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n854), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n932), .ZN(new_n972));
  INV_X1    g547(.A(G1971), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(G8), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(G8), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n960), .A2(new_n932), .A3(new_n963), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n572), .A2(G1976), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(G8), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n572), .B2(G1976), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(KEYINPUT52), .B2(new_n983), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT115), .A4(new_n683), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n579), .A2(new_n499), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT115), .B(G1981), .C1(new_n989), .C2(new_n577), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(KEYINPUT49), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT49), .B1(new_n988), .B2(new_n990), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n981), .A2(new_n994), .A3(G8), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT116), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n980), .A2(new_n987), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n578), .A2(new_n580), .A3(new_n683), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT117), .ZN(new_n999));
  NOR2_X1   g574(.A1(G288), .A2(G1976), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n981), .A2(G8), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n997), .B(KEYINPUT118), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT63), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n961), .B1(new_n960), .B2(new_n963), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n932), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1010), .A2(new_n965), .B1(new_n973), .B2(new_n972), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n977), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(new_n979), .A3(new_n987), .A4(new_n996), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n854), .A2(new_n962), .A3(new_n929), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n962), .B1(new_n854), .B2(new_n929), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n969), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n932), .B1(new_n966), .B2(new_n969), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n765), .ZN(new_n1021));
  INV_X1    g596(.A(G2084), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n964), .A2(new_n1022), .A3(new_n967), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(G8), .A3(new_n566), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1007), .B1(new_n1014), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n978), .B1(new_n975), .B2(G8), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1025), .A2(new_n1007), .A3(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(new_n979), .A3(new_n996), .A4(new_n987), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1005), .A2(new_n1006), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1956), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT56), .B(G2072), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n972), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n552), .A2(new_n1037), .A3(new_n553), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(new_n562), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1032), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1348), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1015), .A2(new_n1016), .A3(KEYINPUT50), .ZN(new_n1043));
  INV_X1    g618(.A(new_n967), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n981), .A2(G2067), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n600), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1040), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n883), .A2(new_n1037), .B1(new_n562), .B2(new_n1038), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT50), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1009), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1956), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1050), .B1(new_n1053), .B2(new_n1035), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1041), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1041), .A3(KEYINPUT61), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1045), .A2(new_n1046), .A3(KEYINPUT60), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1348), .B1(new_n964), .B2(new_n967), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n981), .A2(G2067), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1064), .A3(new_n884), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1045), .A2(new_n1046), .A3(KEYINPUT60), .A4(new_n600), .ZN(new_n1066));
  INV_X1    g641(.A(new_n972), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT58), .B(G1341), .Z(new_n1068));
  AOI22_X1  g643(.A1(new_n1067), .A2(new_n934), .B1(new_n981), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT59), .A3(new_n541), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1069), .B2(new_n540), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1065), .A2(new_n1066), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1049), .B1(new_n1059), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n970), .A2(new_n1076), .A3(new_n971), .A4(new_n932), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1077), .A2(KEYINPUT121), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT121), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g655(.A(G301), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1078), .A2(G2078), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1017), .A2(new_n1082), .A3(new_n1019), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT119), .B(G1961), .Z(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n964), .B2(new_n967), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT120), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1084), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1017), .A2(new_n1019), .A3(new_n1082), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1081), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1077), .A2(KEYINPUT121), .A3(new_n1078), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(G40), .B(new_n1082), .C1(new_n463), .C2(G2105), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n464), .A2(KEYINPUT122), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n466), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n464), .A2(KEYINPUT122), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n971), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n930), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1085), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G301), .B1(new_n1097), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n1092), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(G171), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT54), .B1(new_n1108), .B2(new_n1105), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1111), .B2(G301), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n960), .A2(new_n963), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1018), .B1(new_n1113), .B2(new_n969), .ZN(new_n1114));
  OAI211_X1 g689(.A(G168), .B(new_n1023), .C1(new_n1114), .C2(G1966), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G8), .ZN(new_n1116));
  AOI21_X1  g691(.A(G168), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT51), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1119), .A3(G8), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1107), .A2(new_n1112), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1091), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1089), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1097), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G171), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(KEYINPUT62), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1118), .A2(new_n1128), .A3(new_n1120), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1075), .A2(new_n1121), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1030), .B1(new_n1130), .B2(new_n1014), .ZN(new_n1131));
  AND2_X1   g706(.A1(G290), .A2(G1986), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n933), .B1(new_n1132), .B2(new_n951), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n947), .A2(new_n1133), .A3(new_n949), .A4(new_n950), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT113), .Z(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT123), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1075), .A2(new_n1137), .A3(new_n1126), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1126), .A2(KEYINPUT62), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1125), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n1129), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1014), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(KEYINPUT123), .B(new_n1135), .C1(new_n1142), .C2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n958), .B1(new_n1136), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT125), .B(new_n958), .C1(new_n1136), .C2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g727(.A1(new_n460), .A2(G227), .ZN(new_n1154));
  AND3_X1   g728(.A1(new_n693), .A2(new_n694), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n1155), .A2(new_n652), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1156), .A2(KEYINPUT126), .ZN(new_n1157));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1158));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n652), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g733(.A1(new_n915), .A2(new_n921), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g734(.A1(new_n1160), .A2(KEYINPUT127), .A3(new_n881), .ZN(new_n1161));
  AOI21_X1  g735(.A(KEYINPUT127), .B1(new_n1160), .B2(new_n881), .ZN(new_n1162));
  NOR2_X1   g736(.A1(new_n1161), .A2(new_n1162), .ZN(G308));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n881), .ZN(G225));
endmodule


