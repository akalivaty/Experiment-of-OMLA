//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  INV_X1    g000(.A(G183gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT27), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(KEYINPUT27), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT28), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT26), .B1(new_n209), .B2(new_n210), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n204), .A2(new_n217), .B1(KEYINPUT67), .B2(new_n203), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n217), .B2(new_n204), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n203), .B2(KEYINPUT67), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n207), .B(new_n216), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n208), .A2(KEYINPUT24), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n205), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n202), .A2(new_n205), .A3(KEYINPUT65), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT23), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n232), .A2(new_n234), .A3(new_n214), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n231), .A2(KEYINPUT66), .A3(KEYINPUT25), .A4(new_n235), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n232), .A2(new_n234), .A3(new_n214), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n227), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(KEYINPUT64), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n223), .A2(new_n225), .B1(new_n202), .B2(new_n205), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT25), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n222), .B1(new_n240), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT73), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT1), .B1(new_n251), .B2(KEYINPUT69), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(KEYINPUT69), .B2(new_n251), .ZN(new_n253));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G113gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G113gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(G120gat), .ZN(new_n263));
  OR2_X1    g062(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(G113gat), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n258), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n258), .B2(new_n267), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n256), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n235), .B1(new_n244), .B2(new_n245), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(new_n238), .A3(new_n239), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT73), .A3(new_n222), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n250), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G227gat), .ZN(new_n280));
  INV_X1    g079(.A(G233gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n271), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n269), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n248), .A2(new_n249), .A3(new_n256), .A4(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n279), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n282), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT32), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(new_n288), .B2(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT75), .ZN(new_n296));
  XNOR2_X1  g095(.A(G15gat), .B(G43gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G71gat), .B(G99gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT33), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n290), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n279), .A2(new_n285), .ZN(new_n303));
  INV_X1    g102(.A(new_n282), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n305), .A2(KEYINPUT34), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(KEYINPUT34), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n299), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n309), .A2(KEYINPUT76), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT33), .B1(new_n309), .B2(KEYINPUT76), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n295), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n302), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n302), .A2(new_n312), .ZN(new_n314));
  INV_X1    g113(.A(new_n308), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(new_n319), .B1(G211gat), .B2(G218gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n318), .B2(new_n319), .ZN(new_n321));
  XNOR2_X1  g120(.A(G197gat), .B(G204gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G211gat), .B(G218gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n317), .B1(new_n325), .B2(KEYINPUT29), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT82), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT82), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(G141gat), .B(G148gat), .Z(new_n335));
  OR2_X1    g134(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n336));
  NAND2_X1  g135(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n332), .B1(new_n329), .B2(KEYINPUT2), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n334), .A2(new_n338), .B1(new_n339), .B2(new_n335), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n317), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n325), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G22gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n342), .A2(G22gat), .A3(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G228gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(new_n281), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT31), .B(G50gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT87), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n351), .A2(new_n353), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n355), .A2(new_n361), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n358), .B(KEYINPUT87), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n222), .B(new_n368), .C1(new_n240), .C2(new_n247), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n277), .A2(new_n222), .B1(new_n344), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n325), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n344), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n248), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n325), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n369), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  XOR2_X1   g179(.A(new_n380), .B(KEYINPUT80), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n372), .A2(new_n376), .A3(KEYINPUT30), .A4(new_n380), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n372), .A2(new_n376), .A3(new_n380), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n372), .A2(new_n376), .A3(KEYINPUT81), .A4(new_n380), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n272), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n256), .B(KEYINPUT84), .C1(new_n270), .C2(new_n271), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .A4(new_n343), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n256), .B(new_n340), .C1(new_n270), .C2(new_n271), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n284), .A2(new_n400), .A3(new_n256), .A4(new_n340), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n394), .A2(new_n341), .A3(new_n395), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n405), .A2(new_n398), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT5), .B(new_n404), .C1(new_n406), .C2(new_n403), .ZN(new_n407));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT0), .ZN(new_n409));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n399), .A2(new_n401), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n398), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(KEYINPUT85), .A3(new_n400), .ZN(new_n415));
  INV_X1    g214(.A(new_n403), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n413), .A2(new_n397), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n407), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n411), .B1(new_n407), .B2(new_n418), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n420), .B(new_n411), .C1(new_n407), .C2(new_n418), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n392), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(KEYINPUT35), .ZN(new_n426));
  AND4_X1   g225(.A1(new_n313), .A2(new_n316), .A3(new_n367), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT77), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n316), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n313), .A2(new_n367), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n411), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n403), .B1(new_n405), .B2(new_n398), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT5), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n418), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n420), .A3(new_n419), .ZN(new_n440));
  INV_X1    g239(.A(new_n424), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT86), .A3(new_n392), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n314), .A2(KEYINPUT77), .A3(new_n315), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n427), .B1(new_n446), .B2(KEYINPUT35), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n443), .A3(new_n366), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n423), .A2(new_n424), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT37), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n372), .A2(new_n450), .A3(new_n376), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n381), .A2(KEYINPUT38), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT89), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n377), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n325), .A2(new_n453), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT37), .B1(new_n372), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n451), .B(new_n452), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n380), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n450), .B1(new_n372), .B2(new_n376), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT38), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AND4_X1   g260(.A1(new_n388), .A2(new_n457), .A3(new_n390), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n366), .B1(new_n449), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n405), .A2(new_n398), .A3(new_n403), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT39), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n413), .A2(new_n397), .A3(new_n415), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n416), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(new_n416), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n411), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n465), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n416), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(KEYINPUT39), .A3(new_n466), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(KEYINPUT40), .A3(new_n411), .A4(new_n471), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n439), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n464), .B1(new_n477), .B2(new_n392), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n411), .A3(new_n471), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n422), .B1(new_n479), .B2(new_n465), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n385), .A2(new_n391), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(KEYINPUT88), .A3(new_n481), .A4(new_n476), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n448), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n313), .A2(KEYINPUT36), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n429), .A2(new_n486), .A3(new_n445), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n316), .A2(new_n313), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT78), .B(KEYINPUT36), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n447), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G197gat), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT11), .B(G169gat), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT12), .ZN(new_n497));
  XOR2_X1   g296(.A(G15gat), .B(G22gat), .Z(new_n498));
  INV_X1    g297(.A(KEYINPUT95), .ZN(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT95), .B1(new_n502), .B2(G1gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT94), .ZN(new_n504));
  AND2_X1   g303(.A1(KEYINPUT93), .A2(G1gat), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT16), .B1(KEYINPUT93), .B2(G1gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n501), .B(new_n503), .C1(new_n504), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OR3_X1    g309(.A1(new_n502), .A2(G1gat), .A3(G8gat), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n508), .A2(G8gat), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G43gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(G50gat), .ZN(new_n514));
  INV_X1    g313(.A(G50gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G43gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT90), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(KEYINPUT15), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT14), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(G29gat), .A2(G36gat), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  OR2_X1    g328(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n531));
  AOI21_X1  g330(.A(G50gat), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n514), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n521), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G43gat), .B(G50gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n529), .B1(new_n536), .B2(new_n519), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT91), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n527), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT91), .B1(new_n524), .B2(new_n526), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n518), .B(new_n537), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n512), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT13), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n535), .A2(new_n541), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n535), .B2(new_n541), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n548), .B(new_n512), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n508), .A2(G8gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n510), .A2(new_n511), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n542), .A2(KEYINPUT17), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n535), .A2(new_n541), .A3(new_n549), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n542), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT96), .B1(new_n559), .B2(new_n512), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n552), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n544), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n547), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(KEYINPUT18), .A3(new_n544), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n497), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n497), .A3(new_n565), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G57gat), .B(G64gat), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G57gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G64gat), .ZN(new_n578));
  INV_X1    g377(.A(G64gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G57gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G71gat), .B(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n575), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n576), .A2(new_n584), .A3(KEYINPUT97), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n555), .B1(new_n589), .B2(KEYINPUT21), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT98), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n327), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n576), .A2(new_n584), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G127gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G183gat), .B(G211gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n594), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n606));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G99gat), .B(G106gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT8), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  INV_X1    g416(.A(G92gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n614), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n611), .A2(new_n612), .ZN(new_n621));
  NAND3_X1  g420(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(KEYINPUT7), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n610), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n625));
  AND4_X1   g424(.A1(new_n610), .A2(new_n623), .A3(new_n614), .A4(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT100), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n624), .A2(new_n626), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n627), .B(new_n630), .C1(new_n550), .C2(new_n551), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n542), .A2(new_n628), .B1(KEYINPUT41), .B2(new_n605), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n631), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n631), .A2(new_n633), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT101), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n641), .B2(new_n634), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n609), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n637), .B1(new_n635), .B2(new_n636), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n634), .A3(new_n639), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n608), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n604), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n610), .ZN(new_n650));
  INV_X1    g449(.A(new_n623), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n625), .A2(new_n614), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n620), .A2(new_n610), .A3(new_n623), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(KEYINPUT102), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n595), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n576), .A3(new_n584), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n624), .B2(new_n626), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n628), .A2(KEYINPUT10), .A3(new_n588), .A4(new_n587), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(new_n658), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n662), .A2(KEYINPUT103), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n675), .A3(new_n661), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n663), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n667), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n665), .A2(KEYINPUT104), .A3(new_n666), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n671), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n673), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  NOR4_X1   g482(.A1(new_n492), .A2(new_n570), .A3(new_n649), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n449), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n481), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n684), .A2(KEYINPUT105), .A3(new_n481), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(G8gat), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT106), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n481), .A4(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n689), .B2(new_n690), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n691), .B(new_n695), .C1(new_n696), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g496(.A(G15gat), .ZN(new_n698));
  INV_X1    g497(.A(new_n488), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n487), .A2(new_n490), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n700), .B1(new_n704), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n684), .A2(new_n366), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  OAI21_X1  g507(.A(new_n647), .B1(new_n447), .B2(new_n491), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(KEYINPUT44), .B(new_n647), .C1(new_n447), .C2(new_n491), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n570), .A2(new_n603), .A3(new_n683), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n711), .A2(new_n449), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G29gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n647), .B(new_n713), .C1(new_n447), .C2(new_n491), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n442), .A2(G29gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n709), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n721), .A2(KEYINPUT45), .A3(new_n713), .A4(new_n718), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n715), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1328gat));
  NAND4_X1  g524(.A1(new_n711), .A2(new_n481), .A3(new_n712), .A4(new_n713), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G36gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n392), .A2(G36gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT46), .B1(new_n717), .B2(new_n729), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n717), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT108), .ZN(G1329gat));
  NAND2_X1  g532(.A1(new_n530), .A2(new_n531), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n717), .A2(new_n488), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n711), .A2(new_n702), .A3(new_n712), .A4(new_n713), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n734), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n734), .ZN(new_n743));
  INV_X1    g542(.A(new_n735), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT109), .B1(new_n745), .B2(new_n736), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n735), .B1(new_n738), .B2(new_n734), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT47), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n742), .B1(new_n746), .B2(new_n749), .ZN(G1330gat));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n752));
  OAI21_X1  g551(.A(G50gat), .B1(new_n752), .B2(new_n367), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n721), .A2(new_n515), .A3(new_n366), .A4(new_n713), .ZN(new_n754));
  AOI211_X1 g553(.A(KEYINPUT111), .B(new_n751), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n751), .A2(KEYINPUT111), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(KEYINPUT111), .ZN(new_n757));
  AND4_X1   g556(.A1(new_n756), .A2(new_n753), .A3(new_n757), .A4(new_n754), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n755), .A2(new_n758), .ZN(G1331gat));
  NOR2_X1   g558(.A1(new_n649), .A2(new_n569), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n683), .B(new_n760), .C1(new_n447), .C2(new_n491), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n442), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n577), .ZN(G1332gat));
  NOR3_X1   g562(.A1(new_n492), .A2(new_n569), .A3(new_n649), .ZN(new_n764));
  INV_X1    g563(.A(new_n683), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n392), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT49), .B(G64gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n764), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1333gat));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n764), .A2(new_n774), .A3(new_n699), .A4(new_n683), .ZN(new_n775));
  INV_X1    g574(.A(G71gat), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT113), .B1(new_n761), .B2(new_n488), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n761), .A2(new_n776), .A3(new_n701), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT50), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n782), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1334gat));
  NOR2_X1   g583(.A1(new_n761), .A2(new_n367), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT114), .B(G78gat), .Z(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1335gat));
  NOR3_X1   g586(.A1(new_n603), .A2(new_n569), .A3(new_n765), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n711), .A2(new_n712), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n442), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n603), .A2(new_n569), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n647), .B(new_n791), .C1(new_n447), .C2(new_n491), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n683), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n449), .A2(new_n617), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(G1336gat));
  XNOR2_X1  g596(.A(new_n792), .B(KEYINPUT51), .ZN(new_n798));
  INV_X1    g597(.A(new_n766), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n618), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n392), .A2(new_n618), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n711), .A2(new_n712), .A3(new_n788), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n800), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n803), .B1(new_n800), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(G1337gat));
  OAI21_X1  g609(.A(G99gat), .B1(new_n789), .B2(new_n701), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n488), .A2(G99gat), .A3(new_n765), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT116), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n798), .B2(new_n813), .ZN(G1338gat));
  OAI21_X1  g613(.A(G106gat), .B1(new_n789), .B2(new_n367), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n367), .A2(G106gat), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n795), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n815), .C1(new_n795), .C2(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1339gat));
  NAND3_X1  g621(.A1(new_n648), .A2(new_n570), .A3(new_n765), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT54), .B(new_n666), .C1(new_n660), .C2(new_n661), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT117), .B1(new_n824), .B2(new_n671), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n662), .A2(new_n826), .A3(new_n663), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n672), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n660), .A2(new_n666), .A3(new_n661), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n677), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n543), .A2(new_n546), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n561), .B2(new_n544), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n496), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n647), .A2(new_n568), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n678), .A2(new_n682), .ZN(new_n841));
  AND4_X1   g640(.A1(KEYINPUT118), .A2(new_n830), .A3(KEYINPUT55), .A4(new_n833), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n825), .A2(new_n829), .B1(new_n677), .B2(new_n832), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT118), .B1(new_n843), .B2(KEYINPUT55), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n568), .A2(new_n683), .A3(new_n839), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n568), .A2(new_n839), .A3(new_n683), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n562), .A2(new_n563), .ZN(new_n851));
  INV_X1    g650(.A(new_n547), .ZN(new_n852));
  AND4_X1   g651(.A1(new_n497), .A2(new_n851), .A3(new_n565), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n836), .B1(new_n853), .B2(new_n566), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n848), .B(new_n850), .C1(new_n845), .C2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n647), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n846), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n604), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT120), .B(new_n846), .C1(new_n856), .C2(new_n855), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n823), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n449), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n429), .A2(new_n430), .A3(new_n445), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n392), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n865), .A2(new_n260), .A3(new_n262), .A4(new_n569), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n488), .A2(new_n366), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n442), .A2(new_n481), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n861), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G113gat), .B1(new_n869), .B2(new_n570), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n870), .ZN(G1340gat));
  NAND4_X1  g670(.A1(new_n865), .A2(new_n264), .A3(new_n265), .A4(new_n683), .ZN(new_n872));
  OAI21_X1  g671(.A(G120gat), .B1(new_n869), .B2(new_n765), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n865), .A2(new_n599), .A3(new_n603), .ZN(new_n875));
  OAI21_X1  g674(.A(G127gat), .B1(new_n869), .B2(new_n604), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1342gat));
  NAND2_X1  g676(.A1(new_n392), .A2(new_n647), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(G134gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n869), .B2(new_n856), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G1343gat));
  AND2_X1   g683(.A1(new_n701), .A2(new_n868), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n861), .B2(new_n366), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n847), .B1(new_n845), .B2(new_n854), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n846), .B1(new_n887), .B2(new_n856), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n823), .B1(new_n888), .B2(new_n603), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n366), .A2(KEYINPUT57), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n885), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G141gat), .B1(new_n892), .B2(new_n570), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT58), .B1(new_n893), .B2(KEYINPUT121), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n702), .A2(new_n367), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n862), .A2(new_n895), .A3(new_n392), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n570), .A2(G141gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n894), .B(new_n898), .Z(G1344gat));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n861), .A2(new_n890), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n889), .B2(new_n366), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n683), .B(new_n885), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n683), .B(new_n885), .C1(new_n886), .C2(new_n891), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n901), .A2(G148gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(KEYINPUT122), .A3(new_n907), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n896), .A2(G148gat), .A3(new_n765), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n900), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n913), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n906), .A2(KEYINPUT122), .A3(new_n907), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT122), .B1(new_n906), .B2(new_n907), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT123), .B(new_n915), .C1(new_n918), .C2(new_n905), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n914), .A2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n892), .B2(new_n604), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n603), .A2(new_n327), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n896), .B2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n892), .B2(new_n856), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n878), .A2(G162gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n862), .A2(new_n895), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n449), .A2(new_n392), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n861), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n863), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n209), .A3(new_n569), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n867), .ZN(new_n932));
  OAI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n570), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT124), .ZN(G1348gat));
  AOI21_X1  g734(.A(G176gat), .B1(new_n930), .B2(new_n683), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n929), .A2(G176gat), .A3(new_n867), .A4(new_n683), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(G1349gat));
  NAND4_X1  g740(.A1(new_n930), .A2(new_n203), .A3(new_n204), .A4(new_n603), .ZN(new_n942));
  OAI21_X1  g741(.A(G183gat), .B1(new_n932), .B2(new_n604), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n932), .B2(new_n856), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT61), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n205), .A3(new_n647), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1351gat));
  NAND2_X1  g748(.A1(new_n929), .A2(new_n895), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n569), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n902), .A2(new_n903), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n701), .A2(new_n928), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n569), .A2(G197gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  INV_X1    g756(.A(new_n955), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n958), .B2(new_n765), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n765), .A2(G204gat), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT62), .B1(new_n950), .B2(new_n960), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n950), .A2(KEYINPUT62), .A3(new_n960), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n959), .B(new_n961), .C1(new_n963), .C2(new_n964), .ZN(G1353gat));
  NAND2_X1  g764(.A1(new_n955), .A2(new_n603), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G211gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT63), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n969), .A3(G211gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n950), .A2(G211gat), .A3(new_n604), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT127), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(G218gat), .B1(new_n958), .B2(new_n856), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n856), .A2(G218gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n950), .B2(new_n975), .ZN(G1355gat));
endmodule


