//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT64), .B1(new_n189), .B2(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n192), .A3(G143), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n197), .A2(new_n199), .A3(new_n194), .A4(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G134), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(new_n208), .B2(KEYINPUT11), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT65), .B1(new_n204), .B2(G134), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(G137), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n203), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n189), .A2(G146), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n192), .A2(G143), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n221), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n197), .A2(new_n199), .A3(new_n194), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n216), .B1(new_n211), .B2(new_n212), .ZN(new_n228));
  AOI211_X1 g042(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n204), .C2(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n227), .B1(new_n230), .B2(new_n214), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n188), .B1(new_n219), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(G116), .B(G119), .Z(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n233), .A2(KEYINPUT66), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT2), .B(G113), .Z(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(G116), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n236), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  OAI22_X1  g057(.A1(new_n235), .A2(new_n243), .B1(new_n237), .B2(new_n242), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n224), .A2(new_n226), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n228), .A2(G131), .A3(new_n229), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n210), .B1(new_n209), .B2(new_n213), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n203), .A2(new_n214), .A3(new_n218), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(KEYINPUT30), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n232), .A2(new_n244), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n230), .A2(new_n214), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n196), .A2(new_n202), .B1(G131), .B2(new_n217), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n252), .A2(new_n245), .B1(new_n253), .B2(new_n214), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n237), .A2(new_n242), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT66), .B1(new_n233), .B2(new_n234), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n237), .A2(new_n242), .A3(new_n236), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n251), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT27), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n263), .A2(KEYINPUT26), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(KEYINPUT26), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n264), .A2(G101), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(G101), .B1(new_n264), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT67), .B(KEYINPUT31), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n260), .A2(KEYINPUT68), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n251), .A2(new_n259), .ZN(new_n271));
  INV_X1    g085(.A(new_n268), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT31), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n251), .A2(new_n268), .A3(new_n259), .A4(new_n269), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n270), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n248), .A2(new_n249), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n244), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT69), .B1(new_n254), .B2(new_n258), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n281), .A3(new_n244), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT70), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n278), .B2(new_n244), .ZN(new_n286));
  AOI211_X1 g100(.A(KEYINPUT69), .B(new_n258), .C1(new_n248), .C2(new_n249), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n259), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT28), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n285), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n277), .B1(new_n293), .B2(new_n272), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n272), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n270), .A2(new_n273), .A3(new_n276), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(KEYINPUT32), .A3(new_n295), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n272), .A2(new_n291), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n285), .A2(new_n290), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n271), .B2(new_n272), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT72), .B(G902), .Z(new_n310));
  NAND2_X1  g124(.A1(new_n303), .A2(KEYINPUT29), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n254), .B(new_n244), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(new_n284), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n310), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n307), .A2(new_n309), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n316), .A2(new_n317), .A3(G472), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(new_n316), .B2(G472), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n302), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G137), .ZN(new_n321));
  INV_X1    g135(.A(G953), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(G221), .A3(G234), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G125), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT75), .ZN(new_n332));
  OR3_X1    g146(.A1(new_n330), .A2(KEYINPUT75), .A3(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n329), .A2(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(G146), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G125), .B(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n192), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n239), .B2(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n342), .B(new_n343), .C1(G119), .C2(new_n200), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT76), .B(G110), .ZN(new_n345));
  XNOR2_X1  g159(.A(G119), .B(G128), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT24), .B(G110), .Z(new_n347));
  OAI22_X1  g161(.A1(new_n344), .A2(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n338), .A2(new_n340), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(G110), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n346), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n330), .A2(KEYINPUT75), .A3(G140), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n339), .B2(KEYINPUT75), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT16), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n337), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n192), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n353), .B1(new_n358), .B2(new_n338), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n327), .B1(new_n350), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n338), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n351), .A2(new_n352), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n349), .A3(new_n326), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n310), .ZN(new_n366));
  INV_X1    g180(.A(G234), .ZN(new_n367));
  OAI21_X1  g181(.A(G217), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n368), .B(KEYINPUT74), .Z(new_n369));
  NOR3_X1   g183(.A1(new_n365), .A2(G902), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n366), .B1(new_n360), .B2(new_n364), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI211_X1 g188(.A(KEYINPUT25), .B(new_n366), .C1(new_n360), .C2(new_n364), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n370), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT9), .B(G234), .ZN(new_n378));
  OAI21_X1  g192(.A(G221), .B1(new_n378), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n322), .A2(G227), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g197(.A(new_n252), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n197), .A2(new_n199), .A3(new_n194), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n191), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n202), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT3), .B1(new_n388), .B2(G107), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(G104), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n388), .A2(G107), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n389), .A2(new_n392), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n388), .A2(G107), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n391), .A2(G104), .ZN(new_n397));
  OAI21_X1  g211(.A(G101), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n387), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n389), .A2(new_n392), .A3(new_n394), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n393), .A2(KEYINPUT79), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n406), .B2(new_n395), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT4), .B1(new_n404), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n245), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n196), .B2(new_n202), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n399), .ZN(new_n412));
  AND4_X1   g226(.A1(new_n384), .A2(new_n402), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n400), .A2(new_n401), .B1(new_n399), .B2(new_n411), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n384), .B1(new_n414), .B2(new_n409), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n383), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n384), .A3(new_n409), .ZN(new_n417));
  INV_X1    g231(.A(new_n383), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n395), .A2(new_n398), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n196), .A3(new_n202), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n400), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n421), .A2(KEYINPUT12), .A3(new_n252), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT12), .B1(new_n421), .B2(new_n252), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n417), .B(new_n418), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n366), .B1(new_n416), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G469), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT81), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n429), .A3(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n423), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n421), .A2(KEYINPUT12), .A3(new_n252), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n418), .B1(new_n435), .B2(new_n417), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n417), .A2(new_n418), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n415), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n432), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G469), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n380), .B1(new_n431), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n244), .B1(new_n407), .B2(new_n408), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n447));
  OR2_X1    g261(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n448), .A2(G116), .A3(new_n239), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G113), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n448), .A2(new_n449), .B1(new_n240), .B2(new_n241), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n449), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n242), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(KEYINPUT83), .A3(G113), .A4(new_n450), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n419), .B1(new_n257), .B2(new_n256), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n446), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n446), .A2(new_n459), .A3(new_n461), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n227), .A2(G125), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n196), .A2(new_n330), .A3(new_n202), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n322), .A2(G224), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n471), .A3(new_n462), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n465), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n461), .B(KEYINPUT8), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n256), .A2(new_n257), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n399), .B1(new_n457), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT5), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n450), .B(G113), .C1(new_n233), .C2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT84), .B1(new_n458), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n458), .A2(KEYINPUT84), .A3(new_n479), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n469), .B2(KEYINPUT86), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n468), .B(new_n485), .C1(KEYINPUT86), .C2(new_n469), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n469), .A2(KEYINPUT7), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT85), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n467), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n466), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n467), .A2(new_n488), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n464), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n432), .B1(new_n483), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n445), .B1(new_n473), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n481), .A2(new_n482), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n474), .ZN(new_n497));
  INV_X1    g311(.A(new_n493), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n465), .A2(new_n470), .A3(new_n472), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n444), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n443), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n441), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n388), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n332), .A2(new_n333), .A3(G146), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT88), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n332), .A2(new_n333), .A3(new_n508), .A4(G146), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n340), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n261), .A2(G214), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n189), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n210), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n516));
  AOI21_X1  g330(.A(G143), .B1(new_n261), .B2(G214), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(G131), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n514), .A2(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n510), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n510), .A2(new_n520), .A3(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n514), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n512), .A2(new_n210), .A3(new_n513), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n514), .A2(KEYINPUT17), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n358), .A3(new_n338), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n505), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n505), .B(KEYINPUT91), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n525), .A2(new_n533), .A3(new_n531), .A4(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n510), .A2(new_n520), .A3(KEYINPUT89), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT89), .B1(new_n510), .B2(new_n520), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n531), .B(new_n534), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT92), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n532), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G475), .B1(new_n540), .B2(G902), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n535), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n526), .A2(new_n528), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT19), .ZN(new_n545));
  OR3_X1    g359(.A1(new_n334), .A2(KEYINPUT90), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n339), .A2(new_n545), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT90), .B1(new_n334), .B2(new_n545), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n338), .B(new_n544), .C1(new_n549), .C2(G146), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n505), .B1(new_n525), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n543), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G475), .A2(G902), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n542), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n551), .B1(new_n535), .B2(new_n539), .ZN(new_n556));
  INV_X1    g370(.A(new_n554), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n556), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n541), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT95), .B(G952), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G953), .ZN(new_n562));
  NAND2_X1  g376(.A1(G234), .A2(G237), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n366), .A2(G953), .A3(new_n563), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G116), .B(G122), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n391), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT14), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n238), .A2(KEYINPUT14), .A3(G122), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(G107), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n189), .A2(G128), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT94), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n189), .A2(G128), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n207), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n207), .B1(new_n580), .B2(new_n582), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n574), .B(new_n578), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n573), .A2(new_n391), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n571), .B(KEYINPUT93), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G107), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n583), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n580), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT13), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n581), .B1(new_n580), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n207), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n586), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n378), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n597), .A2(G217), .A3(new_n322), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n586), .B(new_n598), .C1(new_n590), .C2(new_n595), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n310), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G478), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(KEYINPUT15), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n603), .B(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n560), .A2(new_n570), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n503), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n320), .A2(new_n377), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT96), .B(G101), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G3));
  NAND2_X1  g426(.A1(new_n601), .A2(KEYINPUT33), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n598), .B(KEYINPUT97), .Z(new_n615));
  NAND3_X1  g429(.A1(new_n596), .A2(KEYINPUT98), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT98), .B1(new_n596), .B2(new_n615), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT99), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n614), .B(new_n621), .C1(new_n618), .C2(new_n617), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n600), .B2(new_n602), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n366), .A2(new_n604), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n620), .A2(new_n622), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n603), .A2(new_n604), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n559), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n502), .A2(new_n570), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT100), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n630), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n559), .A4(new_n628), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n366), .B1(new_n298), .B2(new_n299), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  OAI22_X1  g451(.A1(new_n636), .A2(new_n637), .B1(new_n294), .B2(new_n296), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n416), .A2(new_n424), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n429), .A2(new_n639), .A3(new_n426), .A4(new_n310), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n429), .B1(new_n425), .B2(new_n426), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n440), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n377), .A3(new_n379), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND3_X1  g461(.A1(new_n553), .A2(new_n542), .A3(new_n554), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT20), .B1(new_n556), .B2(new_n557), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n606), .A3(new_n541), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n630), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n363), .A2(new_n349), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n326), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n369), .A2(G902), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n660), .B1(new_n373), .B2(new_n375), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT101), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n660), .B(new_n663), .C1(new_n373), .C2(new_n375), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n662), .A2(KEYINPUT102), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT102), .B1(new_n662), .B2(new_n664), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n638), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n609), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  INV_X1    g485(.A(new_n667), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n564), .B1(new_n566), .B2(G900), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n650), .A2(new_n606), .A3(new_n541), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n503), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n320), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  AND2_X1   g491(.A1(new_n495), .A2(new_n501), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n662), .A2(new_n664), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n679), .A2(new_n443), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n606), .A3(new_n559), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n673), .B(KEYINPUT39), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n441), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT40), .ZN(new_n685));
  AOI21_X1  g499(.A(G902), .B1(new_n272), .B2(new_n312), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n260), .A2(new_n272), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n297), .A2(new_n301), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n682), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT103), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  NAND3_X1  g508(.A1(new_n628), .A2(new_n559), .A3(new_n673), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n503), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n320), .A2(new_n672), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  NOR2_X1   g512(.A1(new_n425), .A2(new_n426), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n380), .B(new_n699), .C1(new_n428), .C2(new_n430), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n635), .A2(new_n320), .A3(new_n377), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND4_X1  g517(.A1(new_n320), .A2(new_n377), .A3(new_n652), .A4(new_n700), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n502), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n608), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n320), .A2(new_n672), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT104), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n304), .A2(new_n308), .A3(new_n305), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n308), .B1(new_n304), .B2(new_n305), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n711), .A3(new_n314), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT73), .B1(new_n712), .B2(new_n637), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n316), .A2(new_n317), .A3(G472), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n667), .B1(new_n715), .B2(new_n302), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n707), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n709), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n559), .A2(new_n606), .A3(new_n502), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n570), .A3(new_n700), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n313), .A2(new_n291), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n268), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n295), .B1(new_n726), .B2(new_n277), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT105), .B(G472), .Z(new_n728));
  OAI211_X1 g542(.A(new_n727), .B(new_n377), .C1(new_n636), .C2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n721), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n699), .B1(new_n428), .B2(new_n430), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n379), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n722), .A2(new_n732), .A3(new_n569), .ZN(new_n733));
  INV_X1    g547(.A(new_n729), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  OAI211_X1 g551(.A(new_n680), .B(new_n727), .C1(new_n636), .C2(new_n728), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n738), .A2(new_n706), .A3(new_n695), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n330), .ZN(G27));
  NAND2_X1  g554(.A1(new_n297), .A2(new_n301), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n713), .B2(new_n714), .ZN(new_n742));
  INV_X1    g556(.A(new_n377), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n495), .A2(new_n501), .A3(new_n442), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n495), .A2(new_n501), .A3(new_n747), .A4(new_n442), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n379), .A3(new_n642), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n695), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(KEYINPUT42), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n744), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n320), .A2(new_n377), .A3(new_n750), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n752), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  AND2_X1   g572(.A1(new_n674), .A2(KEYINPUT109), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n674), .A2(KEYINPUT109), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n760), .A3(new_n749), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n320), .A3(new_n377), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  INV_X1    g577(.A(new_n436), .ZN(new_n764));
  INV_X1    g578(.A(new_n438), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(KEYINPUT45), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n436), .B2(new_n438), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(G469), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(G469), .A2(G902), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n431), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n379), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n683), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n746), .A2(new_n748), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n559), .B1(new_n627), .B2(new_n626), .ZN(new_n782));
  MUX2_X1   g596(.A(new_n780), .B(new_n781), .S(new_n782), .Z(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n638), .A3(new_n680), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT111), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n204), .ZN(G39));
  XOR2_X1   g603(.A(new_n776), .B(KEYINPUT47), .Z(new_n790));
  NOR3_X1   g604(.A1(new_n695), .A2(new_n778), .A3(new_n377), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n742), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT112), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  AND2_X1   g608(.A1(new_n783), .A2(new_n565), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n778), .A2(new_n732), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n744), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT48), .Z(new_n799));
  AND2_X1   g613(.A1(new_n795), .A2(new_n734), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n502), .A3(new_n700), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n377), .A2(new_n691), .A3(new_n565), .A4(new_n796), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n559), .A3(new_n628), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n562), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n800), .A2(new_n443), .A3(new_n679), .A4(new_n700), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT50), .Z(new_n806));
  AND2_X1   g620(.A1(new_n731), .A2(new_n380), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n790), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n800), .A2(new_n748), .A3(new_n746), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n809), .B2(KEYINPUT118), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(KEYINPUT118), .B2(new_n809), .ZN(new_n811));
  INV_X1    g625(.A(new_n738), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n628), .A2(new_n559), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n797), .A2(new_n812), .B1(new_n802), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n806), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n799), .B(new_n804), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n660), .B(new_n673), .C1(new_n373), .C2(new_n375), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n642), .A2(new_n379), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n722), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n690), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n824), .B1(new_n823), .B2(new_n690), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n739), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n676), .A3(new_n697), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n739), .B1(new_n716), .B2(new_n675), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .A3(new_n697), .A4(new_n827), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT115), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT115), .B1(new_n831), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n736), .A2(new_n701), .A3(new_n704), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n718), .B2(new_n709), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n630), .B1(new_n629), .B2(new_n651), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n668), .A2(new_n609), .B1(new_n644), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n750), .A2(new_n812), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n762), .A2(new_n840), .A3(new_n610), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n754), .B2(new_n756), .ZN(new_n843));
  INV_X1    g657(.A(new_n673), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n749), .A2(new_n606), .A3(new_n559), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n320), .A3(new_n672), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n716), .A2(new_n848), .A3(new_n845), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n838), .A2(new_n843), .A3(KEYINPUT53), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n819), .B1(new_n836), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n842), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n757), .A3(new_n850), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n719), .A2(new_n701), .A3(new_n704), .A4(new_n736), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n857), .B(KEYINPUT117), .C1(new_n835), .C2(new_n834), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n831), .A2(new_n833), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n838), .A3(new_n843), .A4(new_n850), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n860), .A2(KEYINPUT116), .A3(new_n856), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT116), .B1(new_n860), .B2(new_n856), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n852), .B(new_n858), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n836), .A2(new_n855), .A3(new_n854), .ZN(new_n866));
  MUX2_X1   g680(.A(new_n860), .B(new_n866), .S(new_n856), .Z(new_n867));
  OAI21_X1  g681(.A(new_n864), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n818), .A2(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n377), .A2(new_n679), .A3(new_n379), .A4(new_n442), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n731), .B(KEYINPUT49), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n782), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n869), .B1(new_n690), .B2(new_n872), .ZN(G75));
  NAND3_X1  g687(.A1(new_n863), .A2(new_n366), .A3(new_n445), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n465), .A2(new_n472), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n470), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT121), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n877), .A2(KEYINPUT121), .ZN(new_n879));
  XOR2_X1   g693(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n880));
  NAND4_X1  g694(.A1(new_n874), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n322), .A2(G952), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT122), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT56), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n887), .B2(new_n877), .ZN(G51));
  NAND2_X1  g702(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n864), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n770), .B(KEYINPUT57), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n639), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n769), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n863), .A2(new_n366), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n882), .B1(new_n892), .B2(new_n894), .ZN(G54));
  NAND4_X1  g709(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .A4(new_n366), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n896), .A2(new_n556), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n556), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n882), .ZN(G60));
  AND3_X1   g713(.A1(new_n620), .A2(new_n622), .A3(new_n624), .ZN(new_n900));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n883), .B1(new_n890), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n900), .B1(new_n868), .B2(new_n902), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(G63));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT60), .Z(new_n908));
  AND3_X1   g722(.A1(new_n863), .A2(KEYINPUT123), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT123), .B1(new_n863), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n658), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n863), .A2(new_n908), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n863), .A2(KEYINPUT123), .A3(new_n908), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n365), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n911), .A2(new_n916), .A3(new_n883), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n911), .A2(new_n916), .A3(KEYINPUT61), .A4(new_n883), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(G66));
  NAND3_X1  g735(.A1(new_n838), .A2(new_n610), .A3(new_n840), .ZN(new_n922));
  NAND2_X1  g736(.A1(G224), .A2(G953), .ZN(new_n923));
  OAI22_X1  g737(.A1(new_n922), .A2(G953), .B1(new_n568), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT124), .Z(new_n925));
  INV_X1    g739(.A(G898), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n875), .B1(new_n926), .B2(G953), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n925), .B(new_n927), .ZN(G69));
  AND2_X1   g742(.A1(new_n832), .A2(new_n697), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n693), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n793), .A2(new_n787), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n629), .A2(new_n651), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n684), .A2(new_n778), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n744), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT125), .Z(new_n937));
  NAND4_X1  g751(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n322), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n232), .A2(new_n250), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(new_n549), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(G900), .B2(G953), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n776), .A2(new_n777), .A3(new_n722), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n744), .B1(new_n944), .B2(new_n761), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n932), .A2(new_n757), .A3(new_n929), .A4(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n943), .B1(new_n946), .B2(G953), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n322), .B1(G227), .B2(G900), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G72));
  INV_X1    g764(.A(new_n688), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n271), .A2(new_n268), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n637), .A2(new_n432), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT127), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n867), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n956), .B1(new_n946), .B2(new_n922), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n952), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(G952), .B2(new_n322), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n956), .B1(new_n938), .B2(new_n922), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n959), .B(new_n962), .C1(new_n688), .C2(new_n963), .ZN(G57));
endmodule


