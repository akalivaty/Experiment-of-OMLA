//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(G148gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G141gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n204), .A2(G148gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT72), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT2), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n212), .ZN(new_n215));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(G148gat), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n209), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n214), .A2(new_n217), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G197gat), .B(G204gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230));
  INV_X1    g029(.A(G211gat), .ZN(new_n231));
  INV_X1    g030(.A(G218gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n228), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n225), .B1(new_n236), .B2(KEYINPUT29), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT74), .ZN(new_n239));
  INV_X1    g038(.A(new_n217), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(G155gat), .B2(G162gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n209), .A2(new_n210), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(new_n203), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n244), .B2(new_n211), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n222), .B1(new_n209), .B2(new_n220), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n239), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G141gat), .B(G148gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n213), .B1(new_n248), .B2(KEYINPUT72), .ZN(new_n249));
  INV_X1    g048(.A(new_n211), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n217), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n223), .A2(new_n221), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(KEYINPUT74), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n247), .A3(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n237), .A2(G228gat), .A3(G233gat), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G228gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n235), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n234), .B(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n226), .B2(new_n227), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n227), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n224), .B1(new_n260), .B2(new_n225), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n256), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT77), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT31), .B(G50gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  AOI21_X1  g067(.A(new_n202), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT77), .B1(new_n255), .B2(new_n262), .ZN(new_n270));
  INV_X1    g069(.A(new_n268), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n270), .A2(G22gat), .A3(new_n271), .ZN(new_n272));
  OAI22_X1  g071(.A1(new_n269), .A2(new_n272), .B1(new_n264), .B2(new_n263), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n265), .A2(new_n202), .A3(new_n268), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n263), .A2(new_n264), .ZN(new_n275));
  OAI21_X1  g074(.A(G22gat), .B1(new_n270), .B2(new_n271), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT0), .ZN(new_n280));
  XNOR2_X1  g079(.A(G57gat), .B(G85gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G113gat), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G120gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT1), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G127gat), .A2(G134gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT67), .B(G134gat), .ZN(new_n290));
  INV_X1    g089(.A(G127gat), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G127gat), .A2(G134gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT68), .B1(new_n294), .B2(new_n288), .ZN(new_n295));
  INV_X1    g094(.A(G134gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(new_n293), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n289), .A2(new_n292), .B1(new_n300), .B2(new_n287), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n224), .A2(KEYINPUT4), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT4), .B1(new_n224), .B2(new_n301), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n247), .A2(KEYINPUT3), .A3(new_n253), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n301), .B1(new_n224), .B2(new_n225), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n308), .ZN(new_n310));
  INV_X1    g109(.A(new_n301), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n247), .A2(new_n311), .A3(new_n253), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n247), .A2(new_n311), .A3(new_n253), .A4(KEYINPUT75), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n224), .A2(new_n301), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n310), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n309), .B1(new_n318), .B2(KEYINPUT5), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n307), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n320), .A2(new_n321), .A3(new_n310), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n282), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT6), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT5), .ZN(new_n325));
  INV_X1    g124(.A(new_n282), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n312), .A2(new_n313), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(new_n316), .A3(new_n315), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n321), .B1(new_n328), .B2(new_n310), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n325), .B(new_n326), .C1(new_n329), .C2(new_n309), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n319), .A2(new_n322), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(KEYINPUT6), .A3(new_n326), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  AND4_X1   g140(.A1(KEYINPUT25), .A2(new_n338), .A3(new_n339), .A4(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G183gat), .ZN(new_n343));
  INV_X1    g142(.A(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n348));
  AND2_X1   g147(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n345), .B(new_n346), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n352));
  AND3_X1   g151(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n343), .A2(new_n344), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n345), .B(new_n346), .C1(new_n354), .C2(KEYINPUT24), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n352), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT27), .B1(new_n343), .B2(KEYINPUT66), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G183gat), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n357), .B(new_n344), .C1(KEYINPUT66), .C2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT27), .B(G183gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(G190gat), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n360), .A2(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n337), .A2(KEYINPUT26), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n347), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT26), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n339), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(new_n337), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI22_X1  g170(.A1(new_n351), .A2(new_n356), .B1(new_n364), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n336), .B1(new_n372), .B2(new_n227), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n355), .ZN(new_n374));
  INV_X1    g173(.A(new_n352), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n342), .A2(new_n350), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n360), .A2(new_n361), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n362), .A2(new_n363), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n370), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n335), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n236), .B1(new_n373), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G8gat), .B(G36gat), .Z(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT70), .ZN(new_n385));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n336), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT29), .B1(new_n378), .B2(new_n381), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n388), .B(new_n258), .C1(new_n389), .C2(new_n336), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n383), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT71), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT30), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT30), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(KEYINPUT71), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n383), .A2(new_n390), .ZN(new_n396));
  INV_X1    g195(.A(new_n387), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT76), .B1(new_n334), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  AOI211_X1 g201(.A(new_n402), .B(new_n399), .C1(new_n331), .C2(new_n333), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n278), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n387), .B1(new_n396), .B2(KEYINPUT37), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT38), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT37), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n383), .A2(new_n407), .A3(new_n390), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n391), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n405), .B2(new_n408), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(KEYINPUT80), .B2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n411), .A2(KEYINPUT80), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n412), .A2(new_n333), .A3(new_n331), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n320), .A2(new_n310), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n282), .B1(new_n415), .B2(KEYINPUT39), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT78), .B(new_n282), .C1(new_n415), .C2(KEYINPUT39), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT39), .B1(new_n328), .B2(new_n310), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT79), .B(KEYINPUT39), .C1(new_n328), .C2(new_n310), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n415), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT40), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n420), .A2(KEYINPUT40), .A3(new_n425), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n399), .A2(new_n330), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n278), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n372), .A2(new_n301), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n378), .A2(new_n311), .A3(new_n381), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G227gat), .ZN(new_n437));
  INV_X1    g236(.A(G233gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT34), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n436), .A2(new_n440), .B1(KEYINPUT69), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n434), .A2(new_n435), .A3(new_n439), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT32), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(G15gat), .B(G43gat), .Z(new_n448));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n441), .A2(KEYINPUT69), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n450), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n444), .B(KEYINPUT32), .C1(new_n446), .C2(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n451), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n451), .B2(new_n455), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n443), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n452), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n451), .A2(new_n453), .A3(new_n455), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n442), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT36), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n458), .A2(new_n462), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n404), .A2(new_n433), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n401), .A2(new_n403), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n463), .A2(new_n278), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n399), .B1(new_n331), .B2(new_n333), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n470), .A4(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n465), .A2(new_n470), .A3(new_n277), .A4(new_n273), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n334), .A2(new_n400), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT81), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n469), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT82), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n469), .B(new_n483), .C1(new_n473), .C2(new_n480), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G169gat), .B(G197gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT12), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT87), .B(G29gat), .ZN(new_n492));
  INV_X1    g291(.A(G36gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT85), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OR3_X1    g298(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n494), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G50gat), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n502), .A2(G43gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(G43gat), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT84), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  OR2_X1    g309(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n512));
  AOI21_X1  g311(.A(G43gat), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n513), .B2(new_n503), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n501), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n499), .A2(KEYINPUT86), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n497), .B2(new_n498), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n516), .A2(new_n518), .A3(new_n494), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n505), .A2(new_n508), .A3(KEYINPUT15), .A4(new_n500), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n515), .B(KEYINPUT17), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n516), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n518), .A2(new_n494), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n527), .A2(KEYINPUT91), .A3(KEYINPUT17), .A4(new_n515), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n509), .A2(new_n514), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n526), .B1(new_n501), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT89), .B1(new_n531), .B2(KEYINPUT17), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G8gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT16), .ZN(new_n537));
  AOI21_X1  g336(.A(G1gat), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n536), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n527), .A2(new_n515), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT89), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n529), .A2(new_n532), .A3(new_n540), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n539), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n491), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n546), .A4(new_n547), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n540), .A2(new_n531), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n547), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT93), .B(KEYINPUT13), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n546), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n550), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n548), .A2(new_n549), .B1(new_n555), .B2(new_n557), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT94), .B1(new_n548), .B2(new_n549), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n561), .B(new_n553), .C1(new_n562), .C2(new_n491), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G71gat), .B(G78gat), .Z(new_n565));
  XNOR2_X1  g364(.A(G57gat), .B(G64gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n566), .B2(new_n567), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n565), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT96), .ZN(new_n574));
  XOR2_X1   g373(.A(G57gat), .B(G64gat), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT95), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(new_n568), .A3(new_n571), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n565), .ZN(new_n579));
  INV_X1    g378(.A(G64gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G57gat), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT97), .B(G57gat), .Z(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(new_n580), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n565), .A2(new_n570), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n574), .A2(new_n579), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G231gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(new_n438), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n585), .A2(KEYINPUT21), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n587), .B1(new_n585), .B2(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(KEYINPUT99), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(KEYINPUT99), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n539), .B1(new_n585), .B2(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT20), .ZN(new_n600));
  XOR2_X1   g399(.A(G127gat), .B(G155gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G183gat), .B(G211gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n595), .A2(new_n597), .A3(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT7), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  INV_X1    g414(.A(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(KEYINPUT8), .A2(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G99gat), .B(G106gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n529), .A2(new_n532), .A3(new_n544), .A4(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n541), .B2(new_n621), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT100), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n626), .B1(new_n623), .B2(new_n625), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n612), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n631), .A2(KEYINPUT100), .A3(new_n627), .A4(new_n611), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n583), .A2(new_n584), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n573), .A2(KEYINPUT96), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n578), .B1(new_n577), .B2(new_n565), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n622), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n634), .B(new_n621), .C1(new_n635), .C2(new_n636), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT101), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n585), .A2(new_n643), .A3(KEYINPUT10), .A4(new_n621), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n638), .A2(new_n640), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n647), .A2(new_n650), .A3(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n608), .A2(new_n633), .A3(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n485), .A2(new_n564), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n334), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g462(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n664));
  INV_X1    g463(.A(G8gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n660), .A2(new_n399), .A3(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n667), .A2(KEYINPUT103), .A3(KEYINPUT42), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n485), .A2(new_n564), .A3(new_n659), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n400), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT103), .B1(new_n667), .B2(KEYINPUT42), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n668), .B1(new_n673), .B2(new_n674), .ZN(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n670), .B2(new_n468), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n463), .A2(G15gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n670), .B2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n670), .A2(new_n432), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT43), .B(G22gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(new_n608), .ZN(new_n682));
  INV_X1    g481(.A(new_n633), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n682), .A2(new_n683), .A3(new_n658), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n485), .A2(new_n564), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n661), .A2(new_n492), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n685), .A2(KEYINPUT104), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT104), .B1(new_n685), .B2(new_n687), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n683), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n484), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n465), .A2(new_n277), .A3(new_n273), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n401), .A2(new_n403), .A3(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n479), .B(new_n476), .C1(new_n697), .C2(new_n470), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n483), .B1(new_n698), .B2(new_n469), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n694), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n481), .A2(new_n633), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n693), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n608), .B(KEYINPUT105), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n560), .A2(new_n563), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n658), .B(KEYINPUT106), .Z(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n703), .A2(new_n661), .A3(new_n708), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n691), .A2(new_n692), .B1(new_n492), .B2(new_n709), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n685), .A2(G36gat), .A3(new_n400), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n703), .A2(new_n399), .A3(new_n708), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n493), .B2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  INV_X1    g514(.A(new_n468), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n703), .A2(new_n716), .A3(new_n708), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n685), .A2(G43gat), .A3(new_n463), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n715), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  AOI211_X1 g520(.A(KEYINPUT47), .B(new_n719), .C1(new_n717), .C2(G43gat), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  NAND4_X1  g522(.A1(new_n700), .A2(new_n278), .A3(new_n702), .A4(new_n708), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n511), .A2(new_n512), .ZN(new_n725));
  INV_X1    g524(.A(new_n685), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n432), .A2(new_n725), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT107), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n729), .A2(KEYINPUT108), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(KEYINPUT108), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n730), .A2(KEYINPUT108), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n734), .ZN(G1331gat));
  NAND4_X1  g534(.A1(new_n707), .A2(new_n705), .A3(new_n682), .A4(new_n683), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n698), .B2(new_n469), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n661), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n582), .ZN(G1332gat));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n399), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT49), .B(G64gat), .Z(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n737), .A2(new_n744), .A3(new_n465), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n737), .A2(new_n716), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n744), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g547(.A1(new_n737), .A2(new_n278), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  INV_X1    g549(.A(new_n658), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n682), .A2(new_n564), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n700), .A2(new_n702), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT109), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n700), .A2(new_n755), .A3(new_n702), .A4(new_n752), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n661), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT110), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n754), .A2(new_n759), .A3(new_n661), .A4(new_n756), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(G85gat), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n481), .A2(new_n705), .A3(new_n608), .A4(new_n633), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT51), .Z(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n751), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n616), .A3(new_n661), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n761), .A2(new_n766), .ZN(G1336gat));
  NAND3_X1  g566(.A1(new_n754), .A2(new_n399), .A3(new_n756), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n762), .B(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n706), .A2(G92gat), .A3(new_n400), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n768), .A2(G92gat), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n753), .A2(new_n400), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n617), .ZN(new_n775));
  INV_X1    g574(.A(new_n771), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n764), .B2(new_n776), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n772), .A2(new_n773), .B1(new_n775), .B2(new_n777), .ZN(G1337gat));
  INV_X1    g577(.A(G99gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n765), .A2(new_n779), .A3(new_n465), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n754), .A2(new_n716), .A3(new_n756), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(new_n779), .ZN(G1338gat));
  NOR3_X1   g581(.A1(new_n706), .A2(G106gat), .A3(new_n432), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT53), .B1(new_n763), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT112), .B1(new_n753), .B2(new_n432), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G106gat), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n753), .A2(KEYINPUT112), .A3(new_n432), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n754), .A2(new_n278), .A3(new_n756), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n789), .A2(G106gat), .B1(new_n770), .B2(new_n783), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(G1339gat));
  AND2_X1   g591(.A1(new_n641), .A2(new_n644), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n793), .A2(KEYINPUT113), .A3(new_n649), .A4(new_n642), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n645), .B2(new_n646), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n645), .B2(new_n646), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n645), .A2(new_n797), .A3(new_n646), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(new_n655), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n657), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n801), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n564), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n555), .A2(new_n557), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n490), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n550), .A2(new_n491), .A3(new_n553), .A4(new_n558), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n658), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n633), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n806), .A2(new_n657), .A3(new_n802), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n811), .A2(new_n810), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n633), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT114), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n657), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT55), .B1(new_n799), .B2(new_n801), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n633), .A3(new_n816), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n812), .B1(new_n823), .B2(new_n564), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n820), .B(new_n824), .C1(new_n825), .C2(new_n633), .ZN(new_n826));
  INV_X1    g625(.A(new_n704), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n819), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n659), .A2(new_n705), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n334), .A2(new_n399), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n696), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n705), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(new_n285), .ZN(G1340gat));
  NOR3_X1   g635(.A1(new_n834), .A2(new_n283), .A3(new_n706), .ZN(new_n837));
  INV_X1    g636(.A(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n658), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n837), .B1(new_n283), .B2(new_n839), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n834), .B2(new_n827), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n682), .A2(new_n291), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n834), .B2(new_n842), .ZN(G1342gat));
  NOR2_X1   g642(.A1(new_n834), .A2(new_n683), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n296), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n290), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(KEYINPUT56), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(KEYINPUT56), .B2(new_n846), .ZN(G1343gat));
  NAND2_X1  g647(.A1(new_n218), .A2(new_n219), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n716), .A2(new_n832), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n830), .A2(new_n278), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g654(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n856));
  AOI22_X1  g655(.A1(new_n560), .A2(new_n563), .B1(new_n804), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n812), .B1(new_n857), .B2(new_n803), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n633), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(KEYINPUT116), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n824), .B1(new_n859), .B2(KEYINPUT116), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n608), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n829), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n432), .A2(new_n854), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n852), .B1(new_n855), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n850), .B1(new_n866), .B2(new_n564), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n853), .A2(new_n852), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n564), .A2(new_n204), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT117), .Z(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT58), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n830), .B2(new_n278), .ZN(new_n874));
  INV_X1    g673(.A(new_n864), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n862), .B2(new_n829), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n851), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n849), .B1(new_n877), .B2(new_n705), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n879), .A3(new_n871), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n873), .A2(new_n880), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n868), .A2(new_n206), .A3(new_n658), .ZN(new_n882));
  AOI211_X1 g681(.A(KEYINPUT59), .B(new_n206), .C1(new_n866), .C2(new_n658), .ZN(new_n883));
  XNOR2_X1  g682(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n659), .A2(KEYINPUT119), .A3(new_n705), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT119), .B1(new_n659), .B2(new_n705), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n858), .A2(new_n633), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT120), .B1(new_n888), .B2(new_n824), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n824), .B(KEYINPUT120), .C1(new_n858), .C2(new_n633), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n608), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n887), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n892), .B2(new_n278), .ZN(new_n893));
  INV_X1    g692(.A(new_n829), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n813), .B1(new_n815), .B2(new_n705), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n818), .B1(new_n895), .B2(new_n683), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n704), .B1(new_n896), .B2(new_n820), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n894), .B1(new_n897), .B2(new_n819), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n875), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n658), .B(new_n851), .C1(new_n893), .C2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n884), .B1(new_n900), .B2(G148gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n882), .B1(new_n883), .B2(new_n901), .ZN(G1345gat));
  AND3_X1   g701(.A1(new_n866), .A2(G155gat), .A3(new_n704), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n853), .A2(new_n608), .A3(new_n852), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n905));
  AOI21_X1  g704(.A(G155gat), .B1(new_n904), .B2(KEYINPUT121), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(G1346gat));
  AOI21_X1  g706(.A(G162gat), .B1(new_n868), .B2(new_n633), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n633), .A2(G162gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n866), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n661), .A2(new_n400), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n472), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n828), .B2(new_n829), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n564), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(G169gat), .ZN(G1348gat));
  INV_X1    g714(.A(new_n913), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n916), .A2(G176gat), .A3(new_n751), .ZN(new_n917));
  OAI21_X1  g716(.A(G176gat), .B1(new_n916), .B2(new_n706), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1349gat));
  NAND2_X1  g718(.A1(new_n682), .A2(new_n362), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  AOI211_X1 g721(.A(new_n827), .B(new_n912), .C1(new_n828), .C2(new_n829), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n343), .ZN(new_n924));
  XNOR2_X1  g723(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n922), .B(KEYINPUT122), .C1(new_n923), .C2(new_n343), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT123), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n343), .B1(new_n913), .B2(new_n704), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n898), .A2(new_n912), .A3(new_n920), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND4_X1   g733(.A1(KEYINPUT123), .A2(new_n934), .A3(KEYINPUT60), .A4(new_n930), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n926), .B1(new_n931), .B2(new_n935), .ZN(G1350gat));
  OAI22_X1  g735(.A1(new_n916), .A2(new_n683), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(G1351gat));
  OR2_X1    g738(.A1(new_n893), .A2(new_n899), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n468), .A2(new_n911), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT126), .Z(new_n942));
  AND2_X1   g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n705), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n941), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n830), .A2(new_n278), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n564), .A3(new_n950), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n943), .A2(new_n945), .B1(new_n944), .B2(new_n951), .ZN(G1352gat));
  OAI211_X1 g751(.A(new_n707), .B(new_n942), .C1(new_n893), .C2(new_n899), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n751), .A2(G204gat), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n830), .A2(new_n278), .A3(new_n946), .A4(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n954), .A2(KEYINPUT127), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1353gat));
  OAI211_X1 g762(.A(new_n682), .B(new_n946), .C1(new_n893), .C2(new_n899), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n950), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n682), .A2(new_n231), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n965), .A2(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G1354gat));
  NAND3_X1  g768(.A1(new_n940), .A2(new_n633), .A3(new_n942), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G218gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n633), .A2(new_n232), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n967), .B2(new_n972), .ZN(G1355gat));
endmodule


