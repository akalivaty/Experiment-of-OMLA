//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT64), .Z(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(new_n458), .B2(new_n459), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(KEYINPUT66), .A2(G113), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g048(.A(KEYINPUT67), .B(G2105), .C1(new_n465), .C2(new_n470), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n476), .A2(new_n477), .A3(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT3), .B1(new_n476), .B2(new_n477), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n483), .A2(G2104), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G137), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n479), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n475), .A2(new_n489), .ZN(G160));
  NAND3_X1  g065(.A1(new_n480), .A2(new_n485), .A3(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  INV_X1    g068(.A(new_n487), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n486), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n486), .A2(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n480), .A2(new_n485), .A3(G138), .A4(new_n486), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n508), .B(G2104), .C1(G114), .C2(new_n486), .ZN(new_n509));
  INV_X1    g084(.A(G126), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n491), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n507), .A2(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(G543), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n520), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  AND2_X1   g103(.A1(new_n517), .A2(new_n521), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  INV_X1    g105(.A(new_n525), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n530), .A2(new_n532), .A3(new_n533), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n519), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n522), .A2(new_n540), .B1(new_n541), .B2(new_n525), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n519), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n522), .A2(new_n546), .B1(new_n547), .B2(new_n525), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT70), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G188));
  AND3_X1   g131(.A1(new_n517), .A2(G91), .A3(new_n521), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n514), .A2(new_n516), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT72), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G65), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n557), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n519), .A2(KEYINPUT6), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n566), .A2(new_n568), .A3(G53), .A4(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n521), .A2(new_n571), .A3(G53), .A4(G543), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(new_n570), .B2(new_n572), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n565), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  NAND2_X1  g153(.A1(new_n529), .A2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n531), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n517), .A2(KEYINPUT73), .A3(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n558), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G86), .B2(new_n529), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n531), .A2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n519), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n522), .A2(new_n594), .B1(new_n595), .B2(new_n525), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n593), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT72), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT72), .B1(new_n514), .B2(new_n516), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n519), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n531), .A2(G54), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n517), .A2(G92), .A3(new_n521), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT10), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n598), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n486), .ZN(new_n621));
  INV_X1    g196(.A(G135), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n621), .B1(new_n487), .B2(new_n622), .C1(new_n623), .C2(new_n491), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT74), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NOR2_X1   g201(.A1(new_n501), .A2(new_n502), .ZN(new_n627));
  NOR4_X1   g202(.A1(new_n627), .A2(G2105), .A3(new_n477), .A4(new_n476), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT13), .B(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n632), .A3(new_n633), .ZN(G156));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n639), .B2(new_n642), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n643), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n650), .A2(KEYINPUT16), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n645), .B(new_n646), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(new_n643), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT75), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n651), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(KEYINPUT16), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n653), .A2(new_n652), .A3(new_n643), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n637), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n656), .B1(new_n651), .B2(new_n654), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n660), .A3(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n664), .A3(new_n636), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1341), .B(G1348), .Z(new_n667));
  AOI21_X1  g242(.A(new_n635), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n669), .A3(new_n665), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g247(.A1(new_n662), .A2(KEYINPUT78), .A3(new_n669), .A4(new_n665), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  XOR2_X1   g251(.A(G2067), .B(G2678), .Z(new_n677));
  XNOR2_X1  g252(.A(G2084), .B(G2090), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT79), .B(KEYINPUT18), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n677), .B2(new_n678), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT80), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n685), .B(new_n687), .Z(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT20), .Z(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  INV_X1    g271(.A(new_n693), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n690), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n690), .A2(KEYINPUT81), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT82), .B(KEYINPUT83), .Z(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n703), .B(new_n708), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  NAND2_X1  g285(.A1(new_n492), .A2(G119), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n494), .A2(G131), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n486), .A2(G107), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G25), .B(new_n715), .S(G29), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT35), .B(G1991), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G24), .B(G290), .S(G16), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1986), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G23), .ZN(new_n728));
  INV_X1    g303(.A(G288), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT84), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT33), .B(G1976), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n735));
  INV_X1    g310(.A(G22), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G16), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G303), .B2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n737), .B1(new_n739), .B2(new_n735), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G1971), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(G1971), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n730), .A2(KEYINPUT84), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n730), .A2(KEYINPUT84), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n743), .A2(new_n732), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n734), .A2(new_n741), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G6), .B(G305), .S(G16), .Z(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT32), .B(G1981), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n724), .B(new_n726), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n746), .A2(new_n749), .A3(new_n722), .A4(new_n723), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n721), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT87), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(KEYINPUT36), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n753), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G29), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G35), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n498), .B2(G29), .ZN(new_n760));
  MUX2_X1   g335(.A(new_n759), .B(new_n760), .S(KEYINPUT98), .Z(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT29), .Z(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G2090), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n758), .A2(G26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT92), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n492), .A2(G128), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n494), .A2(G140), .ZN(new_n769));
  OR2_X1    g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n486), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n758), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G5), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G171), .B2(G16), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(G1961), .ZN(new_n780));
  NOR2_X1   g355(.A1(G29), .A2(G32), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n478), .A2(G105), .ZN(new_n782));
  INV_X1    g357(.A(G141), .ZN(new_n783));
  INV_X1    g358(.A(G129), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n782), .B1(new_n487), .B2(new_n783), .C1(new_n784), .C2(new_n491), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT94), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT26), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n781), .B1(new_n790), .B2(G29), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT27), .B(G1996), .Z(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n727), .A2(KEYINPUT23), .A3(G20), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT23), .B1(new_n727), .B2(G20), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n794), .B(new_n795), .C1(G299), .C2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1956), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n762), .B2(G2090), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n780), .B(new_n793), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n757), .A2(new_n764), .A3(new_n777), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(G168), .A2(G16), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G16), .B2(G21), .ZN(new_n805));
  INV_X1    g380(.A(G1966), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT88), .B1(G4), .B2(G16), .ZN(new_n808));
  OR3_X1    g383(.A1(KEYINPUT88), .A2(G4), .A3(G16), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n727), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT90), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT89), .B(G1348), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n625), .A2(new_n758), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT95), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n779), .A2(G1961), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT96), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n820));
  NOR2_X1   g395(.A1(KEYINPUT24), .A2(G34), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(KEYINPUT24), .A2(G34), .ZN(new_n823));
  AOI21_X1  g398(.A(G29), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(G160), .A2(G29), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n820), .B2(new_n824), .ZN(new_n826));
  INV_X1    g401(.A(G2084), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n819), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(G27), .A2(G29), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G164), .B2(G29), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT97), .B(G2078), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n817), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n727), .A2(G19), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n549), .B2(new_n727), .ZN(new_n835));
  MUX2_X1   g410(.A(new_n834), .B(new_n835), .S(KEYINPUT91), .Z(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(G1341), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n791), .A2(new_n792), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n815), .A2(new_n833), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G127), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n627), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(G115), .A2(G2104), .ZN(new_n842));
  OAI21_X1  g417(.A(G2105), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n486), .A2(G103), .A3(G2104), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT25), .Z(new_n845));
  INV_X1    g420(.A(G139), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n845), .C1(new_n846), .C2(new_n487), .ZN(new_n847));
  MUX2_X1   g422(.A(G33), .B(new_n847), .S(G29), .Z(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(G2072), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n826), .A2(new_n827), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT30), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(G28), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(G28), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n853), .A3(new_n758), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  NOR4_X1   g430(.A1(new_n803), .A2(new_n807), .A3(new_n839), .A4(new_n855), .ZN(G311));
  INV_X1    g431(.A(new_n803), .ZN(new_n857));
  INV_X1    g432(.A(new_n807), .ZN(new_n858));
  INV_X1    g433(.A(new_n839), .ZN(new_n859));
  INV_X1    g434(.A(new_n855), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n860), .ZN(G150));
  AOI22_X1  g436(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n519), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  INV_X1    g439(.A(G55), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n522), .A2(new_n864), .B1(new_n865), .B2(new_n525), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NOR2_X1   g445(.A1(new_n810), .A2(new_n614), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n549), .ZN(new_n874));
  INV_X1    g449(.A(new_n549), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n873), .B(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n870), .B1(new_n880), .B2(G860), .ZN(G145));
  XNOR2_X1  g456(.A(new_n625), .B(new_n498), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G160), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n492), .A2(G130), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n494), .A2(G142), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n486), .A2(G118), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n715), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n629), .B(new_n847), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n772), .B(G164), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n790), .ZN(new_n894));
  INV_X1    g469(.A(new_n892), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n629), .B(new_n847), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n890), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n893), .A2(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n790), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n897), .A3(new_n894), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n889), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n883), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n900), .A2(new_n904), .A3(new_n883), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n900), .A2(new_n904), .ZN(new_n913));
  INV_X1    g488(.A(new_n883), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n906), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n905), .A2(KEYINPUT102), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n911), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT103), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(G395));
  NOR2_X1   g497(.A1(new_n868), .A2(G868), .ZN(new_n923));
  XOR2_X1   g498(.A(G303), .B(G290), .Z(new_n924));
  XNOR2_X1  g499(.A(G305), .B(new_n729), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT42), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n607), .A2(G299), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n810), .A2(new_n611), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT105), .B1(new_n810), .B2(new_n611), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n930), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n616), .B(new_n877), .Z(new_n939));
  OAI22_X1  g514(.A1(new_n929), .A2(KEYINPUT106), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n933), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n923), .B1(new_n944), .B2(G868), .ZN(G295));
  AOI21_X1  g520(.A(new_n923), .B1(new_n944), .B2(G868), .ZN(G331));
  XOR2_X1   g521(.A(G171), .B(G286), .Z(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(new_n877), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n941), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT108), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n941), .A2(KEYINPUT41), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n934), .A2(new_n935), .ZN(new_n952));
  AOI211_X1 g527(.A(new_n948), .B(new_n951), .C1(new_n952), .C2(KEYINPUT41), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n926), .B(new_n927), .C1(new_n950), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n928), .B(new_n949), .C1(new_n938), .C2(new_n948), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n910), .A4(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n948), .B1(new_n936), .B2(new_n937), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n928), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(new_n949), .ZN(new_n960));
  OR3_X1    g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n910), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n955), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n954), .A2(new_n910), .A3(new_n956), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(new_n967), .B2(new_n955), .ZN(new_n968));
  MUX2_X1   g543(.A(new_n965), .B(new_n968), .S(KEYINPUT44), .Z(G397));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n507), .B2(new_n511), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  OAI211_X1 g549(.A(KEYINPUT109), .B(new_n970), .C1(new_n507), .C2(new_n511), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n475), .A2(new_n978), .A3(new_n489), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT110), .B1(new_n980), .B2(G1996), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n980), .A2(KEYINPUT110), .A3(G1996), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(new_n894), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n772), .B(G2067), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT111), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n894), .A2(G1996), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n980), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR4_X1   g565(.A1(new_n986), .A2(new_n717), .A3(new_n715), .A4(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n772), .A2(G2067), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n981), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n986), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n715), .B(new_n717), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n981), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n990), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n980), .A2(G1986), .A3(G290), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n998), .B(KEYINPUT48), .Z(new_n999));
  NAND4_X1  g574(.A1(new_n994), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n988), .A2(new_n790), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n1001), .A2(new_n980), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n985), .A2(KEYINPUT125), .A3(KEYINPUT46), .ZN(new_n1003));
  NAND2_X1  g578(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n983), .B2(new_n984), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n993), .B(new_n1000), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n565), .A2(new_n576), .A3(KEYINPUT57), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT117), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n565), .A2(new_n576), .A3(new_n1014), .A4(KEYINPUT57), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n519), .B1(new_n562), .B2(new_n563), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n570), .A2(new_n572), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1017), .A2(new_n557), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT116), .B1(new_n1019), .B2(KEYINPUT57), .ZN(new_n1020));
  INV_X1    g595(.A(new_n557), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n570), .A2(new_n572), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n601), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n1022), .C1(new_n1023), .C2(new_n519), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1016), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1031), .B(new_n970), .C1(new_n507), .C2(new_n511), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n979), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n797), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n971), .A2(new_n974), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT45), .B(new_n970), .C1(new_n507), .C2(new_n511), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT56), .B(G2072), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1035), .A2(new_n979), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1029), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1033), .A2(new_n814), .ZN(new_n1040));
  INV_X1    g615(.A(new_n971), .ZN(new_n1041));
  INV_X1    g616(.A(G2067), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n979), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n607), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1029), .A2(KEYINPUT118), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1013), .A2(new_n1015), .B1(new_n1020), .B2(new_n1027), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1045), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(KEYINPUT120), .A3(new_n1047), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1039), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT120), .B1(new_n1050), .B2(new_n1047), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n607), .A2(KEYINPUT121), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1044), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n607), .A2(KEYINPUT121), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(new_n1040), .A3(KEYINPUT60), .A4(new_n1043), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1044), .A2(new_n1059), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1060), .A2(new_n1062), .B1(new_n1063), .B2(new_n1058), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1051), .A2(KEYINPUT61), .A3(new_n1039), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1035), .A2(new_n979), .A3(new_n1036), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(G1996), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(KEYINPUT119), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1068), .A2(new_n1071), .A3(G1996), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT58), .B(G1341), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n979), .B2(new_n1041), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1067), .B1(new_n1075), .B2(new_n875), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1069), .B(KEYINPUT119), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT59), .B(new_n549), .C1(new_n1077), .C2(new_n1074), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1052), .B1(new_n1066), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1961), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1033), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1035), .A2(new_n979), .A3(new_n1084), .A4(new_n1036), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1082), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1083), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1082), .B(KEYINPUT122), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1088), .A2(G301), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n489), .A2(G2078), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n471), .A2(KEYINPUT53), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n976), .A2(new_n1036), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1089), .B(new_n1082), .C1(new_n1095), .C2(new_n978), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1096), .B2(G171), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1091), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G303), .A2(G8), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT55), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT112), .B(G1971), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1068), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1030), .A2(new_n979), .A3(new_n1032), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n1105));
  AOI21_X1  g680(.A(G2090), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1103), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G8), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1100), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n1033), .A2(new_n1111), .A3(G2090), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1033), .B2(G2090), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1102), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1100), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(G8), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT49), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n589), .A2(new_n1118), .A3(new_n590), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n588), .A2(G651), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT114), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G1981), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1109), .B1(new_n979), .B2(new_n1041), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1117), .A2(G1981), .A3(new_n1122), .A4(new_n1119), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n729), .A2(G1976), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT52), .ZN(new_n1130));
  INV_X1    g705(.A(G1976), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT52), .B1(G288), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1125), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1127), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1110), .A2(new_n1116), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1068), .A2(new_n806), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1138), .B(G168), .C1(G2084), .C2(new_n1033), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1139), .B2(G8), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1104), .A2(new_n827), .B1(new_n1068), .B2(new_n806), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1109), .B1(new_n1141), .B2(G168), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT51), .B1(new_n1141), .B2(G168), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1098), .A2(new_n1136), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1096), .A2(G171), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n1147), .B2(G171), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT123), .B1(new_n1148), .B2(KEYINPUT54), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1147), .A2(G171), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1150), .B(new_n1092), .C1(new_n1152), .C2(new_n1146), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1080), .A2(new_n1145), .A3(new_n1149), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1127), .A2(new_n1131), .A3(new_n729), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(G1981), .B2(G305), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1125), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1116), .B2(new_n1134), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1141), .A2(new_n1109), .A3(G286), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1136), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1114), .A2(G8), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1163), .B2(new_n1100), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1164), .A2(new_n1116), .A3(new_n1135), .A4(new_n1160), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1158), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1154), .A2(KEYINPUT124), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT124), .B1(new_n1154), .B2(new_n1166), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1144), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1169), .A2(KEYINPUT62), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(KEYINPUT62), .ZN(new_n1171));
  NOR4_X1   g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n1151), .A4(new_n1136), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1167), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(G290), .B(G1986), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n981), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n994), .A2(new_n1175), .A3(new_n996), .A4(new_n997), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1011), .B1(new_n1173), .B2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1179));
  INV_X1    g753(.A(G227), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n674), .A2(G319), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g757(.A1(new_n674), .A2(KEYINPUT126), .A3(G319), .A4(new_n1180), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1179), .B1(new_n1185), .B2(new_n709), .ZN(new_n1186));
  AOI211_X1 g760(.A(KEYINPUT127), .B(G229), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n908), .B1(new_n907), .B2(new_n911), .ZN(new_n1188));
  AND4_X1   g762(.A1(new_n908), .A2(new_n916), .A3(new_n911), .A4(new_n917), .ZN(new_n1189));
  OAI21_X1  g763(.A(new_n965), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g764(.A1(new_n1186), .A2(new_n1187), .A3(new_n1190), .ZN(G308));
  NAND2_X1  g765(.A1(new_n1185), .A2(new_n709), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1192), .A2(KEYINPUT127), .ZN(new_n1193));
  INV_X1    g767(.A(new_n1190), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n1185), .A2(new_n1179), .A3(new_n709), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(G225));
endmodule


