

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U326 ( .A(n364), .B(n363), .ZN(n365) );
  INV_X1 U327 ( .A(KEYINPUT23), .ZN(n363) );
  INV_X1 U328 ( .A(KEYINPUT103), .ZN(n416) );
  AND2_X1 U329 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  AND2_X1 U330 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U331 ( .A(n398), .B(n443), .ZN(n296) );
  XNOR2_X1 U332 ( .A(n357), .B(n295), .ZN(n358) );
  XNOR2_X1 U333 ( .A(n387), .B(n358), .ZN(n360) );
  INV_X1 U334 ( .A(KEYINPUT94), .ZN(n390) );
  XNOR2_X1 U335 ( .A(n441), .B(n294), .ZN(n442) );
  XNOR2_X1 U336 ( .A(n465), .B(KEYINPUT47), .ZN(n466) );
  XNOR2_X1 U337 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U338 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U339 ( .A(n467), .B(n466), .ZN(n472) );
  XNOR2_X1 U340 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U341 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U342 ( .A(n416), .B(KEYINPUT37), .ZN(n417) );
  XNOR2_X1 U343 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U344 ( .A(n455), .B(n454), .ZN(n460) );
  XOR2_X1 U345 ( .A(n436), .B(n435), .Z(n552) );
  INV_X1 U346 ( .A(G43GAT), .ZN(n483) );
  XNOR2_X1 U347 ( .A(KEYINPUT38), .B(n456), .ZN(n506) );
  XNOR2_X1 U348 ( .A(n480), .B(KEYINPUT124), .ZN(n481) );
  XNOR2_X1 U349 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U350 ( .A(n482), .B(n481), .ZN(G1350GAT) );
  XNOR2_X1 U351 ( .A(n486), .B(n485), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT0), .B(G127GAT), .Z(n298) );
  XNOR2_X1 U353 ( .A(KEYINPUT81), .B(G120GAT), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U355 ( .A(G113GAT), .B(n299), .Z(n373) );
  XNOR2_X1 U356 ( .A(G134GAT), .B(G162GAT), .ZN(n300) );
  XOR2_X1 U357 ( .A(G148GAT), .B(G57GAT), .Z(n437) );
  XNOR2_X1 U358 ( .A(n300), .B(n437), .ZN(n304) );
  XOR2_X1 U359 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n302) );
  XNOR2_X1 U360 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U362 ( .A(n304), .B(n303), .Z(n314) );
  XOR2_X1 U363 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n306) );
  XNOR2_X1 U364 ( .A(KEYINPUT90), .B(KEYINPUT92), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n306), .B(n305), .ZN(n312) );
  XOR2_X1 U366 ( .A(G29GAT), .B(G85GAT), .Z(n321) );
  XOR2_X1 U367 ( .A(G155GAT), .B(KEYINPUT2), .Z(n308) );
  XNOR2_X1 U368 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n359) );
  XOR2_X1 U370 ( .A(n321), .B(n359), .Z(n310) );
  NAND2_X1 U371 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U372 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n373), .B(n315), .ZN(n406) );
  XNOR2_X1 U376 ( .A(KEYINPUT93), .B(n406), .ZN(n523) );
  XOR2_X1 U377 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n317) );
  XNOR2_X1 U378 ( .A(G218GAT), .B(G92GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U380 ( .A(n318), .B(KEYINPUT77), .Z(n320) );
  XOR2_X1 U381 ( .A(G43GAT), .B(G134GAT), .Z(n369) );
  XNOR2_X1 U382 ( .A(G36GAT), .B(n369), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n322) );
  XOR2_X1 U384 ( .A(n322), .B(n321), .Z(n325) );
  XNOR2_X1 U385 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n323), .B(KEYINPUT69), .ZN(n432) );
  XOR2_X1 U387 ( .A(G50GAT), .B(G162GAT), .Z(n357) );
  XNOR2_X1 U388 ( .A(n432), .B(n357), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U390 ( .A(G106GAT), .B(G99GAT), .Z(n327) );
  NAND2_X1 U391 ( .A1(G232GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U393 ( .A(n329), .B(n328), .Z(n334) );
  XOR2_X1 U394 ( .A(KEYINPUT65), .B(KEYINPUT76), .Z(n331) );
  XNOR2_X1 U395 ( .A(KEYINPUT10), .B(KEYINPUT64), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U397 ( .A(G190GAT), .B(n332), .ZN(n333) );
  XOR2_X1 U398 ( .A(n334), .B(n333), .Z(n571) );
  INV_X1 U399 ( .A(n571), .ZN(n560) );
  XOR2_X1 U400 ( .A(KEYINPUT36), .B(n560), .Z(n586) );
  XOR2_X1 U401 ( .A(G211GAT), .B(G155GAT), .Z(n336) );
  XNOR2_X1 U402 ( .A(G127GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U404 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n438) );
  XOR2_X1 U405 ( .A(n337), .B(n438), .Z(n339) );
  XNOR2_X1 U406 ( .A(G183GAT), .B(G71GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n344) );
  XNOR2_X1 U408 ( .A(G15GAT), .B(G22GAT), .ZN(n340) );
  XNOR2_X1 U409 ( .A(n340), .B(G1GAT), .ZN(n431) );
  XOR2_X1 U410 ( .A(n431), .B(KEYINPUT14), .Z(n342) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U412 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U413 ( .A(n344), .B(n343), .Z(n352) );
  XOR2_X1 U414 ( .A(KEYINPUT78), .B(G64GAT), .Z(n346) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(G57GAT), .ZN(n345) );
  XNOR2_X1 U416 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U417 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n348) );
  XNOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n347) );
  XNOR2_X1 U419 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U420 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U421 ( .A(n352), .B(n351), .Z(n558) );
  INV_X1 U422 ( .A(n558), .ZN(n583) );
  XOR2_X1 U423 ( .A(KEYINPUT22), .B(G148GAT), .Z(n354) );
  XNOR2_X1 U424 ( .A(G22GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U425 ( .A(n354), .B(n353), .ZN(n368) );
  XOR2_X1 U426 ( .A(G211GAT), .B(KEYINPUT21), .Z(n356) );
  XNOR2_X1 U427 ( .A(G197GAT), .B(G218GAT), .ZN(n355) );
  XNOR2_X1 U428 ( .A(n356), .B(n355), .ZN(n387) );
  XOR2_X1 U429 ( .A(n360), .B(n359), .Z(n362) );
  XNOR2_X1 U430 ( .A(KEYINPUT89), .B(KEYINPUT24), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U432 ( .A(G106GAT), .B(G78GAT), .Z(n449) );
  XNOR2_X1 U433 ( .A(n449), .B(KEYINPUT88), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n477) );
  XOR2_X1 U435 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n371) );
  XOR2_X1 U436 ( .A(G99GAT), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U437 ( .A(n369), .B(n441), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U439 ( .A(n372), .B(KEYINPUT86), .Z(n375) );
  XNOR2_X1 U440 ( .A(G15GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U442 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n377) );
  NAND2_X1 U443 ( .A1(G227GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U445 ( .A(n379), .B(n378), .Z(n386) );
  XOR2_X1 U446 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n381) );
  XNOR2_X1 U447 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U449 ( .A(n382), .B(G183GAT), .Z(n384) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(G176GAT), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n384), .B(n383), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n395), .B(KEYINPUT20), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n534) );
  XOR2_X1 U454 ( .A(n387), .B(KEYINPUT95), .Z(n389) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U457 ( .A(G36GAT), .B(G8GAT), .Z(n424) );
  XNOR2_X1 U458 ( .A(n424), .B(KEYINPUT78), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n398) );
  XNOR2_X1 U460 ( .A(G92GAT), .B(KEYINPUT72), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n396), .B(G64GAT), .ZN(n397) );
  XOR2_X1 U462 ( .A(G204GAT), .B(n397), .Z(n443) );
  NAND2_X1 U463 ( .A1(n534), .A2(n296), .ZN(n399) );
  NAND2_X1 U464 ( .A1(n477), .A2(n399), .ZN(n400) );
  XNOR2_X1 U465 ( .A(KEYINPUT25), .B(n400), .ZN(n404) );
  NOR2_X1 U466 ( .A1(n477), .A2(n534), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n401), .B(KEYINPUT26), .ZN(n574) );
  XNOR2_X1 U468 ( .A(KEYINPUT27), .B(n296), .ZN(n408) );
  NAND2_X1 U469 ( .A1(n574), .A2(n408), .ZN(n402) );
  XOR2_X1 U470 ( .A(KEYINPUT98), .B(n402), .Z(n403) );
  NOR2_X1 U471 ( .A1(n404), .A2(n403), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n405), .B(KEYINPUT99), .ZN(n407) );
  NAND2_X1 U473 ( .A1(n407), .A2(n406), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n534), .B(KEYINPUT87), .ZN(n412) );
  XOR2_X1 U475 ( .A(KEYINPUT28), .B(n477), .Z(n527) );
  INV_X1 U476 ( .A(n527), .ZN(n410) );
  NAND2_X1 U477 ( .A1(n408), .A2(n523), .ZN(n409) );
  XOR2_X1 U478 ( .A(KEYINPUT96), .B(n409), .Z(n549) );
  NAND2_X1 U479 ( .A1(n410), .A2(n549), .ZN(n533) );
  XNOR2_X1 U480 ( .A(n533), .B(KEYINPUT97), .ZN(n411) );
  NAND2_X1 U481 ( .A1(n412), .A2(n411), .ZN(n413) );
  NAND2_X1 U482 ( .A1(n414), .A2(n413), .ZN(n491) );
  NAND2_X1 U483 ( .A1(n583), .A2(n491), .ZN(n415) );
  NOR2_X1 U484 ( .A1(n586), .A2(n415), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n522) );
  XOR2_X1 U486 ( .A(KEYINPUT68), .B(G197GAT), .Z(n420) );
  XNOR2_X1 U487 ( .A(G113GAT), .B(G141GAT), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n436) );
  XOR2_X1 U489 ( .A(G43GAT), .B(G29GAT), .Z(n422) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(G50GAT), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U492 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U494 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U495 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n428) );
  XNOR2_X1 U496 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n427) );
  XNOR2_X1 U497 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U498 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U501 ( .A(n438), .B(n437), .Z(n440) );
  XNOR2_X1 U502 ( .A(G176GAT), .B(G85GAT), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n455) );
  XOR2_X1 U505 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n447) );
  XNOR2_X1 U506 ( .A(KEYINPUT31), .B(KEYINPUT71), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U508 ( .A(n449), .B(n448), .Z(n453) );
  XOR2_X1 U509 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n451) );
  XNOR2_X1 U510 ( .A(G120GAT), .B(KEYINPUT75), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U512 ( .A1(n552), .A2(n460), .ZN(n493) );
  NOR2_X1 U513 ( .A1(n522), .A2(n493), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n523), .A2(n506), .ZN(n459) );
  XOR2_X1 U515 ( .A(G29GAT), .B(KEYINPUT104), .Z(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT39), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(G1328GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT41), .B(n460), .Z(n563) );
  INV_X1 U519 ( .A(n563), .ZN(n540) );
  NAND2_X1 U520 ( .A1(n540), .A2(n552), .ZN(n461) );
  XNOR2_X1 U521 ( .A(KEYINPUT46), .B(n461), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n462), .A2(n583), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT114), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n560), .A2(n464), .ZN(n467) );
  XNOR2_X1 U525 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n586), .A2(n583), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT45), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n469), .A2(n460), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n470), .A2(n552), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT48), .B(n473), .ZN(n551) );
  INV_X1 U532 ( .A(n551), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n474), .A2(n296), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT54), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n523), .A2(n476), .ZN(n575) );
  NAND2_X1 U536 ( .A1(n575), .A2(n477), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(KEYINPUT55), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n479), .A2(n534), .ZN(n570) );
  NOR2_X1 U539 ( .A1(n583), .A2(n570), .ZN(n482) );
  INV_X1 U540 ( .A(G183GAT), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n534), .A2(n506), .ZN(n486) );
  XOR2_X1 U542 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n484) );
  INV_X1 U543 ( .A(n552), .ZN(n576) );
  NOR2_X1 U544 ( .A1(n576), .A2(n570), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT122), .ZN(n489) );
  INV_X1 U546 ( .A(G169GAT), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1348GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n495) );
  NOR2_X1 U549 ( .A1(n560), .A2(n583), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT16), .ZN(n492) );
  NAND2_X1 U551 ( .A1(n492), .A2(n491), .ZN(n510) );
  NOR2_X1 U552 ( .A1(n493), .A2(n510), .ZN(n501) );
  NAND2_X1 U553 ( .A1(n501), .A2(n523), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U555 ( .A(G1GAT), .B(n496), .Z(G1324GAT) );
  NAND2_X1 U556 ( .A1(n501), .A2(n296), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U559 ( .A1(n501), .A2(n534), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U561 ( .A(G15GAT), .B(n500), .Z(G1326GAT) );
  NAND2_X1 U562 ( .A1(n527), .A2(n501), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT102), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  XOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT105), .Z(n505) );
  NAND2_X1 U566 ( .A1(n296), .A2(n506), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1329GAT) );
  XOR2_X1 U568 ( .A(G50GAT), .B(KEYINPUT107), .Z(n508) );
  NAND2_X1 U569 ( .A1(n506), .A2(n527), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n512) );
  NOR2_X1 U572 ( .A1(n563), .A2(n552), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT109), .ZN(n521) );
  NOR2_X1 U574 ( .A1(n521), .A2(n510), .ZN(n516) );
  NAND2_X1 U575 ( .A1(n516), .A2(n523), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U577 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NAND2_X1 U578 ( .A1(n516), .A2(n296), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n534), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U583 ( .A1(n516), .A2(n527), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT110), .Z(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n523), .A2(n528), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n296), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n534), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n530) );
  NAND2_X1 U596 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1339GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n538) );
  NOR2_X1 U600 ( .A1(n551), .A2(n533), .ZN(n535) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(KEYINPUT117), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n546), .A2(n552), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U607 ( .A1(n546), .A2(n540), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n544) );
  NAND2_X1 U610 ( .A1(n546), .A2(n558), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n545), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n560), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n574), .A2(n549), .ZN(n550) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n561), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U621 ( .A1(n561), .A2(n540), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n561), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n570), .A2(n563), .ZN(n567) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n565) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n569) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT126), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n573) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(n573), .B(n572), .Z(G1351GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n585) );
  NOR2_X1 U640 ( .A1(n576), .A2(n585), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n460), .A2(n585), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

