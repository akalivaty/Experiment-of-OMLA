

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(n818), .A2(n817), .ZN(n521) );
  NOR2_X1 U554 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U555 ( .A1(n798), .A2(n799), .ZN(n809) );
  NOR2_X1 U556 ( .A1(n963), .A2(n753), .ZN(n741) );
  NAND2_X1 U557 ( .A1(n729), .A2(n728), .ZN(n788) );
  XNOR2_X1 U558 ( .A(n553), .B(KEYINPUT91), .ZN(G164) );
  NAND2_X1 U559 ( .A1(n809), .A2(n808), .ZN(n810) );
  AND2_X1 U560 ( .A1(n783), .A2(n782), .ZN(n519) );
  AND2_X1 U561 ( .A1(n821), .A2(n820), .ZN(n520) );
  XNOR2_X1 U562 ( .A(n735), .B(n734), .ZN(n737) );
  INV_X1 U563 ( .A(KEYINPUT99), .ZN(n768) );
  INV_X1 U564 ( .A(KEYINPUT28), .ZN(n740) );
  INV_X1 U565 ( .A(KEYINPUT31), .ZN(n776) );
  AND2_X1 U566 ( .A1(n787), .A2(n519), .ZN(n785) );
  NAND2_X1 U567 ( .A1(G8), .A2(n788), .ZN(n815) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  AND2_X1 U569 ( .A1(n822), .A2(n520), .ZN(n823) );
  XNOR2_X1 U570 ( .A(G543), .B(KEYINPUT0), .ZN(n535) );
  NOR2_X1 U571 ( .A1(n542), .A2(n644), .ZN(n655) );
  NOR2_X1 U572 ( .A1(G2105), .A2(n528), .ZN(n615) );
  BUF_X1 U573 ( .A(n525), .Z(n890) );
  NAND2_X1 U574 ( .A1(n579), .A2(n578), .ZN(n972) );
  NOR2_X1 U575 ( .A1(n532), .A2(n531), .ZN(G160) );
  INV_X1 U576 ( .A(G2104), .ZN(n528) );
  NAND2_X1 U577 ( .A1(G101), .A2(n615), .ZN(n522) );
  XNOR2_X1 U578 ( .A(n522), .B(KEYINPUT23), .ZN(n523) );
  XNOR2_X1 U579 ( .A(n523), .B(KEYINPUT65), .ZN(n527) );
  XOR2_X1 U580 ( .A(KEYINPUT17), .B(n524), .Z(n525) );
  NAND2_X1 U581 ( .A1(G137), .A2(n890), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n532) );
  AND2_X1 U583 ( .A1(n528), .A2(G2105), .ZN(n886) );
  NAND2_X1 U584 ( .A1(G125), .A2(n886), .ZN(n530) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n887) );
  NAND2_X1 U586 ( .A1(G113), .A2(n887), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U588 ( .A1(G543), .A2(G651), .ZN(n533) );
  XNOR2_X1 U589 ( .A(n533), .B(KEYINPUT64), .ZN(n656) );
  NAND2_X1 U590 ( .A1(G90), .A2(n656), .ZN(n534) );
  XNOR2_X1 U591 ( .A(n534), .B(KEYINPUT68), .ZN(n538) );
  INV_X1 U592 ( .A(G651), .ZN(n542) );
  INV_X1 U593 ( .A(n535), .ZN(n536) );
  XNOR2_X1 U594 ( .A(KEYINPUT66), .B(n536), .ZN(n644) );
  NAND2_X1 U595 ( .A1(G77), .A2(n655), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U597 ( .A(n539), .B(KEYINPUT9), .ZN(n541) );
  NOR2_X2 U598 ( .A1(G651), .A2(n644), .ZN(n661) );
  NAND2_X1 U599 ( .A1(G52), .A2(n661), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n541), .A2(n540), .ZN(n546) );
  NOR2_X1 U601 ( .A1(G543), .A2(n542), .ZN(n543) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n543), .Z(n654) );
  NAND2_X1 U603 ( .A1(G64), .A2(n654), .ZN(n544) );
  XNOR2_X1 U604 ( .A(KEYINPUT67), .B(n544), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n546), .A2(n545), .ZN(G171) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U607 ( .A(G57), .ZN(G237) );
  INV_X1 U608 ( .A(G69), .ZN(G235) );
  INV_X1 U609 ( .A(G108), .ZN(G238) );
  INV_X1 U610 ( .A(G120), .ZN(G236) );
  NAND2_X1 U611 ( .A1(n525), .A2(G138), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G114), .A2(n887), .ZN(n548) );
  NAND2_X1 U613 ( .A1(G102), .A2(n615), .ZN(n547) );
  AND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U615 ( .A1(G126), .A2(n886), .ZN(n549) );
  AND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U618 ( .A1(G89), .A2(n656), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  NAND2_X1 U620 ( .A1(G76), .A2(n655), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT5), .B(n557), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n661), .A2(G51), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT75), .B(n558), .Z(n560) );
  NAND2_X1 U625 ( .A1(n654), .A2(G63), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT6), .B(n561), .Z(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT10), .ZN(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT70), .B(n566), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n829) );
  NAND2_X1 U635 ( .A1(n829), .A2(G567), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n567), .B(KEYINPUT71), .ZN(n568) );
  XNOR2_X1 U637 ( .A(KEYINPUT11), .B(n568), .ZN(G234) );
  NAND2_X1 U638 ( .A1(G56), .A2(n654), .ZN(n569) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n569), .Z(n577) );
  NAND2_X1 U640 ( .A1(G81), .A2(n656), .ZN(n570) );
  XOR2_X1 U641 ( .A(KEYINPUT12), .B(n570), .Z(n574) );
  NAND2_X1 U642 ( .A1(n655), .A2(G68), .ZN(n571) );
  XNOR2_X1 U643 ( .A(KEYINPUT72), .B(n571), .ZN(n572) );
  INV_X1 U644 ( .A(n572), .ZN(n573) );
  NOR2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U646 ( .A(n575), .B(KEYINPUT13), .ZN(n576) );
  NOR2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n661), .A2(G43), .ZN(n578) );
  INV_X1 U649 ( .A(G860), .ZN(n603) );
  OR2_X1 U650 ( .A1(n972), .A2(n603), .ZN(G153) );
  XNOR2_X1 U651 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n655), .A2(G79), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G66), .A2(n654), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G92), .A2(n656), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n661), .A2(G54), .ZN(n582) );
  XOR2_X1 U658 ( .A(KEYINPUT74), .B(n582), .Z(n583) );
  NOR2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U661 ( .A(KEYINPUT15), .B(n587), .Z(n956) );
  INV_X1 U662 ( .A(G868), .ZN(n673) );
  NAND2_X1 U663 ( .A1(n956), .A2(n673), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U665 ( .A1(G65), .A2(n654), .ZN(n591) );
  NAND2_X1 U666 ( .A1(G78), .A2(n655), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U668 ( .A1(G91), .A2(n656), .ZN(n592) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n592), .ZN(n593) );
  NOR2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n661), .A2(G53), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(G299) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n597) );
  XOR2_X1 U674 ( .A(KEYINPUT78), .B(n597), .Z(n601) );
  XOR2_X1 U675 ( .A(G868), .B(KEYINPUT76), .Z(n598) );
  NOR2_X1 U676 ( .A1(G286), .A2(n598), .ZN(n599) );
  XNOR2_X1 U677 ( .A(KEYINPUT77), .B(n599), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U679 ( .A(KEYINPUT79), .B(n602), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U681 ( .A(n956), .ZN(n622) );
  NAND2_X1 U682 ( .A1(n604), .A2(n622), .ZN(n605) );
  XNOR2_X1 U683 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U684 ( .A1(n622), .A2(G868), .ZN(n606) );
  NOR2_X1 U685 ( .A1(G559), .A2(n606), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n607), .B(KEYINPUT80), .ZN(n609) );
  NOR2_X1 U687 ( .A1(n972), .A2(G868), .ZN(n608) );
  NOR2_X1 U688 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U689 ( .A1(G123), .A2(n886), .ZN(n610) );
  XOR2_X1 U690 ( .A(KEYINPUT18), .B(n610), .Z(n611) );
  XNOR2_X1 U691 ( .A(n611), .B(KEYINPUT81), .ZN(n613) );
  NAND2_X1 U692 ( .A1(G135), .A2(n890), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U694 ( .A(KEYINPUT82), .B(n614), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G111), .A2(n887), .ZN(n617) );
  BUF_X1 U696 ( .A(n615), .Z(n891) );
  NAND2_X1 U697 ( .A1(G99), .A2(n891), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n932) );
  XNOR2_X1 U700 ( .A(n932), .B(G2096), .ZN(n621) );
  INV_X1 U701 ( .A(G2100), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(G156) );
  NAND2_X1 U703 ( .A1(n622), .A2(G559), .ZN(n670) );
  XOR2_X1 U704 ( .A(KEYINPUT83), .B(n972), .Z(n623) );
  XNOR2_X1 U705 ( .A(n670), .B(n623), .ZN(n624) );
  NOR2_X1 U706 ( .A1(G860), .A2(n624), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G67), .A2(n654), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G55), .A2(n661), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U710 ( .A(KEYINPUT85), .B(n627), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G80), .A2(n655), .ZN(n629) );
  NAND2_X1 U712 ( .A1(G93), .A2(n656), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U714 ( .A(KEYINPUT84), .B(n630), .Z(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n672) );
  XOR2_X1 U716 ( .A(n633), .B(n672), .Z(G145) );
  NAND2_X1 U717 ( .A1(G75), .A2(n655), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G88), .A2(n656), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U720 ( .A(KEYINPUT86), .B(n636), .Z(n640) );
  NAND2_X1 U721 ( .A1(G62), .A2(n654), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G50), .A2(n661), .ZN(n637) );
  AND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(G303) );
  INV_X1 U725 ( .A(G303), .ZN(G166) );
  NAND2_X1 U726 ( .A1(G49), .A2(n661), .ZN(n642) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U729 ( .A1(n654), .A2(n643), .ZN(n646) );
  NAND2_X1 U730 ( .A1(G87), .A2(n644), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U732 ( .A1(G61), .A2(n654), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G86), .A2(n656), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n655), .A2(G73), .ZN(n649) );
  XOR2_X1 U736 ( .A(KEYINPUT2), .B(n649), .Z(n650) );
  NOR2_X1 U737 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U738 ( .A1(n661), .A2(G48), .ZN(n652) );
  NAND2_X1 U739 ( .A1(n653), .A2(n652), .ZN(G305) );
  AND2_X1 U740 ( .A1(n654), .A2(G60), .ZN(n660) );
  NAND2_X1 U741 ( .A1(G72), .A2(n655), .ZN(n658) );
  NAND2_X1 U742 ( .A1(G85), .A2(n656), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U745 ( .A1(n661), .A2(G47), .ZN(n662) );
  NAND2_X1 U746 ( .A1(n663), .A2(n662), .ZN(G290) );
  XNOR2_X1 U747 ( .A(KEYINPUT19), .B(G288), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n664), .B(G305), .ZN(n665) );
  XNOR2_X1 U749 ( .A(G166), .B(n665), .ZN(n667) );
  INV_X1 U750 ( .A(G299), .ZN(n963) );
  XNOR2_X1 U751 ( .A(G290), .B(n963), .ZN(n666) );
  XNOR2_X1 U752 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U753 ( .A(n668), .B(n972), .ZN(n669) );
  XNOR2_X1 U754 ( .A(n669), .B(n672), .ZN(n903) );
  XOR2_X1 U755 ( .A(n903), .B(n670), .Z(n671) );
  NAND2_X1 U756 ( .A1(G868), .A2(n671), .ZN(n675) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XNOR2_X1 U760 ( .A(n676), .B(KEYINPUT20), .ZN(n677) );
  XNOR2_X1 U761 ( .A(n677), .B(KEYINPUT87), .ZN(n678) );
  NAND2_X1 U762 ( .A1(n678), .A2(G2090), .ZN(n679) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n682) );
  NAND2_X1 U767 ( .A1(G132), .A2(G82), .ZN(n681) );
  XNOR2_X1 U768 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U769 ( .A(n683), .B(KEYINPUT88), .ZN(n684) );
  NOR2_X1 U770 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U771 ( .A1(G96), .A2(n685), .ZN(n833) );
  NAND2_X1 U772 ( .A1(n833), .A2(G2106), .ZN(n690) );
  NOR2_X1 U773 ( .A1(G236), .A2(G238), .ZN(n687) );
  NOR2_X1 U774 ( .A1(G235), .A2(G237), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U776 ( .A(KEYINPUT90), .B(n688), .ZN(n834) );
  NAND2_X1 U777 ( .A1(n834), .A2(G567), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n835) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n691) );
  NOR2_X1 U780 ( .A1(n835), .A2(n691), .ZN(n832) );
  NAND2_X1 U781 ( .A1(n832), .A2(G36), .ZN(G176) );
  NAND2_X1 U782 ( .A1(G105), .A2(n891), .ZN(n692) );
  XNOR2_X1 U783 ( .A(n692), .B(KEYINPUT38), .ZN(n699) );
  NAND2_X1 U784 ( .A1(G141), .A2(n890), .ZN(n694) );
  NAND2_X1 U785 ( .A1(G117), .A2(n887), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U787 ( .A1(G129), .A2(n886), .ZN(n695) );
  XNOR2_X1 U788 ( .A(KEYINPUT93), .B(n695), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n871) );
  NOR2_X1 U791 ( .A1(G1996), .A2(n871), .ZN(n927) );
  NOR2_X1 U792 ( .A1(G164), .A2(G1384), .ZN(n728) );
  NAND2_X1 U793 ( .A1(G160), .A2(G40), .ZN(n727) );
  NOR2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n819) );
  NAND2_X1 U795 ( .A1(G119), .A2(n886), .ZN(n701) );
  NAND2_X1 U796 ( .A1(G131), .A2(n890), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n705) );
  NAND2_X1 U798 ( .A1(G107), .A2(n887), .ZN(n703) );
  NAND2_X1 U799 ( .A1(G95), .A2(n891), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n704) );
  OR2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n867) );
  NAND2_X1 U802 ( .A1(G1991), .A2(n867), .ZN(n707) );
  NAND2_X1 U803 ( .A1(G1996), .A2(n871), .ZN(n706) );
  NAND2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n923) );
  NAND2_X1 U805 ( .A1(n819), .A2(n923), .ZN(n821) );
  INV_X1 U806 ( .A(n821), .ZN(n710) );
  NOR2_X1 U807 ( .A1(G1986), .A2(G290), .ZN(n708) );
  NOR2_X1 U808 ( .A1(G1991), .A2(n867), .ZN(n933) );
  NOR2_X1 U809 ( .A1(n708), .A2(n933), .ZN(n709) );
  NOR2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U811 ( .A1(n927), .A2(n711), .ZN(n712) );
  XNOR2_X1 U812 ( .A(KEYINPUT39), .B(n712), .ZN(n723) );
  XNOR2_X1 U813 ( .A(KEYINPUT37), .B(G2067), .ZN(n724) );
  NAND2_X1 U814 ( .A1(G140), .A2(n890), .ZN(n714) );
  NAND2_X1 U815 ( .A1(G104), .A2(n891), .ZN(n713) );
  NAND2_X1 U816 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U817 ( .A(KEYINPUT34), .B(n715), .ZN(n720) );
  NAND2_X1 U818 ( .A1(G128), .A2(n886), .ZN(n717) );
  NAND2_X1 U819 ( .A1(G116), .A2(n887), .ZN(n716) );
  NAND2_X1 U820 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U821 ( .A(KEYINPUT35), .B(n718), .Z(n719) );
  NOR2_X1 U822 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U823 ( .A(KEYINPUT36), .B(n721), .ZN(n873) );
  NOR2_X1 U824 ( .A1(n724), .A2(n873), .ZN(n938) );
  NAND2_X1 U825 ( .A1(n938), .A2(n819), .ZN(n722) );
  XNOR2_X1 U826 ( .A(n722), .B(KEYINPUT92), .ZN(n822) );
  NAND2_X1 U827 ( .A1(n723), .A2(n822), .ZN(n725) );
  NAND2_X1 U828 ( .A1(n724), .A2(n873), .ZN(n924) );
  NAND2_X1 U829 ( .A1(n725), .A2(n924), .ZN(n726) );
  NAND2_X1 U830 ( .A1(n726), .A2(n819), .ZN(n826) );
  XOR2_X1 U831 ( .A(G1981), .B(G305), .Z(n952) );
  INV_X1 U832 ( .A(n727), .ZN(n729) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n730) );
  XNOR2_X1 U834 ( .A(KEYINPUT101), .B(n730), .ZN(n961) );
  NOR2_X1 U835 ( .A1(n815), .A2(n961), .ZN(n731) );
  NAND2_X1 U836 ( .A1(KEYINPUT33), .A2(n731), .ZN(n732) );
  NAND2_X1 U837 ( .A1(n952), .A2(n732), .ZN(n811) );
  INV_X1 U838 ( .A(n811), .ZN(n733) );
  NAND2_X1 U839 ( .A1(n733), .A2(KEYINPUT33), .ZN(n804) );
  INV_X1 U840 ( .A(n788), .ZN(n760) );
  NAND2_X1 U841 ( .A1(n760), .A2(G2072), .ZN(n735) );
  INV_X1 U842 ( .A(KEYINPUT27), .ZN(n734) );
  NAND2_X1 U843 ( .A1(G1956), .A2(n788), .ZN(n736) );
  NAND2_X1 U844 ( .A1(n737), .A2(n736), .ZN(n739) );
  INV_X1 U845 ( .A(KEYINPUT96), .ZN(n738) );
  XNOR2_X1 U846 ( .A(n739), .B(n738), .ZN(n753) );
  XNOR2_X1 U847 ( .A(n741), .B(n740), .ZN(n757) );
  AND2_X1 U848 ( .A1(n760), .A2(G1996), .ZN(n742) );
  XOR2_X1 U849 ( .A(n742), .B(KEYINPUT26), .Z(n744) );
  NAND2_X1 U850 ( .A1(n788), .A2(G1341), .ZN(n743) );
  NAND2_X1 U851 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U852 ( .A1(n972), .A2(n745), .ZN(n749) );
  NAND2_X1 U853 ( .A1(G1348), .A2(n788), .ZN(n747) );
  NAND2_X1 U854 ( .A1(n760), .A2(G2067), .ZN(n746) );
  NAND2_X1 U855 ( .A1(n747), .A2(n746), .ZN(n750) );
  NOR2_X1 U856 ( .A1(n956), .A2(n750), .ZN(n748) );
  OR2_X1 U857 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U858 ( .A1(n956), .A2(n750), .ZN(n751) );
  NAND2_X1 U859 ( .A1(n752), .A2(n751), .ZN(n755) );
  NAND2_X1 U860 ( .A1(n963), .A2(n753), .ZN(n754) );
  NAND2_X1 U861 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U862 ( .A1(n757), .A2(n756), .ZN(n759) );
  XNOR2_X1 U863 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n758) );
  XNOR2_X1 U864 ( .A(n759), .B(n758), .ZN(n765) );
  XNOR2_X1 U865 ( .A(G2078), .B(KEYINPUT25), .ZN(n1006) );
  NOR2_X1 U866 ( .A1(n788), .A2(n1006), .ZN(n762) );
  INV_X1 U867 ( .A(G1961), .ZN(n979) );
  NOR2_X1 U868 ( .A1(n760), .A2(n979), .ZN(n761) );
  NOR2_X1 U869 ( .A1(n762), .A2(n761), .ZN(n773) );
  NAND2_X1 U870 ( .A1(G171), .A2(n773), .ZN(n763) );
  XOR2_X1 U871 ( .A(KEYINPUT95), .B(n763), .Z(n764) );
  NAND2_X1 U872 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U873 ( .A(n766), .B(KEYINPUT98), .ZN(n779) );
  NOR2_X1 U874 ( .A1(G2084), .A2(n788), .ZN(n781) );
  NOR2_X1 U875 ( .A1(G1966), .A2(n815), .ZN(n767) );
  XNOR2_X1 U876 ( .A(KEYINPUT94), .B(n767), .ZN(n780) );
  NOR2_X1 U877 ( .A1(n781), .A2(n780), .ZN(n769) );
  XNOR2_X1 U878 ( .A(n769), .B(n768), .ZN(n770) );
  NAND2_X1 U879 ( .A1(n770), .A2(G8), .ZN(n771) );
  XNOR2_X1 U880 ( .A(n771), .B(KEYINPUT30), .ZN(n772) );
  NOR2_X1 U881 ( .A1(n772), .A2(G168), .ZN(n775) );
  NOR2_X1 U882 ( .A1(G171), .A2(n773), .ZN(n774) );
  NOR2_X1 U883 ( .A1(n775), .A2(n774), .ZN(n777) );
  XNOR2_X1 U884 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U885 ( .A1(n779), .A2(n778), .ZN(n787) );
  INV_X1 U886 ( .A(n780), .ZN(n783) );
  NAND2_X1 U887 ( .A1(G8), .A2(n781), .ZN(n782) );
  INV_X1 U888 ( .A(KEYINPUT100), .ZN(n784) );
  XNOR2_X1 U889 ( .A(n785), .B(n784), .ZN(n799) );
  AND2_X1 U890 ( .A1(G286), .A2(G8), .ZN(n786) );
  NAND2_X1 U891 ( .A1(n787), .A2(n786), .ZN(n795) );
  INV_X1 U892 ( .A(G8), .ZN(n793) );
  NOR2_X1 U893 ( .A1(G1971), .A2(n815), .ZN(n790) );
  NOR2_X1 U894 ( .A1(G2090), .A2(n788), .ZN(n789) );
  NOR2_X1 U895 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U896 ( .A1(n791), .A2(G303), .ZN(n792) );
  OR2_X1 U897 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U898 ( .A1(n795), .A2(n794), .ZN(n797) );
  INV_X1 U899 ( .A(KEYINPUT32), .ZN(n796) );
  XNOR2_X1 U900 ( .A(n797), .B(n796), .ZN(n798) );
  NOR2_X1 U901 ( .A1(G2090), .A2(G303), .ZN(n800) );
  NAND2_X1 U902 ( .A1(G8), .A2(n800), .ZN(n801) );
  NAND2_X1 U903 ( .A1(n809), .A2(n801), .ZN(n802) );
  NAND2_X1 U904 ( .A1(n802), .A2(n815), .ZN(n803) );
  NAND2_X1 U905 ( .A1(n804), .A2(n803), .ZN(n818) );
  NOR2_X1 U906 ( .A1(G1981), .A2(G305), .ZN(n805) );
  XNOR2_X1 U907 ( .A(KEYINPUT24), .B(n805), .ZN(n814) );
  NOR2_X1 U908 ( .A1(G1971), .A2(G303), .ZN(n806) );
  XOR2_X1 U909 ( .A(n806), .B(KEYINPUT102), .Z(n807) );
  AND2_X1 U910 ( .A1(n807), .A2(n961), .ZN(n808) );
  NAND2_X1 U911 ( .A1(G1976), .A2(G288), .ZN(n962) );
  NAND2_X1 U912 ( .A1(n810), .A2(n962), .ZN(n812) );
  NOR2_X1 U913 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U915 ( .A(G1986), .B(G290), .ZN(n958) );
  NAND2_X1 U916 ( .A1(n819), .A2(n958), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n521), .A2(n823), .ZN(n824) );
  XOR2_X1 U918 ( .A(n824), .B(KEYINPUT103), .Z(n825) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n828) );
  XNOR2_X1 U920 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n828), .B(n827), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G82), .ZN(G220) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n835), .ZN(G319) );
  XNOR2_X1 U934 ( .A(G1996), .B(KEYINPUT41), .ZN(n845) );
  XOR2_X1 U935 ( .A(G1981), .B(G1966), .Z(n837) );
  XNOR2_X1 U936 ( .A(G1991), .B(G1986), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(G1976), .B(G1971), .Z(n839) );
  XNOR2_X1 U939 ( .A(G1956), .B(G1961), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U942 ( .A(KEYINPUT108), .B(G2474), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(G229) );
  XOR2_X1 U945 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2678), .B(KEYINPUT43), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2090), .Z(n849) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2096), .B(G2100), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U954 ( .A(G2078), .B(G2084), .Z(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U956 ( .A1(G112), .A2(n887), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G100), .A2(n891), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U959 ( .A1(n886), .A2(G124), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G136), .A2(n890), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT109), .B(n861), .Z(n862) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(G162) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n865) );
  XNOR2_X1 U966 ( .A(KEYINPUT114), .B(KEYINPUT113), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U968 ( .A(G164), .B(G162), .Z(n866) );
  XNOR2_X1 U969 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n875) );
  XOR2_X1 U971 ( .A(G160), .B(n932), .Z(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n899) );
  NAND2_X1 U975 ( .A1(G139), .A2(n890), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G103), .A2(n891), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n885) );
  NAND2_X1 U978 ( .A1(n887), .A2(G115), .ZN(n878) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(n878), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n886), .A2(G127), .ZN(n879) );
  XOR2_X1 U981 ( .A(n879), .B(KEYINPUT110), .Z(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT112), .B(n883), .Z(n884) );
  NOR2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n942) );
  NAND2_X1 U986 ( .A1(G130), .A2(n886), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G118), .A2(n887), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U989 ( .A1(G142), .A2(n890), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G106), .A2(n891), .ZN(n892) );
  NAND2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n894), .Z(n895) );
  NOR2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n942), .B(n897), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U996 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n902) );
  XNOR2_X1 U998 ( .A(G171), .B(G286), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n956), .B(n903), .Z(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U1003 ( .A(G2454), .B(G2435), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G2438), .B(G2427), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n915) );
  XOR2_X1 U1006 ( .A(KEYINPUT105), .B(G2446), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G2443), .B(G2430), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n911), .B(G2451), .Z(n913) );
  XNOR2_X1 U1010 ( .A(G1341), .B(G1348), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n916), .A2(G14), .ZN(n922) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(n922), .ZN(G401) );
  INV_X1 U1022 ( .A(n923), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n931) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n928), .Z(n929) );
  XNOR2_X1 U1027 ( .A(n929), .B(KEYINPUT119), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n941) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(KEYINPUT117), .B(n934), .Z(n936) );
  XNOR2_X1 U1031 ( .A(G160), .B(G2084), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n939), .B(KEYINPUT118), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n947) );
  XOR2_X1 U1036 ( .A(G2072), .B(n942), .Z(n944) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n945), .Z(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n948), .ZN(n950) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n951), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .ZN(n978) );
  XNOR2_X1 U1046 ( .A(G1966), .B(G168), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(n954), .B(KEYINPUT57), .ZN(n976) );
  XNOR2_X1 U1049 ( .A(G1961), .B(G171), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT122), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(G1348), .B(n956), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n970) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n967) );
  XNOR2_X1 U1055 ( .A(G166), .B(G1971), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(n963), .B(G1956), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(KEYINPUT123), .B(n968), .ZN(n969) );
  NOR2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1061 ( .A(KEYINPUT124), .B(n971), .Z(n974) );
  XNOR2_X1 U1062 ( .A(G1341), .B(n972), .ZN(n973) );
  NOR2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1065 ( .A1(n978), .A2(n977), .ZN(n1004) );
  INV_X1 U1066 ( .A(G16), .ZN(n1002) );
  XNOR2_X1 U1067 ( .A(G5), .B(n979), .ZN(n999) );
  XNOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT59), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n980), .B(G4), .ZN(n984) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(G6), .B(G1981), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G20), .B(G1956), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1076 ( .A(KEYINPUT60), .B(n987), .Z(n989) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G21), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n990), .ZN(n997) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G23), .B(G1976), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n994) );
  XOR2_X1 U1083 ( .A(G1986), .B(G24), .Z(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(KEYINPUT58), .B(n995), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(KEYINPUT61), .B(n1000), .Z(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1028) );
  XOR2_X1 U1091 ( .A(G2067), .B(G26), .Z(n1014) );
  XOR2_X1 U1092 ( .A(G1991), .B(G25), .Z(n1005) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(G28), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(G27), .B(n1006), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G1996), .B(G32), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G33), .B(G2072), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(n1015), .B(KEYINPUT53), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(G2084), .B(KEYINPUT54), .Z(n1016) );
  XNOR2_X1 U1103 ( .A(G34), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(KEYINPUT120), .B(G2090), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(G35), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(KEYINPUT55), .B(n1022), .ZN(n1024) );
  INV_X1 U1109 ( .A(G29), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(G11), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(KEYINPUT121), .B(n1026), .Z(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(n1031), .B(KEYINPUT126), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1117 ( .A(G150), .ZN(G311) );
endmodule

