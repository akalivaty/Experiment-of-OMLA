//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT73), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G237), .ZN(new_n192));
  AOI21_X1  g006(.A(G953), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G210), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n194), .B(G101), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(G134), .B2(G137), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT65), .A2(G134), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT65), .A2(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n202), .B2(new_n203), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n206), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n208), .A2(new_n211), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n205), .B1(new_n215), .B2(G131), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .A4(G128), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT1), .B1(new_n219), .B2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n226), .A3(KEYINPUT1), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT68), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT68), .A2(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT64), .B1(new_n217), .B2(G143), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n219), .A3(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n218), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n223), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n216), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n232), .A2(new_n234), .B1(G143), .B2(new_n217), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n211), .A2(new_n214), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT65), .B(G134), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n212), .B1(new_n248), .B2(new_n207), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n200), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n215), .A2(G131), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n246), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n238), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT2), .ZN(new_n255));
  INV_X1    g069(.A(G113), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT69), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(KEYINPUT2), .B2(G113), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT2), .A2(G113), .ZN(new_n261));
  XNOR2_X1  g075(.A(G116), .B(G119), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n262), .B1(new_n260), .B2(new_n261), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n254), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n261), .ZN(new_n267));
  INV_X1    g081(.A(new_n262), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT70), .A3(new_n263), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT74), .B1(new_n253), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n271), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n273), .B(new_n274), .C1(new_n252), .C2(new_n238), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n264), .A2(new_n265), .A3(new_n254), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT70), .B1(new_n269), .B2(new_n263), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT72), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n266), .A2(new_n270), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT71), .B1(new_n216), .B2(new_n237), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n252), .B1(new_n284), .B2(new_n238), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n199), .B1(new_n276), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n266), .A2(new_n270), .A3(new_n280), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n280), .B1(new_n266), .B2(new_n270), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n253), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n199), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT75), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n293), .A3(new_n199), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n198), .B1(new_n287), .B2(new_n295), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n238), .A2(new_n252), .A3(KEYINPUT30), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n231), .A2(new_n236), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n222), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(new_n284), .A3(new_n250), .A4(new_n205), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n250), .A2(new_n251), .ZN(new_n301));
  INV_X1    g115(.A(new_n246), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n303), .A3(new_n283), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n297), .B1(KEYINPUT30), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n286), .B(new_n197), .C1(new_n305), .C2(new_n271), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT31), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT30), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n285), .B2(new_n283), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n273), .B1(new_n309), .B2(new_n297), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT31), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n286), .A4(new_n197), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n296), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  XOR2_X1   g128(.A(new_n314), .B(KEYINPUT76), .Z(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n188), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n307), .A2(new_n312), .ZN(new_n318));
  AOI211_X1 g132(.A(KEYINPUT75), .B(KEYINPUT28), .C1(new_n282), .C2(new_n253), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n293), .B1(new_n290), .B2(new_n199), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n272), .A2(new_n275), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n288), .A2(new_n289), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(new_n304), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT28), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n197), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n188), .B(new_n316), .C1(new_n318), .C2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n187), .B1(new_n317), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n316), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n287), .A2(new_n295), .A3(new_n198), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n310), .A2(new_n286), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n198), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n331), .A2(new_n334), .A3(KEYINPUT29), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n323), .A2(new_n304), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n199), .B1(new_n336), .B2(new_n286), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n295), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT29), .A3(new_n197), .ZN(new_n339));
  INV_X1    g153(.A(G902), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G472), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n329), .A2(new_n330), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n344));
  INV_X1    g158(.A(G119), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G116), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n344), .B(G113), .C1(KEYINPUT5), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n263), .ZN(new_n348));
  INV_X1    g162(.A(G107), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G104), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(G104), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT82), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G104), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G107), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n352), .A2(KEYINPUT82), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G101), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n354), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G101), .B1(new_n356), .B2(new_n350), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n348), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n361), .A2(KEYINPUT83), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n351), .A2(new_n353), .ZN(new_n367));
  INV_X1    g181(.A(new_n350), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n351), .B1(new_n353), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT4), .B(new_n366), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n369), .A2(new_n371), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(new_n361), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n367), .B(new_n368), .C1(new_n376), .C2(new_n351), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(new_n366), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n372), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n365), .B1(new_n273), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G122), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n348), .A2(new_n364), .A3(KEYINPUT87), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n381), .B(KEYINPUT8), .Z(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n348), .A2(new_n364), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n348), .B2(new_n364), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n380), .A2(new_n381), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G224), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT7), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n395));
  INV_X1    g209(.A(G125), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n237), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n246), .A2(G125), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT86), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n394), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n398), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n394), .ZN(new_n404));
  AOI21_X1  g218(.A(G902), .B1(new_n389), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n362), .A2(KEYINPUT4), .B1(new_n377), .B2(new_n366), .ZN(new_n406));
  INV_X1    g220(.A(new_n372), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n385), .B1(new_n408), .B2(new_n271), .ZN(new_n409));
  INV_X1    g223(.A(new_n381), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n385), .B(new_n381), .C1(new_n408), .C2(new_n271), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n403), .A2(KEYINPUT86), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(new_n392), .C1(KEYINPUT86), .C2(new_n400), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n391), .B1(new_n399), .B2(new_n401), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n409), .A2(new_n418), .A3(new_n410), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n405), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n405), .A2(new_n420), .A3(new_n422), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT88), .A3(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n425), .A2(KEYINPUT88), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT9), .B(G234), .ZN(new_n430));
  OAI21_X1  g244(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n431));
  XNOR2_X1  g245(.A(G110), .B(G140), .ZN(new_n432));
  INV_X1    g246(.A(G227), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G953), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n432), .B(new_n434), .Z(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n301), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n302), .B1(new_n406), .B2(new_n407), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT84), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n440), .B(new_n302), .C1(new_n406), .C2(new_n407), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G128), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n222), .B1(new_n444), .B2(new_n239), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n362), .A2(new_n363), .A3(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT85), .B(KEYINPUT10), .Z(new_n447));
  NAND3_X1  g261(.A1(new_n362), .A2(KEYINPUT10), .A3(new_n363), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n446), .A2(new_n447), .B1(new_n237), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n437), .B1(new_n442), .B2(new_n450), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n301), .B(new_n449), .C1(new_n439), .C2(new_n441), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n436), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n449), .B1(new_n439), .B2(new_n441), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n437), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n364), .A2(new_n237), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n362), .A2(new_n363), .A3(new_n445), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n458), .A2(KEYINPUT12), .A3(new_n301), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT12), .B1(new_n458), .B2(new_n301), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n461), .A3(new_n435), .ZN(new_n462));
  AOI211_X1 g276(.A(G469), .B(G902), .C1(new_n453), .C2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n436), .B1(new_n454), .B2(new_n437), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n440), .B1(new_n379), .B2(new_n302), .ZN(new_n465));
  INV_X1    g279(.A(new_n441), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n450), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n301), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n459), .A2(new_n460), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n436), .B1(new_n452), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n471), .A3(G469), .ZN(new_n472));
  NAND2_X1  g286(.A1(G469), .A2(G902), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n431), .B1(new_n463), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G953), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n191), .A2(G237), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n189), .A2(KEYINPUT73), .ZN(new_n479));
  OAI211_X1 g293(.A(G214), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n219), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n193), .A2(G143), .A3(G214), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT18), .A2(G131), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G140), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G125), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n396), .A2(G140), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G146), .ZN(new_n491));
  XNOR2_X1  g305(.A(G125), .B(G140), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n217), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT89), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n484), .A2(new_n486), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n485), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n487), .A3(G125), .ZN(new_n502));
  OAI211_X1 g316(.A(G146), .B(new_n502), .C1(new_n490), .C2(new_n501), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n492), .B(KEYINPUT19), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n505), .B2(new_n217), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n481), .A2(new_n200), .A3(new_n483), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n200), .B1(new_n481), .B2(new_n483), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G113), .B(G122), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n355), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n500), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  INV_X1    g329(.A(new_n509), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n507), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n502), .B1(new_n490), .B2(new_n501), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n217), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n503), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n509), .B2(KEYINPUT17), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n518), .A2(new_n522), .B1(new_n498), .B2(new_n499), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n514), .B(new_n515), .C1(new_n523), .C2(new_n513), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT20), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n522), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n500), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n510), .A2(new_n513), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n530), .A2(new_n512), .B1(new_n531), .B2(new_n500), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n515), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G475), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n513), .A2(KEYINPUT92), .ZN(new_n537));
  AOI21_X1  g351(.A(G902), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n523), .A2(KEYINPUT92), .A3(new_n513), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n543));
  INV_X1    g357(.A(G217), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n430), .A2(new_n544), .A3(G953), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G134), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n219), .A2(G128), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT13), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI211_X1 g365(.A(KEYINPUT93), .B(KEYINPUT13), .C1(new_n219), .C2(G128), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT68), .B(G128), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n443), .A2(G143), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n554), .A2(G143), .B1(KEYINPUT13), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n547), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G122), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G116), .ZN(new_n559));
  INV_X1    g373(.A(G116), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G122), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G107), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n561), .A3(new_n349), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G143), .B1(new_n228), .B2(new_n229), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n248), .A3(new_n549), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n557), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n559), .A2(KEYINPUT14), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n562), .A2(new_n570), .A3(G107), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n559), .B(new_n561), .C1(KEYINPUT14), .C2(new_n349), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n248), .B1(new_n566), .B2(new_n549), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n575), .B2(new_n567), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n546), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT93), .B1(new_n555), .B2(KEYINPUT13), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n549), .A2(new_n548), .A3(new_n550), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n555), .A2(KEYINPUT13), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n578), .A2(new_n566), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G134), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n567), .A3(new_n565), .ZN(new_n583));
  INV_X1    g397(.A(new_n567), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n572), .B(new_n571), .C1(new_n584), .C2(new_n574), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n585), .A3(new_n545), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n577), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G478), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT15), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n543), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n569), .A2(new_n576), .A3(new_n546), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n545), .B1(new_n583), .B2(new_n585), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n340), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT94), .A3(new_n589), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n340), .B(new_n590), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n587), .A2(KEYINPUT95), .A3(new_n590), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT96), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n596), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(G234), .A2(G237), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(G952), .A3(new_n477), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT21), .B(G898), .Z(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(G902), .A3(G953), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n611), .B(KEYINPUT97), .Z(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n542), .A2(new_n606), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n429), .A2(new_n476), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n554), .A2(G119), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n345), .A2(G128), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT24), .B(G110), .Z(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT78), .B(G110), .Z(new_n621));
  NAND3_X1  g435(.A1(new_n616), .A2(KEYINPUT23), .A3(new_n617), .ZN(new_n622));
  OR3_X1    g436(.A1(new_n345), .A2(KEYINPUT23), .A3(G128), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n503), .B(new_n493), .C1(new_n620), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n618), .A2(new_n619), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(G110), .A3(new_n623), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n521), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT80), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT80), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n625), .A2(new_n631), .A3(new_n628), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n477), .A2(G221), .A3(G234), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT79), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT22), .B(G137), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n630), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n629), .A2(KEYINPUT80), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n544), .B1(G234), .B2(new_n340), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT81), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT81), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n640), .A2(new_n645), .A3(new_n642), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n638), .B2(new_n639), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT25), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI211_X1 g463(.A(KEYINPUT25), .B(G902), .C1(new_n638), .C2(new_n639), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n644), .B(new_n646), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n343), .A2(new_n615), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G101), .ZN(G3));
  OAI21_X1  g468(.A(new_n316), .B1(new_n318), .B2(new_n326), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT77), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n327), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n340), .B1(new_n318), .B2(new_n326), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(G472), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n428), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n424), .B2(new_n425), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n475), .A2(new_n651), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n592), .A2(new_n593), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT33), .Z(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(G478), .A3(new_n340), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(G478), .B2(new_n587), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n542), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n665), .A2(new_n613), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G104), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n534), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n532), .A2(KEYINPUT99), .A3(new_n533), .A4(new_n515), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n527), .A3(new_n528), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n540), .A2(KEYINPUT100), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n540), .A2(KEYINPUT100), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n679), .A2(new_n682), .A3(new_n612), .A4(new_n606), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT101), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n680), .A2(new_n681), .B1(new_n603), .B2(new_n605), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n685), .A2(new_n679), .A3(new_n686), .A4(new_n612), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n665), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT102), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT35), .B(G107), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G9));
  NOR2_X1   g505(.A1(new_n637), .A2(KEYINPUT36), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n629), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n642), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n649), .B2(new_n650), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n661), .A2(new_n615), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT37), .B(G110), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  OR2_X1    g512(.A1(new_n610), .A2(G900), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n608), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n685), .A2(new_n679), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n424), .A2(new_n425), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n428), .ZN(new_n703));
  INV_X1    g517(.A(new_n695), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n343), .A2(new_n476), .A3(new_n701), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  AND2_X1   g521(.A1(new_n336), .A2(new_n286), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n306), .B1(new_n197), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n709), .A2(KEYINPUT103), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n340), .B1(new_n709), .B2(KEYINPUT103), .ZN(new_n711));
  OAI21_X1  g525(.A(G472), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n329), .A2(new_n330), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n542), .A2(new_n606), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n426), .A2(new_n427), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT38), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n704), .A2(new_n428), .ZN(new_n718));
  OR4_X1    g532(.A1(new_n714), .A2(new_n715), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n700), .B(KEYINPUT39), .Z(new_n723));
  NOR2_X1   g537(.A1(new_n475), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT40), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  INV_X1    g541(.A(new_n700), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n670), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n343), .A2(new_n476), .A3(new_n705), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT105), .B(G146), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G48));
  NOR2_X1   g546(.A1(new_n670), .A2(new_n613), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n453), .A2(new_n462), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n340), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  INV_X1    g550(.A(G469), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n737), .A3(new_n340), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n431), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n703), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n343), .A2(new_n652), .A3(new_n733), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND2_X1  g557(.A1(new_n684), .A2(new_n687), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n343), .A2(new_n744), .A3(new_n652), .A4(new_n740), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G116), .ZN(G18));
  AND2_X1   g560(.A1(new_n614), .A2(new_n695), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n343), .A2(new_n740), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  AND3_X1   g563(.A1(new_n542), .A2(new_n606), .A3(new_n612), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n737), .B1(new_n734), .B2(new_n340), .ZN(new_n751));
  INV_X1    g565(.A(new_n431), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n751), .A2(new_n463), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n753), .A3(new_n663), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n338), .A2(new_n197), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n316), .B1(new_n755), .B2(new_n318), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n659), .A2(new_n652), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT106), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n542), .A2(new_n606), .A3(new_n612), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n739), .A2(new_n759), .A3(new_n703), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n659), .A2(new_n652), .A3(new_n756), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  AND2_X1   g579(.A1(new_n659), .A2(new_n756), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n740), .A3(new_n695), .A4(new_n729), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  NAND2_X1  g582(.A1(new_n655), .A2(new_n187), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n342), .A2(new_n330), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n652), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n475), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT107), .B(new_n431), .C1(new_n463), .C2(new_n474), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n662), .B1(new_n426), .B2(new_n427), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n771), .A2(KEYINPUT42), .A3(new_n729), .A4(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n343), .A2(new_n652), .A3(new_n776), .A4(new_n729), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT109), .B(G131), .Z(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G33));
  AND2_X1   g599(.A1(new_n343), .A2(new_n652), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n701), .A3(new_n776), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  NAND3_X1  g602(.A1(new_n669), .A2(new_n535), .A3(new_n541), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT43), .Z(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n660), .A3(new_n695), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT44), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(KEYINPUT44), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n775), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n792), .B1(new_n794), .B2(KEYINPUT113), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n469), .B2(new_n471), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n737), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT45), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT46), .B1(new_n799), .B2(new_n473), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT111), .Z(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n473), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT110), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(KEYINPUT110), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n801), .A2(new_n738), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n723), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n431), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT112), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n795), .B(new_n808), .C1(KEYINPUT113), .C2(new_n794), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT114), .B(G137), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n809), .B(new_n810), .ZN(G39));
  NAND2_X1  g625(.A1(new_n805), .A2(new_n431), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n729), .A2(new_n651), .A3(new_n775), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n343), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NOR2_X1   g632(.A1(new_n751), .A2(new_n463), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT49), .Z(new_n820));
  NAND3_X1  g634(.A1(new_n652), .A2(new_n428), .A3(new_n431), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n820), .A2(new_n789), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n714), .A3(new_n717), .ZN(new_n823));
  INV_X1    g637(.A(new_n608), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n790), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n775), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n739), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n771), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT48), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n740), .A3(new_n761), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n830), .A2(G952), .A3(new_n477), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n714), .A2(new_n652), .A3(new_n824), .A4(new_n827), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT123), .Z(new_n833));
  OAI211_X1 g647(.A(new_n829), .B(new_n831), .C1(new_n833), .C2(new_n670), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n825), .A2(new_n761), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n717), .A2(new_n662), .A3(new_n753), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT50), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n825), .A2(new_n695), .A3(new_n766), .A4(new_n827), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n833), .A2(new_n542), .A3(new_n669), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n840), .A2(KEYINPUT51), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n835), .A2(new_n826), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n751), .A2(new_n463), .A3(new_n431), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n814), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n834), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n845), .A2(KEYINPUT122), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(KEYINPUT122), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n847), .A2(new_n841), .A3(new_n840), .A4(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n663), .A2(new_n542), .A3(new_n606), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n475), .A2(new_n695), .A3(new_n728), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n713), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n706), .A2(new_n730), .A3(new_n767), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT117), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n741), .A2(new_n745), .A3(new_n764), .A4(new_n748), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n343), .A2(new_n652), .A3(new_n615), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n664), .A2(new_n657), .A3(new_n659), .ZN(new_n867));
  INV_X1    g681(.A(new_n602), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n670), .B1(new_n542), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n429), .A3(new_n612), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n429), .A2(new_n476), .A3(new_n614), .A4(new_n695), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n867), .A2(new_n870), .B1(new_n871), .B2(new_n660), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT115), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n867), .A2(new_n870), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n653), .A3(new_n696), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n865), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n695), .A2(new_n776), .A3(new_n729), .A4(new_n766), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n679), .A2(new_n868), .A3(new_n682), .A4(new_n700), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n826), .A2(new_n704), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n343), .A3(new_n476), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT116), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n880), .A2(new_n343), .A3(new_n883), .A4(new_n476), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n878), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n877), .A2(new_n783), .A3(new_n787), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n853), .B1(new_n864), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n858), .B(KEYINPUT52), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n886), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n888), .B2(new_n887), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n852), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n891), .B1(new_n886), .B2(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n873), .A2(new_n876), .ZN(new_n897));
  INV_X1    g711(.A(new_n865), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n885), .ZN(new_n899));
  INV_X1    g713(.A(new_n787), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n778), .A2(new_n780), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT108), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n900), .B1(new_n904), .B2(new_n777), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n863), .A2(new_n899), .A3(new_n905), .A4(KEYINPUT53), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n896), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n895), .A2(KEYINPUT120), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT120), .B1(new_n895), .B2(new_n908), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n851), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(G952), .A2(G953), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n823), .B1(new_n911), .B2(new_n912), .ZN(G75));
  INV_X1    g727(.A(new_n417), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n340), .B1(new_n896), .B2(new_n906), .ZN(new_n915));
  AOI211_X1 g729(.A(KEYINPUT55), .B(KEYINPUT56), .C1(new_n915), .C2(G210), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT55), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n907), .A2(G210), .A3(G902), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n413), .A2(new_n419), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  INV_X1    g737(.A(G210), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n924), .B(new_n340), .C1(new_n896), .C2(new_n906), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT55), .B1(new_n925), .B2(KEYINPUT56), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n918), .A2(new_n917), .A3(new_n919), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n927), .A3(new_n417), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n921), .A2(new_n923), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n477), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n923), .B1(new_n921), .B2(new_n928), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G51));
  XNOR2_X1  g748(.A(new_n907), .B(KEYINPUT54), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n473), .B(KEYINPUT57), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n734), .B(KEYINPUT125), .Z(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n915), .A2(new_n798), .A3(new_n797), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n930), .B1(new_n939), .B2(new_n940), .ZN(G54));
  AND3_X1   g755(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n931), .B1(new_n942), .B2(new_n532), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n532), .B2(new_n942), .ZN(G60));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT59), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n935), .A2(new_n667), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n931), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n909), .A2(new_n910), .A3(new_n946), .ZN(new_n949));
  INV_X1    g763(.A(new_n667), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT60), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n896), .B2(new_n906), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n930), .B1(new_n954), .B2(new_n693), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n640), .B2(new_n954), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g771(.A(new_n477), .B1(new_n609), .B2(G224), .ZN(new_n958));
  INV_X1    g772(.A(new_n877), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n477), .ZN(new_n960));
  INV_X1    g774(.A(G898), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n923), .B1(new_n961), .B2(G953), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT126), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n960), .B(new_n963), .ZN(G69));
  AND2_X1   g778(.A1(new_n809), .A2(new_n817), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n706), .A2(new_n730), .A3(new_n767), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n808), .A2(new_n771), .A3(new_n855), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n965), .A2(new_n905), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n477), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n305), .B(new_n505), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(G900), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n726), .A2(new_n966), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT62), .Z(new_n976));
  NAND4_X1  g790(.A1(new_n786), .A2(new_n724), .A3(new_n775), .A4(new_n869), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n965), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n477), .A3(new_n971), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n433), .B2(new_n972), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n978), .B2(new_n959), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n197), .A3(new_n332), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n889), .A2(new_n894), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n333), .B(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n306), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n984), .B1(new_n968), .B2(new_n959), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n991), .A2(new_n286), .A3(new_n198), .A4(new_n310), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n931), .A2(new_n986), .A3(new_n990), .A4(new_n992), .ZN(G57));
endmodule


