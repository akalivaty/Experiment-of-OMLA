//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G134), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT65), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G134), .ZN(new_n194));
  AOI21_X1  g008(.A(G137), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(new_n188), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(new_n194), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(new_n189), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n197), .B2(new_n189), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n196), .A2(KEYINPUT66), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n193), .A2(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n191), .A2(KEYINPUT65), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n188), .B(new_n189), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n190), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(G134), .ZN(new_n209));
  AOI21_X1  g023(.A(G131), .B1(new_n209), .B2(G137), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n203), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n199), .B1(new_n202), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n218), .B2(new_n219), .ZN(new_n223));
  OAI22_X1  g037(.A1(new_n221), .A2(new_n223), .B1(new_n217), .B2(new_n222), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n212), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G116), .B(G119), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(new_n196), .B2(new_n201), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n208), .A2(new_n203), .A3(new_n210), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n233), .A3(G128), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n214), .B(new_n216), .C1(KEYINPUT1), .C2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n189), .A2(G134), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n195), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n232), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n226), .A2(new_n229), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n229), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n224), .B1(new_n232), .B2(new_n199), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n237), .A2(new_n239), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n231), .B2(new_n230), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n242), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT28), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n251), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n248), .A2(new_n250), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n187), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT71), .ZN(new_n261));
  INV_X1    g075(.A(new_n257), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT30), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n226), .A2(KEYINPUT67), .A3(new_n263), .A4(new_n240), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n265), .B(new_n266), .C1(new_n243), .C2(new_n245), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n229), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n241), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n262), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n258), .A3(new_n259), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(new_n187), .C1(new_n258), .C2(new_n259), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n270), .A2(new_n258), .A3(new_n275), .A4(new_n259), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n261), .A2(new_n272), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G472), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n264), .A2(new_n267), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n242), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n241), .A3(new_n257), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT69), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n268), .A2(new_n269), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n257), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(KEYINPUT31), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n257), .B1(new_n248), .B2(new_n250), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n268), .A2(new_n269), .A3(new_n262), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n279), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n293), .ZN(new_n295));
  AOI211_X1 g109(.A(KEYINPUT32), .B(new_n295), .C1(new_n287), .C2(new_n291), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n278), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT20), .ZN(new_n298));
  NOR2_X1   g112(.A1(G475), .A2(G902), .ZN(new_n299));
  XOR2_X1   g113(.A(G113), .B(G122), .Z(new_n300));
  XOR2_X1   g114(.A(KEYINPUT86), .B(G104), .Z(new_n301));
  XOR2_X1   g115(.A(new_n300), .B(new_n301), .Z(new_n302));
  NAND3_X1  g116(.A1(new_n252), .A2(new_n253), .A3(G214), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n215), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n252), .A2(new_n253), .A3(G143), .A4(G214), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT18), .A2(G131), .ZN(new_n308));
  OR3_X1    g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n306), .B2(new_n307), .ZN(new_n310));
  XOR2_X1   g124(.A(G125), .B(G140), .Z(new_n311));
  OR2_X1    g125(.A1(new_n311), .A2(G146), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT74), .A2(G125), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(KEYINPUT74), .A2(G125), .A3(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G146), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n309), .A2(new_n310), .B1(new_n312), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n306), .A2(G131), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n304), .A2(new_n200), .A3(new_n305), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  MUX2_X1   g137(.A(new_n323), .B(new_n321), .S(KEYINPUT17), .Z(new_n324));
  AND3_X1   g138(.A1(new_n315), .A2(KEYINPUT16), .A3(new_n316), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT16), .B1(new_n314), .B2(G125), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n213), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n329));
  OAI21_X1  g143(.A(G146), .B1(new_n325), .B2(new_n326), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(KEYINPUT75), .A3(new_n213), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI211_X1 g147(.A(new_n302), .B(new_n320), .C1(new_n324), .C2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n302), .ZN(new_n335));
  INV_X1    g149(.A(new_n320), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n315), .A2(KEYINPUT19), .A3(new_n316), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n337), .B(new_n338), .C1(new_n311), .C2(KEYINPUT19), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n338), .B2(new_n337), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n213), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n330), .A3(new_n323), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n335), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n298), .B(new_n299), .C1(new_n334), .C2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n334), .A2(new_n343), .ZN(new_n347));
  INV_X1    g161(.A(new_n299), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT20), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n320), .B1(new_n324), .B2(new_n333), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n335), .ZN(new_n351));
  INV_X1    g165(.A(new_n343), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT87), .A3(new_n298), .A4(new_n299), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n346), .A2(new_n349), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n350), .A2(new_n335), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n187), .B1(new_n356), .B2(new_n334), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G475), .ZN(new_n358));
  INV_X1    g172(.A(G952), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G953), .ZN(new_n360));
  NAND2_X1  g174(.A1(G234), .A2(G237), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(G902), .A3(G953), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT21), .B(G898), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G478), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT15), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT88), .B(G122), .ZN(new_n372));
  INV_X1    g186(.A(G116), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n373), .A2(G122), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G107), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n376), .B1(KEYINPUT14), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n215), .A2(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n235), .A2(G143), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT89), .B1(new_n235), .B2(G143), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n197), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n209), .B(new_n379), .C1(new_n382), .C2(new_n383), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT14), .B1(new_n372), .B2(new_n373), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(G107), .C1(new_n374), .C2(new_n375), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n378), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT13), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n379), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n215), .A2(KEYINPUT13), .A3(G128), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n392), .B(new_n393), .C1(new_n382), .C2(new_n383), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G134), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT90), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n386), .A2(KEYINPUT91), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n386), .A2(KEYINPUT91), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n376), .A2(new_n377), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n374), .A2(G107), .A3(new_n375), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n390), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  XOR2_X1   g216(.A(KEYINPUT9), .B(G234), .Z(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT77), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n404), .A2(new_n405), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n390), .B(new_n406), .C1(new_n396), .C2(new_n401), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n371), .B1(new_n410), .B2(new_n187), .ZN(new_n411));
  AOI211_X1 g225(.A(G902), .B(new_n370), .C1(new_n408), .C2(new_n409), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n355), .A2(new_n358), .A3(new_n368), .A4(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G140), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n253), .A2(G227), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT78), .ZN(new_n418));
  INV_X1    g232(.A(G104), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT3), .B1(new_n419), .B2(G107), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n377), .A3(G104), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(G107), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n424), .A2(G101), .ZN(new_n425));
  INV_X1    g239(.A(G101), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n420), .A2(new_n422), .A3(new_n426), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n418), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(G101), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(KEYINPUT78), .A3(KEYINPUT4), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n424), .A2(new_n433), .A3(G101), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT79), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT79), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n424), .A2(new_n436), .A3(new_n433), .A4(G101), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n224), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n198), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n208), .A2(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n230), .A2(new_n231), .B1(new_n441), .B2(G131), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n377), .A3(G104), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT80), .B1(new_n419), .B2(G107), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n377), .A2(G104), .ZN(new_n446));
  OAI211_X1 g260(.A(G101), .B(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n234), .A2(new_n447), .A3(new_n427), .A4(new_n236), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n448), .A2(KEYINPUT10), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(KEYINPUT10), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n439), .A2(new_n442), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n442), .B1(new_n439), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n417), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n432), .A2(new_n438), .B1(new_n449), .B2(new_n450), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n417), .B1(new_n455), .B2(new_n442), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n234), .A2(new_n236), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n447), .A2(new_n427), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n448), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n457), .B1(new_n442), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n212), .A2(KEYINPUT12), .A3(new_n461), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n454), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G469), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n187), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n187), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n439), .A2(new_n451), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n212), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n456), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n417), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n463), .A2(new_n464), .B1(new_n455), .B2(new_n442), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n474), .B(G469), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G221), .B1(new_n404), .B2(G902), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n414), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G210), .B1(G237), .B2(G902), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT83), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT5), .ZN(new_n487));
  INV_X1    g301(.A(G119), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(G116), .ZN(new_n489));
  XOR2_X1   g303(.A(G116), .B(G119), .Z(new_n490));
  OAI211_X1 g304(.A(G113), .B(new_n489), .C1(new_n490), .C2(new_n487), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n490), .A2(new_n228), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n427), .A4(new_n447), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n229), .B1(new_n435), .B2(new_n437), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n432), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G110), .B(G122), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n486), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n432), .A2(new_n495), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n493), .ZN(new_n500));
  INV_X1    g314(.A(new_n497), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n486), .A3(new_n501), .ZN(new_n504));
  INV_X1    g318(.A(G125), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n237), .A2(new_n505), .ZN(new_n506));
  OAI221_X1 g320(.A(G125), .B1(new_n217), .B2(new_n222), .C1(new_n221), .C2(new_n223), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n253), .A2(G224), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n503), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT81), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT82), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n509), .A2(KEYINPUT7), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n506), .A2(KEYINPUT82), .A3(new_n507), .A4(new_n515), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n491), .A2(new_n492), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n459), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n493), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n497), .B(KEYINPUT8), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n522), .A2(new_n523), .B1(new_n508), .B2(new_n516), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n496), .A2(new_n497), .ZN(new_n526));
  AOI21_X1  g340(.A(G902), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n504), .A4(new_n510), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n485), .B1(new_n513), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n511), .A2(new_n512), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n531), .A2(new_n484), .A3(new_n528), .A4(new_n527), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n483), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n481), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n405), .B1(G234), .B2(new_n187), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G110), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n488), .B2(G128), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n539), .A2(KEYINPUT23), .B1(new_n488), .B2(G128), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT23), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n538), .B(new_n541), .C1(new_n488), .C2(G128), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n537), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n544), .B2(new_n543), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT24), .B(G110), .Z(new_n547));
  XNOR2_X1  g361(.A(G119), .B(G128), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n546), .A2(new_n331), .A3(new_n332), .A4(new_n549), .ZN(new_n550));
  OAI22_X1  g364(.A1(new_n543), .A2(G110), .B1(new_n548), .B2(new_n547), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n330), .A3(new_n312), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G137), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n550), .A2(new_n552), .A3(new_n556), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n187), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT25), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n558), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n559), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n536), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n558), .A2(new_n559), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n536), .A2(new_n187), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT76), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n297), .A2(new_n534), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G101), .ZN(G3));
  NAND2_X1  g386(.A1(new_n292), .A2(new_n293), .ZN(new_n573));
  INV_X1    g387(.A(new_n570), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n480), .ZN(new_n575));
  INV_X1    g389(.A(G472), .ZN(new_n576));
  AOI21_X1  g390(.A(G902), .B1(new_n287), .B2(new_n291), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n573), .B(new_n575), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n410), .A2(KEYINPUT92), .A3(KEYINPUT33), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT33), .B1(new_n410), .B2(KEYINPUT92), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n187), .A2(G478), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n408), .B2(new_n409), .ZN(new_n583));
  OAI22_X1  g397(.A1(new_n581), .A2(new_n582), .B1(G478), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n355), .A2(new_n358), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n484), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n513), .B2(new_n529), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n483), .B1(new_n588), .B2(new_n532), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR4_X1   g404(.A1(new_n578), .A2(new_n367), .A3(new_n586), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT93), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT34), .B(G104), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  AOI21_X1  g408(.A(new_n295), .B1(new_n287), .B2(new_n291), .ZN(new_n595));
  INV_X1    g409(.A(new_n577), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(G472), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n367), .B(KEYINPUT94), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n413), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n349), .A2(new_n344), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n358), .A3(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n590), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n597), .A2(new_n575), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  NOR2_X1   g420(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n553), .B(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n608), .A2(new_n568), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n564), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n597), .A2(new_n534), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT37), .B(G110), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G12));
  NOR3_X1   g428(.A1(new_n590), .A2(new_n480), .A3(new_n610), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n297), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G900), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n363), .B1(new_n365), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n602), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G128), .ZN(G30));
  XNOR2_X1  g435(.A(new_n595), .B(new_n279), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n283), .A2(new_n286), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n247), .B2(new_n262), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n624), .B2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n530), .A2(new_n532), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n480), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n618), .B(KEYINPUT39), .Z(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n632), .A2(KEYINPUT40), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n585), .A2(new_n600), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n610), .A2(new_n482), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n634), .B(new_n635), .C1(new_n632), .C2(KEYINPUT40), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n626), .A2(new_n629), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G143), .ZN(G45));
  NOR2_X1   g452(.A1(new_n586), .A2(new_n618), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n616), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT96), .B(G146), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G48));
  NOR2_X1   g456(.A1(new_n468), .A2(KEYINPUT97), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n455), .A2(new_n442), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n473), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n645), .A2(new_n417), .B1(new_n465), .B2(new_n456), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n643), .B1(new_n646), .B2(G902), .ZN(new_n647));
  INV_X1    g461(.A(new_n643), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n467), .A2(new_n187), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n649), .A3(new_n479), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT98), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n647), .A2(new_n649), .A3(new_n652), .A4(new_n479), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n574), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n590), .A2(new_n586), .A3(new_n367), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n297), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT41), .B(G113), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(G15));
  NAND3_X1  g474(.A1(new_n297), .A2(new_n603), .A3(new_n655), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT100), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n297), .A2(new_n603), .A3(new_n663), .A4(new_n655), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G116), .ZN(G18));
  NAND2_X1  g480(.A1(new_n588), .A2(new_n532), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(new_n651), .A3(new_n482), .A4(new_n653), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n589), .A2(new_n670), .A3(new_n653), .A4(new_n651), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n414), .A2(new_n610), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n297), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G119), .ZN(G21));
  NAND3_X1  g489(.A1(new_n589), .A2(new_n585), .A3(new_n600), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n676), .A2(new_n599), .A3(new_n654), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(G472), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n595), .B1(new_n596), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n570), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G122), .ZN(G24));
  INV_X1    g495(.A(new_n678), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n573), .B(new_n611), .C1(new_n577), .C2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n639), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n672), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G125), .ZN(G27));
  AOI21_X1  g501(.A(new_n574), .B1(new_n622), .B2(new_n278), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n477), .A2(new_n471), .ZN(new_n690));
  AOI211_X1 g504(.A(G469), .B(G902), .C1(new_n454), .C2(new_n466), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n469), .A2(KEYINPUT103), .A3(new_n471), .A4(new_n477), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n479), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n627), .A2(new_n483), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n692), .A2(new_n693), .A3(new_n697), .A4(new_n479), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT105), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n688), .A2(new_n703), .A3(new_n639), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n688), .A2(new_n703), .A3(KEYINPUT42), .A4(new_n639), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n706), .A2(KEYINPUT106), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n200), .ZN(G33));
  XNOR2_X1  g527(.A(new_n619), .B(KEYINPUT107), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n688), .A2(new_n703), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G134), .ZN(G36));
  OAI21_X1  g530(.A(new_n474), .B1(new_n476), .B2(new_n475), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT108), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n468), .B1(new_n717), .B2(new_n718), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n722), .A2(new_n723), .A3(new_n470), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n723), .B1(new_n722), .B2(new_n470), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n469), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n726), .A2(new_n479), .A3(new_n631), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n696), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n584), .A2(new_n358), .A3(new_n355), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n585), .B2(KEYINPUT109), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n729), .B(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n732), .A2(new_n611), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n733), .A2(KEYINPUT44), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT44), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n728), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n189), .ZN(G39));
  NAND3_X1  g552(.A1(new_n639), .A2(new_n574), .A3(new_n696), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n726), .A2(new_n479), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n479), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n297), .B(new_n739), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n314), .ZN(G42));
  INV_X1    g559(.A(new_n479), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n574), .A2(new_n483), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n647), .A2(new_n649), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n747), .B(new_n729), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT110), .Z(new_n751));
  INV_X1    g565(.A(new_n626), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n629), .B1(new_n748), .B2(new_n749), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT111), .Z(new_n755));
  INV_X1    g569(.A(new_n696), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n654), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n752), .A2(new_n570), .A3(new_n363), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n360), .B1(new_n758), .B2(new_n586), .ZN(new_n759));
  INV_X1    g573(.A(new_n688), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n732), .A2(new_n363), .A3(new_n757), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT48), .ZN(new_n763));
  AND4_X1   g577(.A1(new_n570), .A2(new_n732), .A3(new_n363), .A4(new_n679), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n759), .B(new_n763), .C1(new_n672), .C2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n629), .A2(new_n482), .A3(new_n654), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT50), .Z(new_n768));
  OR3_X1    g582(.A1(new_n758), .A2(new_n585), .A3(new_n584), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n768), .B(new_n769), .C1(new_n683), .C2(new_n761), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n742), .A2(new_n743), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n746), .B2(new_n749), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n764), .A2(new_n696), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT51), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n771), .A2(KEYINPUT118), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n749), .A2(new_n746), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT119), .Z(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n771), .B2(KEYINPUT118), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n773), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n770), .A2(new_n779), .ZN(new_n780));
  OAI221_X1 g594(.A(new_n765), .B1(new_n770), .B2(new_n774), .C1(new_n780), .C2(KEYINPUT51), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n674), .A2(new_n680), .A3(new_n657), .ZN(new_n784));
  INV_X1    g598(.A(new_n618), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n413), .A2(new_n601), .A3(new_n358), .A4(new_n785), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n756), .A2(new_n480), .A3(new_n610), .A4(new_n786), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n703), .A2(new_n685), .B1(new_n787), .B2(new_n297), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n784), .A2(new_n665), .A3(new_n715), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n586), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n533), .A2(new_n598), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n597), .A2(new_n575), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n571), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT112), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n585), .A2(new_n413), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n533), .A2(new_n598), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n481), .A2(new_n533), .A3(new_n611), .ZN(new_n797));
  OAI22_X1  g611(.A1(new_n578), .A2(new_n796), .B1(new_n734), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT113), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n800));
  OAI221_X1 g614(.A(new_n800), .B1(new_n734), .B2(new_n797), .C1(new_n578), .C2(new_n796), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n571), .A2(new_n792), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n794), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n789), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n807), .A3(new_n710), .A4(new_n711), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n297), .B(new_n615), .C1(new_n619), .C2(new_n639), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n610), .A2(new_n785), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT115), .Z(new_n811));
  INV_X1    g625(.A(new_n676), .ZN(new_n812));
  INV_X1    g626(.A(new_n694), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n686), .B(new_n809), .C1(new_n752), .C2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n626), .A2(new_n812), .A3(new_n813), .A4(new_n811), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(new_n686), .A3(KEYINPUT52), .A4(new_n809), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT116), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n808), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n706), .A2(KEYINPUT106), .A3(new_n707), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT106), .B1(new_n706), .B2(new_n707), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n807), .B1(new_n828), .B2(new_n806), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n783), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n806), .A2(new_n710), .A3(new_n711), .A4(new_n820), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n783), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n782), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n783), .B1(new_n706), .B2(new_n707), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n806), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n836), .A2(new_n824), .B1(new_n831), .B2(new_n783), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n782), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT117), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n782), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n789), .A2(new_n805), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT114), .B1(new_n712), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n808), .A3(new_n824), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n832), .B1(new_n844), .B2(new_n783), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n840), .B(new_n841), .C1(new_n845), .C2(new_n782), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n781), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(G952), .A2(G953), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n755), .B1(new_n847), .B2(new_n848), .ZN(G75));
  NAND2_X1  g663(.A1(new_n503), .A2(new_n504), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(new_n510), .Z(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT55), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(KEYINPUT122), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(KEYINPUT122), .ZN(new_n855));
  XOR2_X1   g669(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n837), .A2(new_n187), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n485), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(KEYINPUT120), .A3(new_n485), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n857), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n359), .A2(G953), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT123), .Z(new_n865));
  AOI21_X1  g679(.A(KEYINPUT56), .B1(new_n858), .B2(G210), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n853), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n863), .A2(new_n867), .ZN(G51));
  INV_X1    g682(.A(new_n865), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n470), .B(KEYINPUT57), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n836), .A2(new_n824), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n831), .A2(new_n783), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n782), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(new_n782), .B2(new_n837), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n837), .B2(new_n782), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n870), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n467), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n858), .A2(new_n722), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n869), .B1(new_n878), .B2(new_n879), .ZN(G54));
  NAND3_X1  g694(.A1(new_n858), .A2(KEYINPUT58), .A3(G475), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n881), .A2(new_n353), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n353), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n869), .B1(new_n882), .B2(new_n883), .ZN(G60));
  NAND2_X1  g698(.A1(G478), .A2(G902), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT59), .Z(new_n886));
  NOR2_X1   g700(.A1(new_n581), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n875), .B2(new_n876), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n865), .ZN(new_n889));
  INV_X1    g703(.A(new_n886), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n839), .A2(new_n846), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n889), .B1(new_n891), .B2(new_n581), .ZN(G63));
  XNOR2_X1  g706(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n893));
  NAND2_X1  g707(.A1(G217), .A2(G902), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n837), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(new_n565), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n608), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n865), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n897), .A2(KEYINPUT61), .A3(new_n865), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G66));
  INV_X1    g717(.A(G224), .ZN(new_n904));
  OAI21_X1  g718(.A(G953), .B1(new_n366), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n784), .A2(new_n665), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n805), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n907), .B2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n850), .B1(G898), .B2(new_n253), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(G69));
  NAND3_X1  g724(.A1(new_n727), .A2(new_n688), .A3(new_n812), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n686), .A2(new_n809), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n715), .A3(new_n912), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n712), .A2(new_n737), .A3(new_n744), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n253), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n280), .B(new_n340), .Z(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(G900), .B2(G953), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n737), .A2(new_n744), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n912), .A2(new_n637), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n920), .A2(KEYINPUT62), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(KEYINPUT62), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n790), .A2(new_n795), .ZN(new_n923));
  OR4_X1    g737(.A1(new_n760), .A2(new_n632), .A3(new_n756), .A4(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n919), .A2(new_n921), .A3(new_n922), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n253), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n916), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT126), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n918), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n918), .A2(KEYINPUT127), .A3(new_n927), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n928), .B1(new_n918), .B2(KEYINPUT127), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G72));
  NAND2_X1  g747(.A1(G472), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT63), .Z(new_n935));
  INV_X1    g749(.A(new_n907), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n925), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n284), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n257), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n935), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n914), .B2(new_n907), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n284), .A2(new_n262), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n939), .B(new_n865), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n623), .B1(new_n262), .B2(new_n938), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n845), .A2(new_n940), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n943), .A2(new_n945), .ZN(G57));
endmodule


