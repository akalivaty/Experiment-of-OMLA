//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n457), .A2(KEYINPUT65), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(KEYINPUT65), .B1(G567), .B2(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n462), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n464), .B2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n472), .A2(G137), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND3_X1  g053(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n473), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI22_X1  g057(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n475), .A2(new_n471), .A3(G2105), .A4(new_n465), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT67), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OR3_X1    g061(.A1(new_n484), .A2(KEYINPUT67), .A3(new_n485), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n475), .A2(new_n471), .A3(new_n490), .A4(new_n465), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n491), .A2(KEYINPUT4), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OR2_X1    g070(.A1(KEYINPUT68), .A2(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT68), .A2(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n473), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n484), .A2(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n494), .A2(new_n500), .ZN(G164));
  XOR2_X1   g076(.A(KEYINPUT5), .B(G543), .Z(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G651), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT6), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n502), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  XOR2_X1   g085(.A(KEYINPUT70), .B(G88), .Z(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n507), .B2(new_n509), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n502), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n503), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n512), .A2(new_n515), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n514), .A2(G51), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n510), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT5), .B(G543), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n525), .A2(new_n526), .A3(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n502), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n521), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n514), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n510), .A2(G90), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n540), .B1(new_n539), .B2(new_n538), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n502), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(new_n521), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT72), .ZN(new_n549));
  AOI22_X1  g124(.A1(G43), .A2(new_n514), .B1(new_n510), .B2(G81), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT6), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n519), .B2(new_n520), .ZN(new_n559));
  OAI21_X1  g134(.A(G543), .B1(new_n559), .B2(new_n508), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n507), .A2(new_n509), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n563), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n502), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n510), .A2(G91), .B1(new_n569), .B2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G168), .ZN(G286));
  NAND2_X1  g147(.A1(new_n514), .A2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n510), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n510), .A2(G86), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n502), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n530), .A2(KEYINPUT74), .A3(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(new_n521), .B1(G48), .B2(new_n514), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n578), .A2(new_n585), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n502), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(new_n521), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(G47), .A2(new_n514), .B1(new_n510), .B2(G85), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n510), .A2(G92), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT77), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n597), .A2(KEYINPUT77), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(KEYINPUT77), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n560), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(new_n560), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n530), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n505), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(new_n608), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n600), .A2(new_n603), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT80), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n596), .B1(new_n620), .B2(G868), .ZN(G284));
  XNOR2_X1  g196(.A(G284), .B(KEYINPUT81), .ZN(G321));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(G299), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(G168), .ZN(G297));
  OAI21_X1  g200(.A(new_n624), .B1(new_n623), .B2(G168), .ZN(G280));
  XNOR2_X1  g201(.A(KEYINPUT82), .B(G559), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n620), .B1(G860), .B2(new_n628), .ZN(G148));
  NAND2_X1  g204(.A1(new_n549), .A2(new_n550), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n623), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n619), .A2(new_n627), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(new_n623), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n484), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(G111), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(new_n479), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G135), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n492), .A2(new_n469), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT13), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(G2096), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n650), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2451), .B(G2454), .Z(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n665), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(KEYINPUT17), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n673), .B1(new_n675), .B2(new_n671), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT85), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  OR2_X1    g254(.A1(new_n670), .A2(new_n671), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n679), .C1(new_n675), .C2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2096), .B(G2100), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n689));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n686), .A2(new_n687), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n691), .B2(new_n688), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n691), .A2(KEYINPUT87), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT88), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n703), .A2(new_n705), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n685), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n708), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n710), .A2(new_n684), .A3(new_n706), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(G229));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G24), .ZN(new_n714));
  INV_X1    g289(.A(G290), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1986), .ZN(new_n717));
  INV_X1    g292(.A(G119), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n473), .A2(G107), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n720));
  OAI22_X1  g295(.A1(new_n484), .A2(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n642), .B2(G131), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT89), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G25), .B2(new_n725), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  AOI21_X1  g303(.A(new_n717), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n713), .A2(G6), .ZN(new_n730));
  INV_X1    g305(.A(G305), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n713), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT32), .B(G1981), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n713), .A2(G22), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT90), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n713), .ZN(new_n737));
  INV_X1    g312(.A(G1971), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n713), .A2(G23), .ZN(new_n740));
  INV_X1    g315(.A(G288), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(new_n713), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT33), .B(G1976), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n734), .A2(new_n739), .A3(new_n744), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n729), .B1(new_n727), .B2(new_n728), .C1(KEYINPUT34), .C2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(KEYINPUT34), .B2(new_n745), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n725), .A2(G32), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n642), .A2(G141), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT26), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n754), .A2(new_n755), .B1(G105), .B2(new_n469), .ZN(new_n756));
  INV_X1    g331(.A(G129), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n484), .B2(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n750), .B1(new_n760), .B2(new_n725), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT27), .B(G1996), .Z(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n764), .B2(KEYINPUT24), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(KEYINPUT24), .B2(new_n764), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n477), .B2(new_n725), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n713), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n713), .ZN(new_n772));
  INV_X1    g347(.A(G2072), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n492), .A2(G127), .ZN(new_n774));
  INV_X1    g349(.A(G115), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n462), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT93), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n473), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n777), .B2(new_n776), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n642), .B2(G139), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n725), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n725), .B2(G33), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n770), .B1(G1966), .B2(new_n772), .C1(new_n773), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n725), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  INV_X1    g364(.A(G128), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n473), .A2(G116), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  OAI22_X1  g367(.A1(new_n484), .A2(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n642), .B2(G140), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(new_n725), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2067), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT31), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G11), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(G11), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT30), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n800), .A2(G28), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n725), .B1(new_n800), .B2(G28), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n798), .B(new_n799), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n644), .B2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n713), .A2(G19), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n551), .B2(new_n713), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n804), .B1(new_n806), .B2(G1341), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n787), .A2(new_n796), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n725), .A2(G27), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n725), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT94), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G2078), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n713), .A2(G5), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G171), .B2(new_n713), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G1961), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n786), .A2(new_n773), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n772), .A2(G1966), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n761), .A2(new_n762), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n806), .A2(G1341), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n713), .A2(G20), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT23), .Z(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G299), .B2(G16), .ZN(new_n823));
  INV_X1    g398(.A(G1956), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n808), .A2(new_n812), .A3(new_n815), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n713), .A2(G4), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n620), .B2(new_n713), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1348), .ZN(new_n830));
  NOR2_X1   g405(.A1(G29), .A2(G35), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G162), .B2(G29), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G2090), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n827), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n749), .A2(new_n836), .ZN(G150));
  INV_X1    g412(.A(G150), .ZN(G311));
  NAND2_X1  g413(.A1(new_n510), .A2(G93), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n514), .A2(G55), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n504), .A2(new_n506), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  INV_X1    g420(.A(G559), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n847));
  OR3_X1    g422(.A1(new_n619), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n551), .B(new_n843), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n619), .B2(new_n846), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n848), .B2(new_n850), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT39), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT39), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n854), .A2(KEYINPUT97), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT97), .B1(new_n854), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(G145));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n760), .B(new_n784), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n722), .B(KEYINPUT100), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n648), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n860), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n500), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n865));
  AOI221_X4 g440(.A(new_n865), .B1(new_n492), .B2(new_n493), .C1(new_n491), .C2(KEYINPUT4), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n492), .A2(new_n493), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT99), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n864), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n794), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n642), .A2(G142), .ZN(new_n872));
  INV_X1    g447(.A(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n473), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  OAI221_X1 g450(.A(new_n872), .B1(new_n873), .B2(new_n484), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n871), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n863), .B(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n477), .B(KEYINPUT98), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(G162), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n644), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n878), .A2(KEYINPUT101), .A3(new_n881), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT101), .B1(new_n878), .B2(new_n881), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n859), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(G395));
  NAND2_X1  g462(.A1(new_n843), .A2(new_n623), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n630), .B(new_n843), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n632), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n849), .B1(new_n619), .B2(new_n627), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n614), .A2(KEYINPUT103), .A3(G299), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n612), .B1(new_n598), .B2(new_n599), .ZN(new_n894));
  OR2_X1    g469(.A1(G299), .A2(KEYINPUT103), .ZN(new_n895));
  NAND2_X1  g470(.A1(G299), .A2(KEYINPUT103), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n603), .A4(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n893), .A2(KEYINPUT41), .A3(new_n897), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT41), .B1(new_n893), .B2(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n892), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  XNOR2_X1  g479(.A(G288), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n715), .ZN(new_n906));
  XNOR2_X1  g481(.A(G288), .B(KEYINPUT104), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G290), .ZN(new_n908));
  NAND2_X1  g483(.A1(G305), .A2(G166), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n731), .A2(G303), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n906), .A2(new_n908), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n906), .A2(new_n908), .B1(new_n910), .B2(new_n909), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n911), .A3(KEYINPUT105), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n912), .A2(KEYINPUT42), .A3(new_n913), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n899), .B(new_n902), .C1(new_n920), .C2(KEYINPUT106), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n899), .A2(new_n902), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT106), .B1(new_n918), .B2(new_n919), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n921), .A2(new_n924), .B1(KEYINPUT106), .B2(new_n920), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n888), .B1(new_n925), .B2(new_n623), .ZN(G295));
  OAI21_X1  g501(.A(new_n888), .B1(new_n925), .B2(new_n623), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g504(.A1(G301), .A2(KEYINPUT107), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(new_n537), .C1(new_n541), .C2(new_n542), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n930), .A2(G168), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(G168), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n849), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n932), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G286), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n930), .A2(G168), .A3(new_n932), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n889), .A3(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n849), .B(KEYINPUT108), .C1(new_n933), .C2(new_n934), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n937), .A2(new_n898), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n900), .A2(new_n901), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n935), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n914), .A2(new_n916), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n948), .A2(new_n859), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n943), .A2(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n917), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n929), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n935), .A2(new_n941), .A3(new_n898), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n944), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n948), .B(new_n859), .C1(new_n955), .C2(new_n947), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n928), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n928), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n949), .A2(new_n929), .A3(new_n951), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n959), .A2(KEYINPUT109), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT109), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(G397));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(G1384), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n870), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n468), .A2(G2105), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n469), .A2(G101), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n476), .A3(G40), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT111), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n470), .A2(new_n971), .A3(G40), .A4(new_n476), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT112), .Z(new_n975));
  INV_X1    g550(.A(G2067), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n794), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT113), .ZN(new_n979));
  INV_X1    g554(.A(new_n975), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n760), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n974), .A2(G1996), .ZN(new_n982));
  OAI22_X1  g557(.A1(new_n981), .A2(new_n982), .B1(G1996), .B2(new_n760), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n722), .B(new_n728), .Z(new_n984));
  OAI211_X1 g559(.A(new_n979), .B(new_n983), .C1(new_n980), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n974), .ZN(new_n986));
  XNOR2_X1  g561(.A(G290), .B(G1986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n989));
  NAND2_X1  g564(.A1(G303), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  NAND4_X1  g568(.A1(G303), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(G8), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT118), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n494), .B2(new_n500), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT115), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n999), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n973), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n870), .A2(new_n1003), .A3(new_n998), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT114), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n870), .A2(new_n1006), .A3(new_n1003), .A4(new_n998), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1002), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G2090), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n997), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n970), .A2(new_n972), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1000), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n999), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1011), .A2(new_n1015), .A3(new_n997), .A4(new_n1009), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n999), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n973), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n738), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n996), .B(G8), .C1(new_n1010), .C2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1021), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1003), .B1(new_n870), .B2(new_n998), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1003), .B(new_n998), .C1(new_n494), .C2(new_n500), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n970), .A2(new_n972), .A3(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1025), .A2(new_n1027), .A3(G2090), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n995), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G305), .A2(G1981), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n700), .B1(new_n585), .B2(new_n577), .ZN(new_n1033));
  OR3_X1    g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n870), .A2(new_n970), .A3(new_n998), .A4(new_n972), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n741), .A2(G1976), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1023), .A2(new_n1030), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT125), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT125), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1023), .A2(new_n1046), .A3(new_n1049), .A4(new_n1030), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n999), .A2(new_n1018), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n870), .A2(new_n998), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n973), .B(new_n1051), .C1(new_n1052), .C2(KEYINPUT45), .ZN(new_n1053));
  INV_X1    g628(.A(G1966), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(G2084), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1057), .B2(G286), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1008), .A2(new_n768), .ZN(new_n1059));
  AOI21_X1  g634(.A(G168), .B1(new_n1059), .B2(new_n1055), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT51), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(G8), .C1(new_n1057), .C2(G286), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1020), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n1056), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(KEYINPUT53), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1053), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(G301), .B(KEYINPUT54), .ZN(new_n1072));
  INV_X1    g647(.A(new_n966), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n969), .A2(new_n1070), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1017), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1071), .A2(new_n1072), .B1(new_n1069), .B2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1048), .A2(new_n1050), .A3(new_n1064), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1348), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1035), .A2(G2067), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT121), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1080), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1082), .B(new_n1083), .C1(new_n1008), .C2(G1348), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT60), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1081), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n615), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1088), .B2(new_n615), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1086), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(G299), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT120), .B(new_n1095), .C1(new_n566), .C2(new_n570), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n824), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n973), .A2(new_n1017), .A3(new_n1019), .A4(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1094), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1096), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1098), .A2(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n1106));
  INV_X1    g681(.A(G1996), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n973), .A2(new_n1017), .A3(new_n1107), .A4(new_n1019), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1035), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1106), .B1(new_n1111), .B2(new_n551), .ZN(new_n1112));
  AOI211_X1 g687(.A(KEYINPUT59), .B(new_n630), .C1(new_n1108), .C2(new_n1110), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1105), .A2(KEYINPUT61), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1116), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT61), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1114), .A2(new_n1122), .A3(KEYINPUT123), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT61), .B1(new_n1126), .B2(new_n1120), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1119), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1104), .A2(new_n1116), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1130), .A4(new_n1120), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1124), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1123), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1088), .A2(new_n615), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT124), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1086), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1088), .A2(new_n1089), .A3(new_n615), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1092), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1129), .B(new_n1130), .C1(new_n1085), .C2(new_n614), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1120), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1078), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n741), .A2(new_n1042), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT119), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1036), .B1(new_n1145), .B2(new_n1031), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1023), .B2(new_n1045), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1057), .A2(G8), .A3(G168), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1023), .A2(new_n1046), .A3(new_n1030), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(G8), .B1(new_n1010), .B2(new_n1022), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n995), .ZN(new_n1153));
  AND4_X1   g728(.A1(KEYINPUT63), .A2(new_n1057), .A3(G8), .A4(G168), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1153), .A2(new_n1023), .A3(new_n1046), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1147), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1064), .A2(KEYINPUT62), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1061), .A2(new_n1158), .A3(new_n1063), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1071), .A2(G171), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1156), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n988), .B1(new_n1142), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n975), .B1(new_n759), .B2(new_n977), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT126), .Z(new_n1166));
  INV_X1    g741(.A(KEYINPUT47), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n982), .B(KEYINPUT46), .Z(new_n1168));
  AND3_X1   g743(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n974), .A2(G1986), .A3(G290), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT48), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n1169), .A2(new_n1170), .B1(new_n985), .B2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n983), .A2(new_n979), .A3(new_n724), .A4(new_n728), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n794), .A2(new_n976), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n980), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1164), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g753(.A1(G227), .A2(new_n460), .A3(G401), .ZN(new_n1180));
  NOR2_X1   g754(.A1(G229), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1181), .A2(new_n885), .ZN(new_n1182));
  NOR2_X1   g756(.A1(new_n952), .A2(new_n957), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n1183), .ZN(G308));
  OAI211_X1 g758(.A(new_n1181), .B(new_n885), .C1(new_n952), .C2(new_n957), .ZN(G225));
endmodule


