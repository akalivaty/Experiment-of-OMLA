//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT0), .B(G128), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G146), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n196), .A2(KEYINPUT0), .A3(G128), .A4(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI22_X1  g017(.A1(KEYINPUT66), .A2(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G134), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n201), .B1(new_n206), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n207), .A2(G134), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(new_n208), .B2(new_n210), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n203), .A2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n209), .A2(KEYINPUT11), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n219), .A3(KEYINPUT67), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(new_n220), .A3(G131), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n206), .A2(new_n212), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n205), .B(new_n204), .C1(new_n228), .C2(new_n208), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n229), .B2(new_n201), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n222), .A3(new_n220), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n226), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n227), .B1(new_n226), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n200), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n196), .A2(new_n197), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n238));
  INV_X1    g052(.A(new_n191), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n194), .B1(new_n239), .B2(new_n193), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n237), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n223), .A2(new_n224), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n216), .B2(new_n214), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n234), .A2(KEYINPUT30), .A3(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(G116), .B(G119), .Z(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n226), .A2(new_n200), .A3(new_n231), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n244), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT70), .B(G237), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(G210), .A3(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n256), .B(KEYINPUT27), .Z(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n244), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT68), .B1(new_n229), .B2(G131), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n220), .B2(new_n230), .ZN(new_n262));
  AND4_X1   g076(.A1(new_n222), .A2(new_n213), .A3(new_n220), .A4(G131), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT69), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n226), .A2(new_n227), .A3(new_n231), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n260), .B1(new_n266), .B2(new_n200), .ZN(new_n267));
  INV_X1    g081(.A(new_n248), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n259), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n253), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n253), .B2(new_n269), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n250), .A2(new_n248), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n267), .B2(new_n268), .ZN(new_n276));
  AND4_X1   g090(.A1(new_n275), .A2(new_n234), .A3(new_n268), .A4(new_n244), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n259), .ZN(new_n279));
  AOI211_X1 g093(.A(KEYINPUT32), .B(new_n189), .C1(new_n273), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n253), .A2(new_n269), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT31), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n253), .A2(new_n269), .A3(new_n270), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n285), .B2(new_n188), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G472), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n234), .A2(new_n268), .A3(new_n244), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(KEYINPUT28), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  INV_X1    g105(.A(new_n259), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n274), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n292), .B(new_n274), .C1(new_n276), .C2(new_n277), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT71), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n253), .A2(new_n289), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n296), .B2(new_n259), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n276), .A2(new_n277), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n267), .A2(new_n268), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n292), .A2(KEYINPUT29), .ZN(new_n302));
  AOI21_X1  g116(.A(G902), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n288), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n187), .B1(new_n287), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G116), .B(G122), .ZN(new_n306));
  INV_X1    g120(.A(G107), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n193), .A2(G128), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT13), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n235), .A2(G143), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n309), .A2(new_n310), .ZN(new_n314));
  OAI21_X1  g128(.A(G134), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(new_n312), .A3(new_n203), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT9), .B(G234), .ZN(new_n318));
  INV_X1    g132(.A(G217), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n318), .A2(new_n319), .A3(G953), .ZN(new_n320));
  INV_X1    g134(.A(G116), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G122), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT14), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n321), .A2(G122), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n324), .B2(KEYINPUT14), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n325), .B2(KEYINPUT94), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(KEYINPUT94), .B2(new_n325), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n327), .A2(G107), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n306), .A2(new_n307), .ZN(new_n329));
  INV_X1    g143(.A(new_n316), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n203), .B1(new_n309), .B2(new_n312), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n317), .B(new_n320), .C1(new_n328), .C2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n320), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n327), .B2(G107), .ZN(new_n335));
  INV_X1    g149(.A(new_n317), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(G902), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT95), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n338), .A2(new_n339), .ZN(new_n342));
  INV_X1    g156(.A(G478), .ZN(new_n343));
  OAI22_X1  g157(.A1(new_n341), .A2(new_n342), .B1(KEYINPUT15), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(G234), .A2(G237), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n345), .A2(G952), .A3(new_n255), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n345), .A2(G902), .A3(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT21), .B(G898), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT15), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n340), .A2(new_n351), .A3(G478), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n344), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(G475), .A2(G902), .ZN(new_n354));
  XNOR2_X1  g168(.A(G113), .B(G122), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n254), .A2(G214), .A3(new_n255), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(new_n193), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G131), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(G143), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n224), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT92), .ZN(new_n364));
  XNOR2_X1  g178(.A(G125), .B(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT16), .ZN(new_n366));
  INV_X1    g180(.A(G125), .ZN(new_n367));
  OR3_X1    g181(.A1(new_n367), .A2(KEYINPUT16), .A3(G140), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(G146), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n360), .A2(new_n362), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n365), .B(KEYINPUT19), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n191), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n364), .A2(new_n369), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT18), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(new_n224), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n191), .A2(new_n365), .ZN(new_n378));
  INV_X1    g192(.A(G146), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n365), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n361), .A2(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n361), .A2(KEYINPUT91), .A3(new_n377), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n359), .B2(new_n376), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n357), .B1(new_n374), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n361), .A2(new_n224), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n366), .A2(new_n368), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n379), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(new_n369), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n388), .B(new_n391), .C1(new_n363), .C2(KEYINPUT17), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n357), .B(KEYINPUT93), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n392), .A2(new_n385), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n354), .B1(new_n386), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT20), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n397), .B(new_n354), .C1(new_n386), .C2(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G902), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n392), .A2(new_n385), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(new_n357), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G475), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n353), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n196), .A2(new_n197), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n407));
  OAI21_X1  g221(.A(G128), .B1(new_n194), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n237), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n356), .A2(G107), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n356), .A2(G107), .ZN(new_n413));
  OAI21_X1  g227(.A(G101), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT3), .B1(new_n356), .B2(G107), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n307), .A3(G104), .ZN(new_n417));
  INV_X1    g231(.A(G101), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n415), .A2(new_n417), .A3(new_n418), .A4(new_n411), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n410), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT10), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n420), .B1(new_n409), .B2(new_n237), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n426), .B2(KEYINPUT10), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n420), .A2(new_n423), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n241), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n241), .A2(KEYINPUT84), .A3(new_n428), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n424), .A2(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n415), .A2(new_n417), .A3(new_n411), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G101), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n419), .A2(KEYINPUT4), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n438), .A3(G101), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT82), .A4(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n435), .A2(KEYINPUT4), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n200), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n433), .A2(new_n264), .A3(new_n265), .A4(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G140), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n255), .A2(G227), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n447), .A2(KEYINPUT85), .A3(new_n451), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n433), .A2(new_n446), .B1(new_n264), .B2(new_n265), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n450), .B(KEYINPUT80), .Z(new_n459));
  INV_X1    g273(.A(new_n447), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n422), .B1(new_n241), .B2(new_n421), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT12), .B1(new_n266), .B2(new_n461), .ZN(new_n462));
  AND4_X1   g276(.A1(KEYINPUT12), .A2(new_n461), .A3(new_n226), .A4(new_n231), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n459), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(G469), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G469), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n447), .B(new_n451), .C1(new_n462), .C2(new_n463), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n451), .B1(new_n457), .B2(new_n447), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n467), .B(new_n400), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n467), .A2(new_n400), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G221), .B1(new_n318), .B2(G902), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT78), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT79), .Z(new_n477));
  NAND3_X1  g291(.A1(new_n405), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT5), .ZN(new_n479));
  INV_X1    g293(.A(G119), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n480), .A3(G116), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT87), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n482), .B(G113), .C1(new_n479), .C2(new_n246), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n246), .A2(new_n247), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n421), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n445), .A2(new_n248), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n486), .B1(new_n444), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G110), .B(G122), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT88), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n487), .B1(new_n442), .B2(new_n443), .ZN(new_n493));
  INV_X1    g307(.A(new_n490), .ZN(new_n494));
  NOR4_X1   g308(.A1(new_n493), .A2(new_n486), .A3(KEYINPUT88), .A4(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n241), .A2(G125), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n199), .A2(G125), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT89), .B(G224), .Z(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G953), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n490), .B(KEYINPUT8), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n421), .B1(new_n483), .B2(new_n484), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n506), .B1(new_n486), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n500), .A2(new_n504), .A3(new_n502), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n497), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n500), .B(new_n502), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n489), .A2(KEYINPUT6), .A3(new_n490), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n489), .B2(new_n490), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(new_n495), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT6), .B1(new_n489), .B2(new_n490), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n513), .B(new_n514), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G210), .B1(G237), .B2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n512), .A2(new_n519), .A3(new_n521), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n526));
  OAI21_X1  g340(.A(G214), .B1(G237), .B2(G902), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT86), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n512), .A2(new_n519), .A3(new_n521), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n521), .B1(new_n512), .B2(new_n519), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT90), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n478), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n298), .A2(new_n303), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G472), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n537), .B(KEYINPUT72), .C1(new_n286), .C2(new_n280), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT22), .B(G137), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT74), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT74), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n541), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n543), .B1(new_n541), .B2(new_n547), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n390), .A2(new_n369), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n480), .B2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n553), .B(new_n554), .C1(G119), .C2(new_n235), .ZN(new_n555));
  XNOR2_X1  g369(.A(G119), .B(G128), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT24), .B(G110), .Z(new_n557));
  AOI22_X1  g371(.A1(new_n555), .A2(G110), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n369), .A2(new_n378), .ZN(new_n560));
  OAI22_X1  g374(.A1(new_n555), .A2(G110), .B1(new_n556), .B2(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT76), .B1(new_n550), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n547), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n542), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n541), .A2(new_n543), .A3(new_n547), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n551), .A2(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT76), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(new_n569), .B2(new_n570), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n563), .A2(KEYINPUT75), .A3(new_n568), .A4(new_n567), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n577), .A3(new_n400), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT25), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n573), .A2(new_n577), .A3(new_n580), .A4(new_n400), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n319), .B1(G234), .B2(new_n400), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT77), .ZN(new_n584));
  OR3_X1    g398(.A1(new_n578), .A2(new_n584), .A3(new_n582), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n584), .B1(new_n578), .B2(new_n582), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n305), .A2(new_n535), .A3(new_n538), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  AND3_X1   g403(.A1(new_n474), .A2(new_n587), .A3(new_n477), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n285), .A2(new_n400), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n591), .A2(G472), .B1(new_n188), .B2(new_n285), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n525), .A2(new_n527), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n399), .A2(new_n404), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n333), .A2(new_n337), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n333), .A2(new_n337), .A3(KEYINPUT96), .A4(new_n599), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n343), .A2(G902), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n604), .A2(KEYINPUT97), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT97), .B1(new_n604), .B2(new_n605), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n338), .A2(G478), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n597), .A2(new_n610), .A3(new_n350), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n596), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT34), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  AOI22_X1  g428(.A1(new_n396), .A2(new_n398), .B1(new_n403), .B2(G475), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n344), .A2(new_n352), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n350), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n596), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT98), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT35), .B(G107), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  NAND2_X1  g435(.A1(new_n534), .A2(new_n530), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n405), .A2(new_n474), .A3(new_n477), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n569), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n570), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n569), .A2(new_n625), .A3(new_n563), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n582), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n400), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n578), .B2(KEYINPUT25), .ZN(new_n633));
  AOI211_X1 g447(.A(new_n624), .B(new_n632), .C1(new_n633), .C2(new_n581), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT99), .B1(new_n583), .B2(new_n631), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n622), .A2(new_n623), .A3(new_n592), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n474), .A3(new_n477), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n347), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n346), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n615), .A2(new_n616), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n640), .A2(new_n594), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n305), .A2(new_n538), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  NAND2_X1  g462(.A1(new_n296), .A2(new_n292), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  INV_X1    g464(.A(new_n289), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n292), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n649), .B(new_n650), .C1(new_n300), .C2(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n300), .A2(new_n651), .A3(new_n292), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n259), .B1(new_n253), .B2(new_n289), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT100), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n654), .A2(new_n400), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(KEYINPUT101), .A3(G472), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n659), .B1(new_n286), .B2(new_n280), .ZN(new_n660));
  AOI21_X1  g474(.A(KEYINPUT101), .B1(new_n658), .B2(G472), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n399), .A2(new_n404), .B1(new_n344), .B2(new_n352), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n583), .A2(new_n631), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n664), .A2(new_n527), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n644), .B(KEYINPUT39), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n474), .A2(new_n477), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n667), .B1(new_n669), .B2(KEYINPUT40), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n525), .B(KEYINPUT38), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n663), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT102), .B(G143), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G45));
  NAND3_X1  g489(.A1(new_n597), .A2(new_n610), .A3(new_n644), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n640), .A2(new_n594), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n305), .A2(new_n538), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT103), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n305), .A2(new_n677), .A3(new_n538), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  OAI21_X1  g497(.A(new_n450), .B1(new_n460), .B2(new_n456), .ZN(new_n684));
  AOI21_X1  g498(.A(G902), .B1(new_n684), .B2(new_n468), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n467), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n476), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n685), .A2(new_n688), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(new_n594), .A3(new_n611), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n305), .A2(new_n538), .A3(new_n587), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NOR3_X1   g510(.A1(new_n692), .A2(new_n594), .A3(new_n617), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n305), .A2(new_n538), .A3(new_n587), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT105), .B(G116), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G18));
  NOR2_X1   g514(.A1(new_n692), .A2(new_n594), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n636), .A2(new_n405), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n305), .A2(new_n538), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  NAND3_X1  g518(.A1(new_n525), .A2(new_n664), .A3(new_n527), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n692), .A3(new_n349), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n259), .B1(new_n299), .B2(new_n300), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n189), .B1(new_n273), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n591), .B2(G472), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n587), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  AND2_X1   g525(.A1(new_n709), .A2(new_n665), .ZN(new_n712));
  INV_X1    g526(.A(new_n644), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n615), .A2(new_n609), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n714), .A3(new_n701), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT106), .B(G125), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G27));
  NAND2_X1  g531(.A1(new_n474), .A2(new_n690), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n718), .A2(new_n719), .A3(new_n676), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n305), .A2(new_n538), .A3(new_n587), .A4(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n286), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n285), .A2(new_n281), .A3(new_n188), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n304), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n472), .B1(new_n685), .B2(new_n467), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n476), .B1(new_n727), .B2(new_n466), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n729), .A4(new_n714), .ZN(new_n730));
  INV_X1    g544(.A(new_n587), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n726), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT107), .B1(new_n723), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n735), .B(new_n732), .C1(new_n721), .C2(new_n722), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NOR3_X1   g552(.A1(new_n718), .A2(new_n719), .A3(new_n645), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n305), .A2(new_n538), .A3(new_n587), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  AND2_X1   g555(.A1(new_n458), .A2(new_n465), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n742), .B2(KEYINPUT45), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n458), .A2(KEYINPUT45), .A3(new_n465), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT46), .B1(new_n746), .B2(new_n473), .ZN(new_n747));
  INV_X1    g561(.A(new_n471), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n473), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n476), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n668), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n610), .A2(new_n615), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT108), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n592), .A2(new_n666), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n758), .A2(KEYINPUT44), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n719), .B1(new_n758), .B2(KEYINPUT44), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n752), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT109), .B(G137), .Z(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G39));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n751), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n305), .A2(new_n538), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n731), .A3(new_n714), .A4(new_n729), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(G140), .Z(G42));
  NAND2_X1  g583(.A1(new_n689), .A2(new_n691), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n765), .B1(new_n477), .B2(new_n770), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n587), .A2(new_n755), .A3(new_n346), .A4(new_n709), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n729), .A3(new_n772), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n692), .A2(new_n731), .A3(new_n719), .A4(new_n643), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n662), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n615), .A2(new_n609), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n672), .A2(new_n527), .A3(new_n692), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT50), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n755), .A2(new_n346), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n692), .A3(new_n719), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n777), .B(new_n780), .C1(new_n712), .C2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n773), .A2(KEYINPUT51), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n773), .B2(new_n783), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n597), .A2(new_n610), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n775), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n726), .A2(new_n731), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT48), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT115), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(KEYINPUT115), .ZN(new_n792));
  OR3_X1    g606(.A1(new_n789), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n791), .ZN(new_n794));
  INV_X1    g608(.A(G952), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n795), .B(G953), .C1(new_n772), .C2(new_n701), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  OR4_X1    g611(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n611), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n526), .B1(new_n525), .B2(new_n529), .ZN(new_n800));
  AOI211_X1 g614(.A(KEYINPUT90), .B(new_n528), .C1(new_n523), .C2(new_n524), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n622), .A2(KEYINPUT110), .A3(new_n799), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n593), .A3(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(new_n694), .A3(new_n698), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n588), .A2(new_n703), .A3(new_n710), .ZN(new_n808));
  INV_X1    g622(.A(new_n617), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n622), .A2(new_n592), .A3(new_n590), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n637), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT111), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n637), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n615), .A2(new_n344), .A3(new_n352), .A4(new_n644), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n640), .A2(new_n816), .A3(new_n719), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n305), .A2(new_n817), .A3(new_n538), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n712), .A2(new_n714), .A3(new_n729), .A4(new_n728), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n740), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n807), .A2(new_n808), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n734), .A3(new_n736), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n644), .B(KEYINPUT113), .Z(new_n824));
  NAND2_X1  g638(.A1(new_n666), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n705), .A2(new_n718), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n660), .B2(new_n661), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n647), .A2(new_n715), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n682), .A2(new_n823), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n647), .A2(new_n715), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT112), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n647), .A2(new_n832), .A3(new_n715), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n682), .A2(new_n831), .A3(new_n827), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n829), .B1(KEYINPUT52), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n822), .B2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n807), .A2(new_n808), .A3(new_n815), .A4(new_n820), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n682), .A2(new_n828), .A3(new_n823), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n682), .A2(new_n828), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT52), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n737), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n836), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n842), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n723), .A2(new_n733), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n821), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n835), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n844), .B1(KEYINPUT54), .B2(new_n850), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n798), .A2(new_n851), .B1(G952), .B2(G953), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n770), .A2(KEYINPUT49), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n770), .A2(KEYINPUT49), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n587), .A2(new_n529), .A3(new_n477), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n753), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n672), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n662), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n852), .A2(new_n858), .ZN(G75));
  NOR2_X1   g673(.A1(new_n255), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n841), .A2(new_n842), .B1(new_n835), .B2(new_n848), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n400), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n863), .B2(G210), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT116), .Z(new_n866));
  XNOR2_X1  g680(.A(new_n513), .B(KEYINPUT55), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT117), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n866), .B(new_n868), .Z(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n861), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n850), .A2(G902), .ZN(new_n873));
  INV_X1    g687(.A(G210), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT118), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n860), .B1(new_n875), .B2(new_n869), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n864), .A2(new_n870), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n881), .ZN(G51));
  XNOR2_X1  g696(.A(new_n850), .B(KEYINPUT54), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n472), .B(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n470), .B2(new_n469), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n863), .A2(new_n745), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n860), .B1(new_n886), .B2(new_n887), .ZN(G54));
  NAND2_X1  g702(.A1(KEYINPUT58), .A2(G475), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT119), .Z(new_n890));
  NOR2_X1   g704(.A1(new_n873), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n386), .A2(new_n394), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n861), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT120), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n891), .A2(new_n892), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n861), .A4(new_n893), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n896), .A2(new_n899), .ZN(G60));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT59), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n883), .A2(new_n604), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n604), .B1(new_n851), .B2(new_n903), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n904), .A2(new_n860), .A3(new_n905), .ZN(G63));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n907));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT60), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n842), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n823), .B1(new_n682), .B2(new_n828), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n829), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n822), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n848), .A2(new_n838), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n910), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n573), .A2(new_n577), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT122), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n860), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n629), .B(new_n910), .C1(new_n914), .C2(new_n916), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n907), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n919), .B1(new_n862), .B2(new_n909), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n907), .A2(new_n923), .A3(new_n861), .A4(new_n921), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n909), .B1(new_n845), .B2(new_n849), .ZN(new_n926));
  INV_X1    g740(.A(new_n919), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n861), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n922), .A2(new_n924), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n861), .B1(new_n926), .B2(new_n927), .ZN(new_n932));
  INV_X1    g746(.A(new_n921), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT123), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n923), .A2(new_n921), .A3(new_n907), .A4(new_n861), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n934), .A2(new_n935), .B1(new_n929), .B2(new_n928), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n931), .A2(new_n936), .ZN(G66));
  NOR2_X1   g751(.A1(new_n501), .A2(new_n348), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n255), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n807), .A2(new_n808), .A3(new_n815), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n255), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n866), .B1(G898), .B2(new_n255), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(G69));
  AOI21_X1  g757(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n255), .A2(G900), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n245), .A2(new_n252), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n372), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n761), .B1(new_n765), .B2(new_n767), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n752), .A2(new_n595), .A3(new_n664), .A4(new_n788), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n740), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n682), .A2(new_n831), .A3(new_n833), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n952), .A2(new_n737), .A3(new_n953), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n946), .B(new_n948), .C1(new_n954), .C2(new_n255), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n766), .A2(new_n731), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n615), .A2(new_n616), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n719), .B(new_n669), .C1(new_n786), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n949), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n953), .A2(new_n673), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n948), .A2(new_n255), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(KEYINPUT125), .B(new_n945), .C1(new_n955), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n954), .A2(new_n255), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n948), .A2(new_n946), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n963), .A2(new_n964), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n966), .A2(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n963), .B2(new_n940), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n656), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n954), .B2(new_n940), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n652), .A2(new_n253), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT126), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n836), .A2(new_n843), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n649), .A2(new_n976), .A3(new_n980), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR4_X1   g799(.A1(new_n978), .A2(new_n982), .A3(new_n860), .A4(new_n985), .ZN(G57));
endmodule


