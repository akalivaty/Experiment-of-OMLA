//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT11), .B(G169gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G15gat), .B(G22gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G1gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT16), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT88), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n213), .A2(KEYINPUT88), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n216), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n209), .A2(new_n212), .A3(new_n218), .A4(new_n214), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT87), .B(G36gat), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G29gat), .A2(G36gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT14), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n221), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT14), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n225), .B(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n229), .B(KEYINPUT15), .C1(new_n223), .C2(new_n222), .ZN(new_n230));
  XNOR2_X1  g029(.A(G43gat), .B(G50gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n224), .A2(new_n226), .ZN(new_n233));
  INV_X1    g032(.A(new_n231), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT15), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n232), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n232), .B2(new_n235), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n220), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(new_n235), .ZN(new_n241));
  AOI211_X1 g040(.A(KEYINPUT88), .B(new_n213), .C1(new_n209), .C2(new_n212), .ZN(new_n242));
  INV_X1    g041(.A(new_n219), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n240), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n239), .A2(KEYINPUT18), .A3(new_n240), .A4(new_n245), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n220), .A2(new_n232), .A3(new_n235), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT90), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n245), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n240), .B(KEYINPUT13), .Z(new_n255));
  NAND3_X1  g054(.A1(new_n241), .A2(new_n244), .A3(KEYINPUT90), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n254), .A2(KEYINPUT91), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT91), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n256), .ZN(new_n260));
  INV_X1    g059(.A(new_n255), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT89), .A3(new_n247), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n250), .A2(new_n258), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n258), .A2(new_n262), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n207), .B1(new_n247), .B2(new_n246), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n207), .A2(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G113gat), .ZN(new_n268));
  INV_X1    g067(.A(G120gat), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(new_n268), .B2(new_n269), .ZN(new_n271));
  XNOR2_X1  g070(.A(G127gat), .B(G134gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n270), .B(new_n272), .C1(new_n277), .C2(new_n268), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n274), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n274), .B2(new_n278), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283));
  INV_X1    g082(.A(G155gat), .ZN(new_n284));
  INV_X1    g083(.A(G162gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G141gat), .B(G148gat), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n283), .B(new_n286), .C1(new_n287), .C2(KEYINPUT2), .ZN(new_n288));
  INV_X1    g087(.A(G141gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G148gat), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G141gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(new_n283), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n283), .A2(KEYINPUT2), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT76), .B1(new_n288), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n288), .A2(KEYINPUT76), .A3(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT4), .B1(new_n282), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n288), .A2(new_n296), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(new_n274), .A3(new_n278), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n274), .A2(new_n278), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n296), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(KEYINPUT3), .ZN(new_n309));
  OAI22_X1  g108(.A1(new_n302), .A2(new_n304), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR4_X1   g111(.A1(new_n301), .A2(new_n310), .A3(KEYINPUT5), .A4(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G57gat), .B(G85gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT79), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G1gat), .B(G29gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT70), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n274), .A2(new_n278), .A3(new_n279), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n288), .A2(KEYINPUT76), .A3(new_n296), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n297), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n322), .B(KEYINPUT4), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n328), .B(new_n311), .C1(new_n306), .C2(new_n309), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n302), .B1(new_n282), .B2(new_n300), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT77), .B1(new_n304), .B2(KEYINPUT4), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n303), .B(new_n307), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT5), .B1(new_n334), .B2(new_n311), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n314), .B(new_n321), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n330), .A2(new_n331), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n311), .B1(new_n306), .B2(new_n309), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n330), .B2(new_n322), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n320), .B1(new_n340), .B2(new_n313), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n336), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT6), .B(new_n320), .C1(new_n340), .C2(new_n313), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n346), .B(KEYINPUT74), .Z(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G169gat), .ZN(new_n349));
  INV_X1    g148(.A(G176gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT66), .ZN(new_n352));
  OAI22_X1  g151(.A1(new_n349), .A2(new_n350), .B1(new_n352), .B2(KEYINPUT23), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n352), .A2(KEYINPUT23), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G183gat), .ZN(new_n359));
  INV_X1    g158(.A(G190gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT23), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n355), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT25), .ZN(new_n367));
  AND2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT26), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(new_n364), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT68), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n351), .B2(KEYINPUT26), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n364), .A2(KEYINPUT68), .A3(new_n369), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT27), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G183gat), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n360), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n377), .A3(new_n360), .ZN(new_n381));
  INV_X1    g180(.A(new_n379), .ZN(new_n382));
  NAND2_X1  g181(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n374), .A2(new_n380), .A3(new_n356), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n358), .A2(KEYINPUT64), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT64), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n356), .A2(new_n387), .A3(new_n357), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n386), .A2(new_n361), .A3(new_n362), .A4(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n365), .A2(KEYINPUT65), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT25), .B1(new_n365), .B2(KEYINPUT65), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n389), .A2(new_n355), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n367), .A2(new_n385), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n348), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G197gat), .B(G204gat), .ZN(new_n397));
  INV_X1    g196(.A(G218gat), .ZN(new_n398));
  INV_X1    g197(.A(G211gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT72), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT72), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G211gat), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n398), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n397), .B1(new_n403), .B2(KEYINPUT22), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n399), .A2(G218gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n398), .A2(G211gat), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT73), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n398), .A2(G211gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n399), .A2(G218gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT73), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT22), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT72), .B(G211gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n398), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n416), .A2(new_n397), .A3(new_n407), .A4(new_n411), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n393), .A2(new_n348), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(new_n419), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n395), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT75), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n420), .A2(new_n423), .A3(KEYINPUT30), .A4(new_n427), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n430), .B1(new_n429), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n418), .B1(new_n396), .B2(new_n419), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n422), .A2(new_n395), .A3(new_n421), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n427), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n345), .A2(new_n434), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n303), .A2(new_n305), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n418), .B1(new_n442), .B2(new_n394), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G228gat), .ZN(new_n445));
  INV_X1    g244(.A(G233gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT3), .B1(new_n418), .B2(new_n394), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n444), .B(new_n447), .C1(new_n303), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT81), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n413), .B2(new_n417), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n327), .B1(new_n451), .B2(KEYINPUT3), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n443), .B1(new_n452), .B2(KEYINPUT80), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n327), .B(new_n454), .C1(new_n451), .C2(KEYINPUT3), .ZN(new_n455));
  AOI211_X1 g254(.A(new_n450), .B(new_n447), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT80), .B1(new_n448), .B2(new_n300), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n455), .A3(new_n444), .ZN(new_n458));
  INV_X1    g257(.A(new_n447), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT81), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n449), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G22gat), .ZN(new_n462));
  INV_X1    g261(.A(G22gat), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n463), .B(new_n449), .C1(new_n456), .C2(new_n460), .ZN(new_n464));
  XNOR2_X1  g263(.A(G78gat), .B(G106gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT31), .B(G50gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n458), .A2(new_n459), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n450), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n458), .A2(KEYINPUT81), .A3(new_n459), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n463), .B1(new_n473), .B2(new_n449), .ZN(new_n474));
  INV_X1    g273(.A(new_n464), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n441), .A2(new_n468), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G43gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(G71gat), .B(G99gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G227gat), .A2(G233gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n393), .A2(new_n325), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n393), .A2(new_n325), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n486), .B2(KEYINPUT32), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT71), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n282), .A2(new_n367), .A3(new_n385), .A4(new_n392), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n393), .A2(new_n325), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n482), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n488), .B1(new_n491), .B2(KEYINPUT33), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT33), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n486), .A2(KEYINPUT71), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n486), .B(KEYINPUT32), .C1(new_n493), .C2(new_n481), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n490), .ZN(new_n498));
  OR3_X1    g297(.A1(new_n498), .A2(KEYINPUT34), .A3(new_n483), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT34), .B1(new_n498), .B2(new_n483), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n495), .A2(new_n500), .A3(new_n499), .A4(new_n496), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n477), .A2(new_n478), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n478), .B1(new_n477), .B2(new_n508), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n476), .A2(new_n468), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n312), .B1(new_n301), .B2(new_n310), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT39), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n334), .B2(new_n311), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT40), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n512), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n513), .B(new_n312), .C1(new_n301), .C2(new_n310), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT83), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n321), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n321), .B2(new_n518), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n515), .B2(new_n516), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n429), .A2(new_n431), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n440), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n515), .A2(new_n516), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n517), .B(new_n526), .C1(new_n520), .C2(new_n521), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n523), .A2(new_n525), .A3(new_n341), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT38), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n428), .B1(new_n424), .B2(KEYINPUT37), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(KEYINPUT85), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT37), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n427), .B1(new_n437), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n424), .A2(KEYINPUT37), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n343), .A2(new_n344), .A3(new_n438), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n532), .A2(new_n536), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n529), .A2(new_n540), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n509), .A2(new_n510), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n502), .A2(new_n503), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n467), .B1(new_n462), .B2(new_n464), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548));
  INV_X1    g347(.A(new_n525), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n345), .A4(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n511), .A2(KEYINPUT86), .A3(new_n543), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n441), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n550), .B1(new_n554), .B2(new_n548), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n267), .B1(new_n542), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(KEYINPUT41), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT7), .ZN(new_n563));
  NOR2_X1   g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(KEYINPUT8), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G99gat), .ZN(new_n568));
  INV_X1    g367(.A(G106gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n565), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n563), .A2(new_n572), .A3(new_n566), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n241), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n557), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n237), .A2(new_n238), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT98), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n580), .B(new_n576), .C1(new_n577), .C2(new_n575), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n579), .B2(new_n581), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n561), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n560), .A3(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G71gat), .B(G78gat), .Z(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  INV_X1    g392(.A(G71gat), .ZN(new_n594));
  INV_X1    g393(.A(G78gat), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n592), .B1(KEYINPUT94), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(G57gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT93), .B(G57gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(new_n598), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n596), .A2(KEYINPUT94), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G57gat), .B(G64gat), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n604), .A2(KEYINPUT92), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n596), .B1(new_n604), .B2(KEYINPUT92), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n592), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n244), .B1(KEYINPUT21), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT97), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT95), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n611), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n609), .A2(KEYINPUT21), .ZN(new_n618));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n591), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n574), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n603), .A2(new_n607), .A3(new_n573), .A4(new_n571), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(KEYINPUT99), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n630), .A3(new_n575), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n632), .B2(new_n635), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n633), .B(KEYINPUT100), .Z(new_n638));
  OAI21_X1  g437(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT101), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n639), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT10), .B1(new_n629), .B2(new_n631), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n633), .B1(new_n649), .B2(new_n636), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n642), .A3(new_n634), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n626), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n556), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n345), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n211), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n654), .A2(new_n549), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n213), .B2(new_n657), .ZN(new_n660));
  MUX2_X1   g459(.A(new_n659), .B(new_n660), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g460(.A(G15gat), .B1(new_n654), .B2(new_n508), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n504), .A2(G15gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n654), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT102), .Z(G1326gat));
  NOR2_X1   g464(.A1(new_n654), .A2(new_n511), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT43), .B(G22gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  NAND2_X1  g467(.A1(new_n264), .A2(new_n207), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n266), .A2(new_n258), .A3(new_n262), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n652), .ZN(new_n672));
  INV_X1    g471(.A(new_n625), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n591), .ZN(new_n675));
  INV_X1    g474(.A(new_n345), .ZN(new_n676));
  NOR4_X1   g475(.A1(new_n546), .A2(KEYINPUT35), .A3(new_n676), .A4(new_n525), .ZN(new_n677));
  INV_X1    g476(.A(new_n441), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n546), .A2(new_n551), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT86), .B1(new_n511), .B2(new_n543), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n681), .B2(KEYINPUT35), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n509), .A2(new_n510), .A3(new_n541), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n671), .B(new_n675), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n223), .A3(new_n676), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT45), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n590), .A2(KEYINPUT44), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n682), .B2(new_n683), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n267), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT103), .Z(new_n691));
  OAI211_X1 g490(.A(new_n477), .B(new_n508), .C1(new_n529), .C2(new_n540), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n591), .B1(new_n555), .B2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n689), .B(new_n691), .C1(new_n693), .C2(KEYINPUT44), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n345), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n687), .A2(new_n695), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n685), .A2(new_n222), .A3(new_n525), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT46), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(KEYINPUT46), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n694), .A2(new_n549), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n698), .B(new_n699), .C1(new_n222), .C2(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702));
  OAI21_X1  g501(.A(G43gat), .B1(new_n694), .B2(new_n508), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n684), .A2(G43gat), .A3(new_n504), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1330gat));
  NOR2_X1   g506(.A1(new_n511), .A2(G50gat), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT108), .B1(new_n684), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n556), .A2(new_n711), .A3(new_n675), .A4(new_n708), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n710), .A2(new_n712), .A3(KEYINPUT48), .ZN(new_n713));
  OAI21_X1  g512(.A(G50gat), .B1(new_n694), .B2(new_n511), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n713), .A2(KEYINPUT109), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT109), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n684), .B2(new_n709), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n685), .A2(KEYINPUT107), .A3(new_n708), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n714), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n715), .A2(new_n716), .B1(new_n720), .B2(new_n721), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n555), .A2(new_n692), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n626), .A2(new_n671), .A3(new_n672), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT110), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n676), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n600), .ZN(G1332gat));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n725), .B(new_n729), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n730), .A2(new_n549), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT49), .B(G64gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n726), .A2(new_n525), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1333gat));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n504), .A2(G71gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n726), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n508), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n594), .B1(new_n726), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n735), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G71gat), .B1(new_n730), .B2(new_n508), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(KEYINPUT50), .A3(new_n737), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1334gat));
  INV_X1    g543(.A(new_n511), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g546(.A1(new_n625), .A2(new_n671), .ZN(new_n748));
  AND4_X1   g547(.A1(KEYINPUT51), .A2(new_n723), .A3(new_n590), .A4(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT51), .B1(new_n693), .B2(new_n748), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR4_X1    g550(.A1(G85gat), .A2(new_n751), .A3(new_n345), .A4(new_n672), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n748), .A2(new_n652), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n689), .B(new_n753), .C1(new_n693), .C2(KEYINPUT44), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n345), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(G1336gat));
  NOR2_X1   g555(.A1(new_n549), .A2(G92gat), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n652), .B(new_n757), .C1(new_n749), .C2(new_n750), .ZN(new_n758));
  OAI21_X1  g557(.A(G92gat), .B1(new_n754), .B2(new_n549), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(KEYINPUT111), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n761), .A3(KEYINPUT52), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n758), .B(new_n759), .C1(KEYINPUT111), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n754), .B2(new_n508), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n652), .A2(new_n568), .A3(new_n543), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT112), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n751), .B2(new_n768), .ZN(G1338gat));
  OAI21_X1  g568(.A(G106gat), .B1(new_n754), .B2(new_n511), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n745), .A2(new_n569), .A3(new_n652), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n770), .B(new_n771), .C1(new_n751), .C2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n772), .B(KEYINPUT113), .Z(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n749), .B2(new_n750), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT114), .B1(new_n776), .B2(KEYINPUT53), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n778), .B(new_n771), .C1(new_n770), .C2(new_n775), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n773), .B1(new_n777), .B2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781));
  INV_X1    g580(.A(new_n651), .ZN(new_n782));
  INV_X1    g581(.A(new_n638), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n783), .B(new_n784), .C1(new_n649), .C2(new_n636), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n643), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n650), .A2(KEYINPUT54), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n637), .A2(new_n638), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n782), .B1(new_n789), .B2(KEYINPUT55), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n785), .A2(new_n643), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(KEYINPUT54), .A3(new_n650), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT116), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n796), .B(KEYINPUT55), .C1(new_n791), .C2(new_n792), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n671), .B(new_n790), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n240), .B1(new_n239), .B2(new_n245), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n255), .B1(new_n254), .B2(new_n256), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n205), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n670), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n652), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n590), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n590), .A2(new_n790), .A3(new_n803), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n795), .A2(new_n797), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n781), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n796), .B1(new_n789), .B2(KEYINPUT55), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n793), .A2(KEYINPUT116), .A3(new_n794), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(new_n590), .A3(new_n803), .A4(new_n790), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n802), .B1(new_n648), .B2(new_n651), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n651), .B1(new_n793), .B2(new_n794), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n267), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n812), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT117), .B(new_n813), .C1(new_n817), .C2(new_n590), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n809), .A2(new_n673), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n653), .A2(new_n267), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n345), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n547), .A3(new_n549), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(new_n268), .A3(new_n267), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n676), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n679), .A2(new_n680), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n825), .A2(new_n826), .A3(new_n525), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n671), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n823), .B1(new_n828), .B2(new_n268), .ZN(G1340gat));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n277), .A3(new_n652), .ZN(new_n830));
  OAI21_X1  g629(.A(G120gat), .B1(new_n822), .B2(new_n672), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1341gat));
  INV_X1    g631(.A(G127gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n827), .A2(new_n833), .A3(new_n625), .ZN(new_n834));
  OAI21_X1  g633(.A(G127gat), .B1(new_n822), .B2(new_n673), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1342gat));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n825), .A2(new_n826), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n591), .A2(G134gat), .A3(new_n525), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT119), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n837), .A3(new_n839), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n842), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n822), .B2(new_n591), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  NOR3_X1   g645(.A1(new_n739), .A2(new_n345), .A3(new_n525), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n511), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n793), .A2(new_n794), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n671), .A2(new_n790), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n590), .B1(new_n804), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n673), .B1(new_n853), .B2(new_n808), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n850), .B1(new_n854), .B2(new_n820), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT120), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n824), .B2(new_n745), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n671), .B(new_n847), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G141gat), .ZN(new_n859));
  NOR2_X1   g658(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n739), .A2(new_n511), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n267), .A2(G141gat), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n821), .A2(new_n549), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n859), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n861), .B1(new_n859), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(G1344gat));
  AND2_X1   g668(.A1(new_n821), .A2(new_n862), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(new_n291), .A3(new_n549), .A4(new_n652), .ZN(new_n871));
  INV_X1    g670(.A(new_n847), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n855), .B(KEYINPUT120), .Z(new_n873));
  NAND2_X1  g672(.A1(new_n824), .A2(new_n745), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n848), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT59), .B(new_n291), .C1(new_n876), .C2(new_n652), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n850), .B1(new_n819), .B2(new_n820), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n854), .A2(new_n820), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n745), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n652), .B(new_n847), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n871), .B1(new_n877), .B2(new_n883), .ZN(G1345gat));
  NAND2_X1  g683(.A1(new_n870), .A2(new_n549), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n673), .ZN(new_n886));
  AOI21_X1  g685(.A(G155gat), .B1(new_n886), .B2(KEYINPUT122), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n885), .B2(new_n673), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n673), .A2(new_n284), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n887), .A2(new_n889), .B1(new_n876), .B2(new_n890), .ZN(G1346gat));
  NAND4_X1  g690(.A1(new_n870), .A2(new_n285), .A3(new_n549), .A4(new_n590), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n590), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n894), .B2(new_n285), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n676), .A2(new_n549), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n819), .B2(new_n820), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n547), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n899), .A2(new_n349), .A3(new_n267), .ZN(new_n900));
  AOI211_X1 g699(.A(new_n826), .B(new_n897), .C1(new_n819), .C2(new_n820), .ZN(new_n901));
  AOI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n671), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n902), .ZN(G1348gat));
  INV_X1    g702(.A(new_n899), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(G176gat), .A3(new_n652), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT123), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(KEYINPUT123), .ZN(new_n907));
  AOI21_X1  g706(.A(G176gat), .B1(new_n901), .B2(new_n652), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G1349gat));
  OAI21_X1  g708(.A(G183gat), .B1(new_n899), .B2(new_n673), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n901), .A2(new_n378), .A3(new_n625), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n901), .A2(new_n360), .A3(new_n590), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n904), .A2(new_n590), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(G190gat), .ZN(new_n917));
  AOI211_X1 g716(.A(KEYINPUT61), .B(new_n360), .C1(new_n904), .C2(new_n590), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(G1351gat));
  NOR2_X1   g718(.A1(new_n739), .A2(new_n897), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n874), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(KEYINPUT124), .B(G197gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n671), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n879), .A2(new_n881), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n921), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n671), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n930), .B2(new_n923), .ZN(G1352gat));
  NOR4_X1   g730(.A1(new_n874), .A2(G204gat), .A3(new_n672), .A4(new_n921), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n928), .A2(new_n652), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G204gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n934), .A2(new_n935), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n415), .A3(new_n625), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n625), .B(new_n920), .C1(new_n879), .C2(new_n881), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT127), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n940), .B(new_n946), .C1(new_n942), .C2(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1354gat));
  NAND3_X1  g747(.A1(new_n922), .A2(new_n398), .A3(new_n590), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n928), .A2(new_n590), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(new_n398), .ZN(G1355gat));
endmodule


