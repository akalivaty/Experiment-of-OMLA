//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G58), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  INV_X1    g0020(.A(new_n201), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(new_n219), .A2(new_n220), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n227), .B1(new_n220), .B2(new_n219), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n217), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n209), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT64), .Z(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(G97), .B(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n210), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G351));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT8), .A2(G58), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT65), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT8), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n225), .A2(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n224), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(new_n265), .B2(new_n261), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n267), .A2(G50), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n265), .A2(new_n202), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n262), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT68), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n273), .A2(new_n277), .A3(new_n274), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n262), .A2(KEYINPUT9), .A3(new_n271), .A4(new_n272), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT69), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n259), .A2(new_n261), .B1(new_n202), .B2(new_n265), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n283), .A2(KEYINPUT69), .A3(KEYINPUT9), .A4(new_n271), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G77), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n287), .B1(new_n288), .B2(new_n285), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  OAI211_X1 g0093(.A(G1), .B(G13), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G274), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n298), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n294), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n300), .B1(new_n303), .B2(G226), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n282), .A2(new_n284), .B1(new_n306), .B2(G190), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n279), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT70), .B1(new_n305), .B2(G200), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n312), .A2(KEYINPUT10), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n279), .A2(new_n307), .A3(new_n310), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT71), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT10), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n316), .B2(KEYINPUT10), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n305), .A2(new_n321), .B1(new_n271), .B2(new_n283), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G179), .B2(new_n305), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n210), .A2(G20), .ZN(new_n325));
  INV_X1    g0125(.A(new_n248), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n325), .B1(new_n258), .B2(new_n288), .C1(new_n326), .C2(new_n202), .ZN(new_n327));
  XOR2_X1   g0127(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n328));
  AND3_X1   g0128(.A1(new_n327), .A2(new_n261), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n327), .B2(new_n261), .ZN(new_n330));
  INV_X1    g0130(.A(new_n261), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G68), .A3(new_n268), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n265), .A2(KEYINPUT12), .A3(new_n210), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT12), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n264), .B2(G68), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n329), .A2(new_n330), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n292), .A2(KEYINPUT3), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n339), .A2(new_n341), .A3(G232), .A4(G1698), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n285), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n339), .A2(new_n341), .A3(G226), .A4(new_n286), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n344), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT73), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n347), .A2(new_n346), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT73), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n345), .A4(new_n344), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n295), .A3(new_n352), .ZN(new_n353));
  XOR2_X1   g0153(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n354));
  AOI21_X1  g0154(.A(new_n300), .B1(new_n303), .B2(G238), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  INV_X1    g0157(.A(new_n355), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n294), .B1(new_n348), .B2(KEYINPUT73), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n352), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n356), .B(G179), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT76), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n361), .B(new_n362), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n365));
  OAI21_X1  g0165(.A(G169), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(G169), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n338), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n257), .A2(new_n265), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(new_n257), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n252), .A2(new_n254), .A3(G68), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n225), .B1(new_n376), .B2(new_n221), .ZN(new_n377));
  INV_X1    g0177(.A(G159), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n326), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT77), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n339), .A2(new_n341), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n381), .B2(new_n225), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n383), .B(G20), .C1(new_n339), .C2(new_n341), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT77), .ZN(new_n386));
  INV_X1    g0186(.A(new_n379), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT65), .B(G58), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n201), .B1(new_n388), .B2(G68), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n386), .B(new_n387), .C1(new_n389), .C2(new_n225), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n380), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT16), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n380), .A2(new_n385), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n380), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n380), .A2(new_n385), .A3(new_n390), .A4(new_n395), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n398), .A2(new_n261), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n375), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n299), .B1(new_n302), .B2(new_n209), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  XOR2_X1   g0202(.A(new_n402), .B(KEYINPUT79), .Z(new_n403));
  NAND3_X1  g0203(.A1(new_n285), .A2(G223), .A3(new_n286), .ZN(new_n404));
  INV_X1    g0204(.A(G226), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n403), .B(new_n404), .C1(new_n405), .C2(new_n289), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n401), .B1(new_n406), .B2(new_n295), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n407), .A2(G179), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n321), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n372), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n397), .A2(new_n399), .ZN(new_n412));
  INV_X1    g0212(.A(new_n375), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n410), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT18), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n407), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(G190), .B2(new_n407), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT17), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n400), .A2(new_n422), .A3(new_n419), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n411), .A2(new_n416), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g0224(.A(KEYINPUT8), .B(G58), .Z(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n258), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n261), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT67), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n331), .A2(G77), .A3(new_n268), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n288), .B2(new_n265), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G107), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n289), .A2(new_n211), .B1(new_n434), .B2(new_n285), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n381), .A2(new_n209), .A3(G1698), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n295), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n300), .B1(new_n303), .B2(G244), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G179), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n321), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n433), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n440), .A2(new_n417), .ZN(new_n446));
  INV_X1    g0246(.A(G190), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n433), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(G200), .B1(new_n364), .B2(new_n365), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n356), .B(G190), .C1(new_n357), .C2(new_n360), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n337), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n371), .A2(new_n424), .A3(new_n450), .A4(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n324), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n263), .B(G45), .C1(new_n293), .C2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(G274), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G41), .ZN(new_n459));
  OR3_X1    g0259(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n294), .B(G270), .C1(new_n456), .C2(new_n459), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n339), .A2(new_n341), .A3(G264), .A4(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT82), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n285), .A2(new_n465), .A3(G264), .A4(G1698), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n381), .A2(G303), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n285), .A2(G257), .A3(new_n286), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n464), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n462), .B1(new_n469), .B2(new_n295), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT80), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n263), .B2(G33), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n292), .A2(KEYINPUT80), .A3(G1), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n266), .A2(new_n474), .A3(G116), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n263), .A2(new_n476), .A3(G13), .A4(G20), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT83), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n260), .A2(new_n224), .B1(G20), .B2(new_n476), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n225), .C1(G33), .C2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT20), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n475), .B(new_n478), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n470), .A2(G179), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n470), .A2(KEYINPUT84), .A3(new_n485), .A4(G179), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n339), .A2(new_n341), .A3(G257), .A4(G1698), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT86), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n285), .A2(KEYINPUT86), .A3(G257), .A4(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G294), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n285), .A2(G250), .A3(new_n286), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n295), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n456), .A2(new_n459), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(KEYINPUT87), .A3(G264), .A4(new_n294), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n294), .B(G264), .C1(new_n456), .C2(new_n459), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(new_n460), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n321), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n266), .A2(new_n474), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n264), .A2(G107), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n509), .A2(KEYINPUT25), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(KEYINPUT25), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n508), .A2(G107), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n225), .B2(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n434), .A2(KEYINPUT23), .A3(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n292), .A2(new_n476), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n225), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n339), .A2(new_n341), .A3(new_n225), .A4(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT22), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n285), .A2(new_n522), .A3(new_n225), .A4(G87), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n519), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n261), .B1(new_n524), .B2(KEYINPUT24), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(new_n523), .ZN(new_n526));
  INV_X1    g0326(.A(new_n519), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n526), .A2(KEYINPUT24), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n512), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n295), .A2(new_n497), .B1(new_n500), .B2(new_n503), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n441), .A3(new_n460), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n506), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n470), .ZN(new_n533));
  NOR2_X1   g0333(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n533), .A2(G169), .A3(new_n485), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n485), .A2(G169), .ZN(new_n537));
  AND2_X1   g0337(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n537), .A2(new_n470), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n490), .A2(new_n532), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n505), .A2(G200), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n530), .A2(G190), .A3(new_n460), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n526), .A2(new_n527), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n524), .A2(KEYINPUT24), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n261), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n541), .A2(new_n542), .A3(new_n547), .A4(new_n512), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(new_n286), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT4), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n480), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n295), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n294), .B(G257), .C1(new_n456), .C2(new_n459), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n460), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n321), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n248), .A2(G77), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n434), .A2(G97), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT6), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n563), .B2(new_n240), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n561), .B1(new_n565), .B2(new_n225), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n383), .B1(new_n285), .B2(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n381), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n434), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n261), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n264), .A2(G97), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n507), .B2(new_n481), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n557), .B1(new_n554), .B2(new_n295), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n441), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n560), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n559), .A2(G200), .ZN(new_n579));
  OAI21_X1  g0379(.A(G107), .B1(new_n382), .B2(new_n384), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n481), .A2(G107), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n562), .A2(new_n581), .A3(new_n563), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n563), .B2(new_n562), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G20), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n584), .A3(new_n561), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n573), .B1(new_n585), .B2(new_n261), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n576), .A2(G190), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n579), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n548), .A2(new_n578), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n225), .B1(new_n346), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(G87), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n481), .A3(new_n434), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n339), .A2(new_n341), .A3(new_n225), .A4(G68), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n590), .B1(new_n258), .B2(new_n481), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n261), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n427), .A2(new_n265), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(new_n427), .C2(new_n507), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n339), .A2(new_n341), .A3(G238), .A4(new_n286), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(G1698), .ZN(new_n602));
  INV_X1    g0402(.A(new_n517), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n295), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT81), .B1(new_n297), .B2(G1), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT81), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n263), .A3(G45), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(G33), .A2(G41), .ZN(new_n610));
  OAI21_X1  g0410(.A(G250), .B1(new_n610), .B2(new_n224), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n263), .A2(G45), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n609), .A2(new_n611), .B1(new_n457), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(new_n614), .A3(new_n441), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n295), .B2(new_n604), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n600), .B(new_n615), .C1(G169), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n605), .A2(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G200), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(G190), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n597), .A2(new_n261), .B1(new_n265), .B2(new_n427), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n266), .A2(new_n474), .A3(G87), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n485), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n533), .B2(new_n447), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n470), .A2(new_n417), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n617), .B(new_n623), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n540), .A2(new_n589), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n455), .A2(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n323), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n416), .A2(new_n411), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n361), .A2(KEYINPUT76), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n361), .A2(KEYINPUT76), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n367), .B(new_n369), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n338), .B1(new_n453), .B2(new_n445), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n421), .A2(new_n423), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n631), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n320), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n638), .B2(new_n639), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n630), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n455), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT91), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n623), .A2(new_n617), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT26), .B1(new_n646), .B2(new_n578), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n617), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n616), .B2(new_n417), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n618), .A2(KEYINPUT88), .A3(G200), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n620), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n621), .A2(new_n622), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT89), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT89), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n621), .A2(new_n655), .A3(new_n622), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n617), .B1(new_n652), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n578), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n645), .B1(new_n648), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n617), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n654), .A2(new_n656), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n650), .A2(new_n651), .A3(new_n620), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(new_n578), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(KEYINPUT91), .A3(new_n617), .A4(new_n647), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n536), .A2(new_n539), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n490), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT90), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT90), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(new_n672), .A3(new_n490), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n532), .A3(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n588), .A2(new_n578), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(new_n664), .A3(new_n548), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n660), .A2(new_n668), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n643), .B1(new_n644), .B2(new_n678), .ZN(G369));
  NOR2_X1   g0479(.A1(new_n625), .A2(new_n626), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n225), .A2(G13), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n263), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n624), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n670), .A2(new_n680), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n671), .A2(new_n673), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT93), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n529), .A2(new_n687), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n548), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n532), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n532), .A2(new_n687), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n687), .B1(new_n669), .B2(new_n490), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n702), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n704), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n218), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n593), .A2(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n222), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT26), .B1(new_n658), .B2(new_n578), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n646), .A2(new_n578), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n661), .B1(new_n718), .B2(new_n665), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n490), .A2(new_n532), .A3(new_n536), .A4(new_n539), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n717), .B(new_n719), .C1(new_n676), .C2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT95), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n721), .A2(new_n722), .A3(new_n688), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n721), .B2(new_n688), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT29), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n678), .B2(new_n687), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n548), .A2(new_n578), .A3(new_n588), .ZN(new_n729));
  INV_X1    g0529(.A(new_n627), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n720), .A2(new_n729), .A3(new_n730), .A4(new_n688), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT31), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n616), .A2(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n533), .A2(new_n505), .A3(new_n559), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT94), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n734), .B(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n530), .A2(new_n576), .A3(new_n616), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n470), .A2(G179), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n470), .A2(G179), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n498), .A2(new_n504), .A3(new_n616), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT30), .A4(new_n576), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n687), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n732), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n748), .B(new_n688), .C1(new_n744), .C2(new_n734), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n697), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n728), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n716), .B1(new_n754), .B2(G1), .ZN(G364));
  INV_X1    g0555(.A(new_n696), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n263), .B1(new_n681), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n711), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n696), .A2(new_n697), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n710), .A2(new_n381), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n764), .A2(G355), .B1(new_n476), .B2(new_n710), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n246), .A2(new_n297), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n710), .A2(new_n285), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G45), .B2(new_n222), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n765), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n224), .B1(G20), .B2(new_n321), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n761), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT96), .Z(new_n776));
  NOR2_X1   g0576(.A1(new_n225), .A2(new_n447), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n441), .A3(G200), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT100), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT100), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n225), .A2(G190), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n441), .A3(new_n417), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G303), .A2(new_n782), .B1(new_n788), .B2(G329), .ZN(new_n789));
  INV_X1    g0589(.A(new_n783), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n790), .A2(G179), .A3(new_n417), .ZN(new_n791));
  NOR4_X1   g0591(.A1(new_n225), .A2(new_n441), .A3(new_n447), .A4(G200), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n791), .A2(G283), .B1(G322), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n790), .A2(new_n441), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n381), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n447), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n225), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n797), .B1(G294), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n441), .A2(new_n417), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n777), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n783), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G326), .A2(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n789), .A2(new_n793), .A3(new_n801), .A4(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n803), .A2(new_n202), .B1(new_n805), .B2(new_n210), .ZN(new_n810));
  INV_X1    g0610(.A(new_n791), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n285), .B1(new_n481), .B2(new_n799), .C1(new_n811), .C2(new_n434), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n810), .B(new_n812), .C1(G77), .C2(new_n794), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n782), .A2(G87), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n792), .B(KEYINPUT97), .Z(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n813), .B(new_n814), .C1(new_n255), .C2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT99), .B(G159), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n788), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT32), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n809), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n776), .B1(new_n821), .B2(new_n773), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n772), .B(KEYINPUT101), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n756), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n763), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n660), .A2(new_n668), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n674), .A2(new_n677), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n687), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n444), .A2(new_n687), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n688), .B1(new_n430), .B2(new_n432), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n449), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(new_n444), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n830), .B(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(new_n752), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT104), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(KEYINPUT104), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n835), .A2(new_n752), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n837), .A2(new_n761), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n773), .A2(new_n770), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n761), .B1(new_n288), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n773), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n794), .A2(new_n818), .B1(new_n804), .B2(G137), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  INV_X1    g0645(.A(G143), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n844), .B1(new_n845), .B2(new_n805), .C1(new_n816), .C2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT34), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n787), .A2(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n285), .B1(new_n255), .B2(new_n799), .C1(new_n811), .C2(new_n210), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n850), .B(new_n851), .C1(G50), .C2(new_n782), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n781), .A2(new_n434), .B1(new_n787), .B2(new_n796), .ZN(new_n853));
  INV_X1    g0653(.A(G303), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n381), .B1(new_n803), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n795), .A2(new_n476), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n791), .A2(G87), .ZN(new_n857));
  INV_X1    g0657(.A(G283), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n805), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n853), .A2(new_n855), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n800), .A2(G97), .B1(G294), .B2(new_n792), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT103), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n848), .A2(new_n852), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n842), .B1(new_n843), .B2(new_n863), .C1(new_n834), .C2(new_n771), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n840), .A2(new_n864), .ZN(G384));
  OAI211_X1 g0665(.A(G116), .B(new_n226), .C1(new_n583), .C2(KEYINPUT35), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(KEYINPUT35), .B2(new_n583), .ZN(new_n867));
  XOR2_X1   g0667(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n223), .A2(G77), .A3(new_n376), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n263), .B(G13), .C1(new_n870), .C2(new_n242), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n831), .B1(new_n830), .B2(new_n834), .ZN(new_n873));
  INV_X1    g0673(.A(new_n453), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n634), .B2(new_n338), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n688), .A2(new_n337), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n367), .A2(new_n369), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n361), .B(KEYINPUT76), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n337), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n875), .A2(new_n877), .B1(new_n880), .B2(new_n687), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n392), .A2(new_n394), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n375), .B1(new_n884), .B2(new_n261), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n685), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n424), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n412), .A2(new_n413), .A3(new_n419), .ZN(new_n889));
  INV_X1    g0689(.A(new_n685), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n408), .A2(new_n409), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n420), .B(new_n894), .C1(new_n400), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n883), .B1(new_n888), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT38), .B(new_n896), .C1(new_n424), .C2(new_n887), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n882), .A2(new_n900), .B1(new_n631), .B2(new_n890), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n371), .A2(new_n687), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(KEYINPUT107), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n631), .A2(new_n636), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n886), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT107), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT38), .A4(new_n896), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n400), .A2(new_n891), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n889), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n895), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n414), .A2(new_n890), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n631), .B2(new_n636), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT106), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n424), .A2(KEYINPUT106), .A3(new_n913), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n883), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n909), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n898), .A2(new_n899), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT39), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n903), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n901), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n725), .A2(new_n455), .A3(new_n727), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT108), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT108), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n725), .A2(new_n455), .A3(new_n727), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n643), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n924), .B(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n909), .A2(new_n918), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n688), .B1(new_n736), .B2(new_n744), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n731), .B2(KEYINPUT31), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n746), .A2(new_n748), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n833), .A2(new_n444), .ZN(new_n938));
  INV_X1    g0738(.A(new_n831), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n881), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n932), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n934), .A2(KEYINPUT31), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n748), .B1(new_n628), .B2(new_n688), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n934), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n874), .B(new_n876), .C1(new_n634), .C2(new_n338), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n634), .A2(new_n338), .A3(new_n687), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n945), .B(new_n834), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(G330), .B1(new_n942), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n697), .B1(new_n747), .B2(new_n943), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n455), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n941), .A2(new_n932), .A3(new_n921), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n949), .B1(new_n909), .B2(new_n918), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n956), .B2(new_n932), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(new_n455), .A3(new_n945), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n931), .A2(new_n959), .B1(new_n263), .B2(new_n681), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n960), .A2(KEYINPUT109), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n931), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n960), .B2(KEYINPUT109), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n872), .B1(new_n961), .B2(new_n963), .ZN(G367));
  OAI211_X1 g0764(.A(new_n588), .B(new_n578), .C1(new_n586), .C2(new_n688), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n666), .A2(new_n687), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n708), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT44), .ZN(new_n970));
  INV_X1    g0770(.A(new_n968), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n971), .A2(new_n706), .A3(new_n707), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n704), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(KEYINPUT113), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT113), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n704), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n977), .A3(new_n704), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n703), .A2(new_n705), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n706), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n757), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n698), .B1(new_n706), .B2(new_n982), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n753), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n711), .B(KEYINPUT41), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n758), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n704), .A2(new_n971), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n662), .A2(new_n688), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n661), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n658), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT112), .Z(new_n996));
  XNOR2_X1  g0796(.A(new_n991), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n706), .A2(new_n968), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT111), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n578), .B1(new_n966), .B2(new_n532), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n688), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n998), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n997), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n990), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n767), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n237), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n774), .B1(new_n218), .B2(new_n427), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n760), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(G294), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n795), .A2(new_n858), .B1(new_n1015), .B2(new_n805), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n811), .A2(new_n481), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n381), .B1(new_n803), .B2(new_n796), .C1(new_n799), .C2(new_n434), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(G317), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n787), .C1(new_n854), .C2(new_n816), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT114), .B1(new_n781), .B2(new_n476), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1022), .A2(KEYINPUT46), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT46), .B2(new_n1022), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n811), .A2(new_n288), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n806), .B2(new_n818), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n792), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1027), .B1(new_n846), .B2(new_n803), .C1(new_n845), .C2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n285), .B1(new_n210), .B2(new_n799), .C1(new_n795), .C2(new_n202), .ZN(new_n1030));
  INV_X1    g0830(.A(G137), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n781), .A2(new_n255), .B1(new_n787), .B2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1025), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(new_n843), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1034), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1014), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n994), .A2(new_n823), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1010), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT116), .ZN(G387));
  AND3_X1   g0842(.A1(new_n986), .A2(KEYINPUT117), .A3(new_n759), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT117), .B1(new_n986), .B2(new_n759), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n984), .A2(new_n985), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n753), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n986), .A2(new_n754), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n711), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n794), .A2(G68), .B1(new_n804), .B2(G159), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n202), .B2(new_n1028), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n799), .A2(new_n427), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1051), .A2(new_n381), .A3(new_n1017), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n257), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n806), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n788), .A2(G150), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n782), .A2(G77), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n788), .A2(G326), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n285), .B1(new_n791), .B2(G116), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n794), .A2(G303), .B1(new_n804), .B2(G322), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n796), .B2(new_n805), .C1(new_n816), .C2(new_n1020), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT48), .Z(new_n1063));
  OAI22_X1  g0863(.A1(new_n781), .A2(new_n1015), .B1(new_n858), .B2(new_n799), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1059), .B(new_n1060), .C1(new_n1065), .C2(KEYINPUT49), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(KEYINPUT49), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1058), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT118), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n843), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1011), .B1(new_n233), .B2(G45), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n713), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n764), .ZN(new_n1074));
  AOI21_X1  g0874(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n425), .A2(new_n202), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n713), .B(new_n1075), .C1(new_n1076), .C2(KEYINPUT50), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(KEYINPUT50), .B2(new_n1076), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1074), .A2(new_n1078), .B1(G107), .B2(new_n218), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n761), .B1(new_n1079), .B2(new_n774), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1071), .B(new_n1080), .C1(new_n703), .C2(new_n823), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1045), .A2(new_n1049), .A3(new_n1081), .ZN(G393));
  INV_X1    g0882(.A(new_n1048), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n981), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n979), .A2(new_n1048), .A3(new_n980), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n711), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n971), .A2(new_n772), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n241), .A2(new_n1011), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n774), .B1(new_n481), .B2(new_n218), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n760), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n795), .A2(new_n1015), .B1(new_n854), .B2(new_n805), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n285), .B(new_n1091), .C1(G107), .C2(new_n791), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G283), .A2(new_n782), .B1(new_n788), .B2(G322), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n476), .C2(new_n799), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n804), .A2(G317), .B1(new_n792), .B2(G311), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1028), .A2(new_n378), .B1(new_n803), .B2(new_n845), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n210), .B2(new_n781), .C1(new_n846), .C2(new_n787), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n794), .A2(new_n425), .B1(new_n806), .B2(G50), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n799), .A2(new_n288), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1100), .A2(new_n285), .A3(new_n857), .A4(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1094), .A2(new_n1096), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1090), .B1(new_n1104), .B2(new_n773), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n981), .A2(new_n759), .B1(new_n1087), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1086), .A2(new_n1106), .ZN(G390));
  OAI21_X1  g0907(.A(new_n903), .B1(new_n873), .B2(new_n881), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n920), .A3(new_n922), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n371), .A2(new_n453), .A3(new_n877), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n947), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n751), .A2(new_n1111), .A3(new_n834), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n902), .B1(new_n909), .B2(new_n918), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n676), .A2(new_n720), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n719), .A2(new_n717), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n688), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT95), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n721), .A2(new_n722), .A3(new_n688), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1118), .A3(new_n939), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n938), .A3(new_n1111), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1113), .A2(KEYINPUT119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT119), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1109), .B(new_n1112), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1108), .A2(new_n920), .A3(new_n922), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1113), .A2(new_n1120), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1113), .A2(KEYINPUT119), .A3(new_n1120), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n940), .B1(new_n1110), .B2(new_n947), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n952), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1123), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(new_n758), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n920), .A2(new_n770), .A3(new_n922), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n841), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n760), .B1(new_n1135), .B2(new_n1054), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n795), .A2(new_n481), .B1(new_n434), .B2(new_n805), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1028), .A2(new_n476), .B1(new_n803), .B2(new_n858), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n285), .B(new_n1101), .C1(G68), .C2(new_n791), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n788), .A2(G294), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1139), .A2(new_n814), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n782), .A2(G150), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n788), .A2(G125), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n285), .B1(new_n1028), .B2(new_n849), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G159), .B2(new_n800), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  AOI22_X1  g0948(.A1(new_n794), .A2(new_n1148), .B1(new_n806), .B2(G137), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n791), .A2(G50), .B1(new_n804), .B2(G128), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1145), .A2(new_n1147), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1142), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1136), .B1(new_n1152), .B2(new_n773), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1134), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1133), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1119), .A2(new_n938), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1112), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1111), .B1(new_n952), .B2(new_n834), .ZN(new_n1158));
  OAI211_X1 g0958(.A(G330), .B(new_n834), .C1(new_n935), .C2(new_n749), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1130), .A2(new_n952), .B1(new_n881), .B2(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1157), .A2(new_n1158), .B1(new_n1160), .B2(new_n873), .ZN(new_n1161));
  AND4_X1   g0961(.A1(new_n643), .A2(new_n1161), .A3(new_n929), .A4(new_n953), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(new_n1123), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n711), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n929), .A3(new_n643), .A4(new_n953), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1164), .A2(KEYINPUT120), .B1(new_n1132), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT120), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1163), .A2(new_n1167), .A3(new_n711), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1155), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(G378));
  NAND3_X1  g0970(.A1(new_n929), .A2(new_n643), .A3(new_n953), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1163), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n324), .A2(new_n273), .A3(new_n890), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n273), .A2(new_n890), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n320), .A2(new_n323), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1174), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n957), .A2(G330), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n957), .B2(G330), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n924), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1182), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n951), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n901), .A2(new_n923), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n957), .A2(G330), .A3(new_n1182), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1185), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1173), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT123), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1163), .A2(new_n1172), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1196));
  OAI21_X1  g0996(.A(KEYINPUT123), .B1(new_n1196), .B2(KEYINPUT57), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n712), .B1(new_n1196), .B2(KEYINPUT57), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1186), .A2(new_n770), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n760), .B1(new_n1135), .B2(G50), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n794), .A2(G137), .B1(new_n806), .B2(G132), .ZN(new_n1202));
  INV_X1    g1002(.A(G128), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n1203), .B2(new_n1028), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n800), .A2(G150), .B1(new_n804), .B2(G125), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT122), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n782), .C2(new_n1148), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT59), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n788), .A2(G124), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n791), .C2(new_n818), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n285), .A2(G41), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G50), .B(new_n1214), .C1(new_n292), .C2(new_n293), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n811), .A2(new_n255), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n795), .A2(new_n427), .B1(new_n481), .B2(new_n805), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G116), .C2(new_n804), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1214), .B1(new_n1028), .B2(new_n434), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G68), .B2(new_n800), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n788), .A2(G283), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1057), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1223));
  AOI21_X1  g1023(.A(new_n1215), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1213), .B(new_n1224), .C1(new_n1223), .C2(new_n1222), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1201), .B1(new_n1225), .B2(new_n773), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1191), .A2(new_n759), .B1(new_n1200), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1199), .A2(new_n1227), .ZN(G375));
  INV_X1    g1028(.A(new_n1161), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1171), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n988), .A3(new_n1165), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1161), .A2(new_n759), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1111), .A2(new_n771), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n760), .B1(new_n1135), .B2(G68), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1026), .A2(new_n285), .A3(new_n1052), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G116), .A2(new_n806), .B1(new_n792), .B2(G283), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n1015), .B2(new_n803), .C1(new_n434), .C2(new_n795), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n781), .A2(new_n481), .B1(new_n787), .B2(new_n854), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT125), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G132), .A2(new_n804), .B1(new_n806), .B2(new_n1148), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n845), .B2(new_n795), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n799), .A2(new_n202), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1245), .A2(new_n381), .A3(new_n1216), .A4(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G159), .A2(new_n782), .B1(new_n815), .B2(G137), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n1203), .C2(new_n787), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(KEYINPUT125), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1243), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1236), .B1(new_n1251), .B2(new_n773), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1234), .A2(new_n1235), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1232), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1231), .A2(new_n1255), .ZN(G381));
  NAND3_X1  g1056(.A1(new_n1199), .A2(new_n1169), .A3(new_n1227), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1045), .A2(new_n826), .A3(new_n1049), .A4(new_n1081), .ZN(new_n1258));
  OR4_X1    g1058(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1258), .ZN(new_n1259));
  OR3_X1    g1059(.A1(G387), .A2(new_n1257), .A3(new_n1259), .ZN(G407));
  OAI211_X1 g1060(.A(G407), .B(G213), .C1(G343), .C2(new_n1257), .ZN(G409));
  INV_X1    g1061(.A(new_n1049), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1081), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1263));
  OAI21_X1  g1063(.A(G396), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1258), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G390), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT116), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1264), .B2(new_n1258), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(G390), .B2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1010), .A2(new_n1040), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1041), .B(new_n1266), .C1(G390), .C2(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1165), .A2(KEYINPUT60), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n712), .B1(new_n1274), .B2(new_n1230), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1171), .A2(new_n1229), .A3(KEYINPUT60), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1275), .A2(KEYINPUT126), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT126), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1255), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G384), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1274), .A2(new_n1230), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n711), .A3(new_n1276), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1275), .A2(KEYINPUT126), .A3(new_n1276), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G384), .A3(new_n1255), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n686), .A2(G213), .A3(G2897), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1281), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1289), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G384), .B1(new_n1287), .B2(new_n1255), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n1280), .B(new_n1254), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1169), .B1(new_n1199), .B2(new_n1227), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1164), .A2(KEYINPUT120), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1132), .A2(new_n1165), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1168), .A3(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1133), .A2(new_n1154), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1196), .A2(new_n988), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1227), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n686), .A2(G213), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1290), .B(new_n1294), .C1(new_n1295), .C2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1281), .A2(new_n1288), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1295), .A2(new_n1303), .A3(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1304), .B(new_n1305), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G375), .A2(G378), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1303), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1306), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(KEYINPUT62), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1273), .B1(new_n1309), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1273), .B1(KEYINPUT63), .B2(new_n1307), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1313), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1315), .A2(new_n1320), .ZN(G405));
  NAND2_X1  g1121(.A1(new_n1310), .A2(new_n1257), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1306), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1310), .A2(new_n1257), .A3(new_n1312), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1271), .A2(new_n1272), .A3(KEYINPUT127), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT127), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1327), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1329), .A2(new_n1323), .A3(new_n1324), .A4(new_n1325), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(G402));
endmodule


