

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U555 ( .A1(n527), .A2(n524), .ZN(n769) );
  XNOR2_X1 U556 ( .A(n748), .B(KEYINPUT104), .ZN(n753) );
  NAND2_X1 U557 ( .A1(n625), .A2(n624), .ZN(n1016) );
  INV_X1 U558 ( .A(G2104), .ZN(n584) );
  NAND2_X1 U559 ( .A1(n546), .A2(KEYINPUT40), .ZN(n544) );
  INV_X1 U560 ( .A(G2105), .ZN(n558) );
  NOR2_X1 U561 ( .A1(n853), .A2(n852), .ZN(n547) );
  NOR2_X1 U562 ( .A1(n735), .A2(n1016), .ZN(n736) );
  NOR2_X1 U563 ( .A1(n620), .A2(n619), .ZN(n622) );
  INV_X1 U564 ( .A(KEYINPUT75), .ZN(n621) );
  AND2_X1 U565 ( .A1(n558), .A2(G2104), .ZN(n929) );
  NAND2_X1 U566 ( .A1(n558), .A2(n584), .ZN(n583) );
  NOR2_X1 U567 ( .A1(n548), .A2(n544), .ZN(n543) );
  NAND2_X1 U568 ( .A1(n862), .A2(n545), .ZN(n539) );
  INV_X1 U569 ( .A(n544), .ZN(n541) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n933) );
  XNOR2_X1 U571 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U572 ( .A1(n551), .A2(n558), .ZN(n550) );
  NOR2_X1 U573 ( .A1(n553), .A2(n552), .ZN(n551) );
  INV_X1 U574 ( .A(G101), .ZN(n552) );
  AND2_X1 U575 ( .A1(n557), .A2(n555), .ZN(n554) );
  NAND2_X1 U576 ( .A1(G2105), .A2(KEYINPUT23), .ZN(n557) );
  NAND2_X1 U577 ( .A1(n556), .A2(KEYINPUT23), .ZN(n555) );
  NAND2_X1 U578 ( .A1(G101), .A2(G2104), .ZN(n556) );
  XNOR2_X1 U579 ( .A(n534), .B(n522), .ZN(n533) );
  AND2_X1 U580 ( .A1(n791), .A2(n790), .ZN(n792) );
  INV_X1 U581 ( .A(KEYINPUT23), .ZN(n549) );
  INV_X1 U582 ( .A(KEYINPUT0), .ZN(n560) );
  XNOR2_X1 U583 ( .A(n622), .B(n621), .ZN(n625) );
  NOR2_X1 U584 ( .A1(n543), .A2(n538), .ZN(n537) );
  NOR2_X1 U585 ( .A1(n592), .A2(n591), .ZN(G164) );
  NOR2_X1 U586 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U587 ( .A1(G164), .A2(G1384), .ZN(n830) );
  XOR2_X1 U588 ( .A(KEYINPUT65), .B(KEYINPUT26), .Z(n522) );
  OR2_X1 U589 ( .A1(G301), .A2(n765), .ZN(n523) );
  XOR2_X1 U590 ( .A(n768), .B(KEYINPUT31), .Z(n524) );
  XNOR2_X1 U591 ( .A(n583), .B(KEYINPUT17), .ZN(n601) );
  AND2_X1 U592 ( .A1(n554), .A2(n550), .ZN(n525) );
  AND2_X1 U593 ( .A1(n830), .A2(n531), .ZN(n526) );
  INV_X1 U594 ( .A(n862), .ZN(n546) );
  INV_X1 U595 ( .A(KEYINPUT40), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n528), .A2(n523), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n528) );
  INV_X1 U598 ( .A(KEYINPUT29), .ZN(n529) );
  NAND2_X1 U599 ( .A1(n757), .A2(n756), .ZN(n530) );
  NAND2_X1 U600 ( .A1(n734), .A2(n830), .ZN(n771) );
  NAND2_X1 U601 ( .A1(n526), .A2(n734), .ZN(n534) );
  INV_X1 U602 ( .A(n981), .ZN(n531) );
  NAND2_X1 U603 ( .A1(n533), .A2(n532), .ZN(n735) );
  NAND2_X1 U604 ( .A1(n771), .A2(G1341), .ZN(n532) );
  NAND2_X1 U605 ( .A1(n537), .A2(n535), .ZN(G329) );
  NAND2_X1 U606 ( .A1(n548), .A2(n536), .ZN(n535) );
  AND2_X1 U607 ( .A1(n547), .A2(n545), .ZN(n536) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n538) );
  NAND2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n540) );
  INV_X1 U610 ( .A(n547), .ZN(n542) );
  OR2_X2 U611 ( .A1(n801), .A2(n800), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(G2104), .ZN(n553) );
  NOR2_X2 U613 ( .A1(n738), .A2(n829), .ZN(n759) );
  BUF_X1 U614 ( .A(n737), .Z(n829) );
  XNOR2_X2 U615 ( .A(n609), .B(KEYINPUT67), .ZN(G160) );
  XOR2_X1 U616 ( .A(KEYINPUT15), .B(n636), .Z(n559) );
  INV_X1 U617 ( .A(KEYINPUT77), .ZN(n627) );
  XNOR2_X1 U618 ( .A(KEYINPUT78), .B(n631), .ZN(n635) );
  NOR2_X1 U619 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U620 ( .A1(n690), .A2(G56), .ZN(n613) );
  NOR2_X1 U621 ( .A1(n687), .A2(G651), .ZN(n626) );
  INV_X1 U622 ( .A(KEYINPUT97), .ZN(n585) );
  INV_X1 U623 ( .A(KEYINPUT68), .ZN(n604) );
  INV_X1 U624 ( .A(KEYINPUT1), .ZN(n561) );
  BUF_X1 U625 ( .A(n626), .Z(n692) );
  NAND2_X1 U626 ( .A1(n608), .A2(n525), .ZN(n609) );
  XNOR2_X2 U627 ( .A(n560), .B(G543), .ZN(n687) );
  NAND2_X1 U628 ( .A1(G51), .A2(n692), .ZN(n564) );
  INV_X1 U629 ( .A(G651), .ZN(n566) );
  NOR2_X1 U630 ( .A1(G543), .A2(n566), .ZN(n562) );
  XNOR2_X2 U631 ( .A(n562), .B(n561), .ZN(n690) );
  NAND2_X1 U632 ( .A1(G63), .A2(n690), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U634 ( .A(KEYINPUT6), .B(n565), .Z(n574) );
  NOR2_X2 U635 ( .A1(n687), .A2(n566), .ZN(n696) );
  NAND2_X1 U636 ( .A1(n696), .A2(G76), .ZN(n567) );
  XNOR2_X1 U637 ( .A(KEYINPUT81), .B(n567), .ZN(n570) );
  NOR2_X4 U638 ( .A1(G543), .A2(G651), .ZN(n693) );
  NAND2_X1 U639 ( .A1(n693), .A2(G89), .ZN(n568) );
  XOR2_X1 U640 ( .A(n568), .B(KEYINPUT4), .Z(n569) );
  NOR2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U642 ( .A(KEYINPUT82), .B(n571), .Z(n572) );
  XNOR2_X1 U643 ( .A(KEYINPUT5), .B(n572), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U645 ( .A(KEYINPUT7), .B(n575), .ZN(G168) );
  XOR2_X1 U646 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U647 ( .A1(G88), .A2(n693), .ZN(n577) );
  NAND2_X1 U648 ( .A1(G75), .A2(n696), .ZN(n576) );
  NAND2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U650 ( .A1(G50), .A2(n692), .ZN(n579) );
  NAND2_X1 U651 ( .A1(G62), .A2(n690), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT90), .ZN(G166) );
  INV_X1 U655 ( .A(G166), .ZN(G303) );
  INV_X1 U656 ( .A(G96), .ZN(G221) );
  INV_X1 U657 ( .A(G120), .ZN(G236) );
  NAND2_X1 U658 ( .A1(n601), .A2(G138), .ZN(n588) );
  AND2_X4 U659 ( .A1(n584), .A2(G2105), .ZN(n657) );
  NAND2_X1 U660 ( .A1(G126), .A2(n657), .ZN(n586) );
  XNOR2_X1 U661 ( .A(n586), .B(n585), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G102), .A2(n929), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G114), .A2(n933), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U666 ( .A1(G52), .A2(n692), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G64), .A2(n690), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G90), .A2(n693), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G77), .A2(n696), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT70), .B(n597), .Z(n598) );
  XNOR2_X1 U673 ( .A(KEYINPUT9), .B(n598), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G171) );
  NAND2_X1 U675 ( .A1(G137), .A2(n601), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G113), .A2(n933), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U678 ( .A1(G125), .A2(n657), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G94), .A2(G452), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n610), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U681 ( .A1(G7), .A2(G661), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U683 ( .A(G223), .ZN(n872) );
  NAND2_X1 U684 ( .A1(n872), .A2(G567), .ZN(n612) );
  XOR2_X1 U685 ( .A(KEYINPUT11), .B(n612), .Z(G234) );
  XOR2_X1 U686 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(n620) );
  NAND2_X1 U688 ( .A1(G68), .A2(n696), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n693), .A2(G81), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n615), .B(KEYINPUT12), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U692 ( .A(KEYINPUT13), .B(n618), .Z(n619) );
  NAND2_X1 U693 ( .A1(n692), .A2(G43), .ZN(n623) );
  XNOR2_X1 U694 ( .A(KEYINPUT76), .B(n623), .ZN(n624) );
  INV_X1 U695 ( .A(G860), .ZN(n649) );
  OR2_X1 U696 ( .A1(n1016), .A2(n649), .ZN(G153) );
  INV_X1 U697 ( .A(G171), .ZN(G301) );
  NAND2_X1 U698 ( .A1(n626), .A2(G54), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n696), .A2(G79), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U702 ( .A1(G66), .A2(n690), .ZN(n633) );
  NAND2_X1 U703 ( .A1(G92), .A2(n693), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X2 U705 ( .A(KEYINPUT79), .B(n559), .Z(n1012) );
  OR2_X1 U706 ( .A1(n1012), .A2(G868), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT80), .ZN(n639) );
  NAND2_X1 U708 ( .A1(G868), .A2(G301), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n639), .A2(n638), .ZN(G284) );
  NAND2_X1 U710 ( .A1(G53), .A2(n692), .ZN(n641) );
  NAND2_X1 U711 ( .A1(G65), .A2(n690), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U713 ( .A(KEYINPUT72), .B(n642), .ZN(n646) );
  NAND2_X1 U714 ( .A1(G91), .A2(n693), .ZN(n644) );
  NAND2_X1 U715 ( .A1(G78), .A2(n696), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n1002) );
  XNOR2_X1 U718 ( .A(n1002), .B(KEYINPUT73), .ZN(G299) );
  NAND2_X1 U719 ( .A1(G286), .A2(G868), .ZN(n648) );
  INV_X1 U720 ( .A(G868), .ZN(n713) );
  NAND2_X1 U721 ( .A1(G299), .A2(n713), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(G297) );
  NAND2_X1 U723 ( .A1(n649), .A2(G559), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n650), .A2(n1012), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U726 ( .A1(G868), .A2(n1016), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n1012), .A2(G868), .ZN(n652) );
  NOR2_X1 U728 ( .A1(G559), .A2(n652), .ZN(n653) );
  NOR2_X1 U729 ( .A1(n654), .A2(n653), .ZN(G282) );
  NAND2_X1 U730 ( .A1(G99), .A2(n929), .ZN(n656) );
  NAND2_X1 U731 ( .A1(G111), .A2(n933), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n657), .A2(G123), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n658), .B(KEYINPUT18), .ZN(n660) );
  BUF_X1 U735 ( .A(n601), .Z(n930) );
  NAND2_X1 U736 ( .A1(G135), .A2(n930), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U738 ( .A(KEYINPUT83), .B(n661), .Z(n662) );
  NOR2_X1 U739 ( .A1(n663), .A2(n662), .ZN(n950) );
  XOR2_X1 U740 ( .A(n950), .B(G2096), .Z(n664) );
  XNOR2_X1 U741 ( .A(KEYINPUT84), .B(n664), .ZN(n665) );
  NOR2_X1 U742 ( .A1(G2100), .A2(n665), .ZN(n666) );
  XNOR2_X1 U743 ( .A(KEYINPUT85), .B(n666), .ZN(G156) );
  NAND2_X1 U744 ( .A1(G80), .A2(n696), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n667), .B(KEYINPUT86), .ZN(n674) );
  NAND2_X1 U746 ( .A1(G67), .A2(n690), .ZN(n669) );
  NAND2_X1 U747 ( .A1(G93), .A2(n693), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n669), .A2(n668), .ZN(n672) );
  NAND2_X1 U749 ( .A1(G55), .A2(n692), .ZN(n670) );
  XNOR2_X1 U750 ( .A(KEYINPUT87), .B(n670), .ZN(n671) );
  NOR2_X1 U751 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n714) );
  NAND2_X1 U753 ( .A1(n1012), .A2(G559), .ZN(n710) );
  XNOR2_X1 U754 ( .A(n1016), .B(n710), .ZN(n675) );
  NOR2_X1 U755 ( .A1(G860), .A2(n675), .ZN(n676) );
  XOR2_X1 U756 ( .A(n714), .B(n676), .Z(G145) );
  NAND2_X1 U757 ( .A1(G47), .A2(n692), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G60), .A2(n690), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U760 ( .A(KEYINPUT69), .B(n679), .ZN(n683) );
  NAND2_X1 U761 ( .A1(G85), .A2(n693), .ZN(n681) );
  NAND2_X1 U762 ( .A1(G72), .A2(n696), .ZN(n680) );
  AND2_X1 U763 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U764 ( .A1(n683), .A2(n682), .ZN(G290) );
  NAND2_X1 U765 ( .A1(G49), .A2(n692), .ZN(n685) );
  NAND2_X1 U766 ( .A1(G74), .A2(G651), .ZN(n684) );
  NAND2_X1 U767 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U768 ( .A1(n690), .A2(n686), .ZN(n689) );
  NAND2_X1 U769 ( .A1(n687), .A2(G87), .ZN(n688) );
  NAND2_X1 U770 ( .A1(n689), .A2(n688), .ZN(G288) );
  NAND2_X1 U771 ( .A1(G61), .A2(n690), .ZN(n691) );
  XNOR2_X1 U772 ( .A(n691), .B(KEYINPUT88), .ZN(n701) );
  NAND2_X1 U773 ( .A1(G48), .A2(n692), .ZN(n695) );
  NAND2_X1 U774 ( .A1(G86), .A2(n693), .ZN(n694) );
  NAND2_X1 U775 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U776 ( .A1(n696), .A2(G73), .ZN(n697) );
  XOR2_X1 U777 ( .A(KEYINPUT2), .B(n697), .Z(n698) );
  NOR2_X1 U778 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U779 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U780 ( .A(KEYINPUT89), .B(n702), .Z(G305) );
  XNOR2_X1 U781 ( .A(KEYINPUT19), .B(G290), .ZN(n703) );
  XNOR2_X1 U782 ( .A(n703), .B(G288), .ZN(n706) );
  XNOR2_X1 U783 ( .A(G303), .B(G305), .ZN(n704) );
  XNOR2_X1 U784 ( .A(n704), .B(n714), .ZN(n705) );
  XNOR2_X1 U785 ( .A(n706), .B(n705), .ZN(n708) );
  XNOR2_X1 U786 ( .A(G299), .B(KEYINPUT91), .ZN(n707) );
  XNOR2_X1 U787 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U788 ( .A(n709), .B(n1016), .ZN(n880) );
  XNOR2_X1 U789 ( .A(KEYINPUT92), .B(n880), .ZN(n711) );
  XNOR2_X1 U790 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U791 ( .A1(n712), .A2(G868), .ZN(n716) );
  NAND2_X1 U792 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U793 ( .A1(n716), .A2(n715), .ZN(G295) );
  NAND2_X1 U794 ( .A1(G2078), .A2(G2084), .ZN(n717) );
  XOR2_X1 U795 ( .A(KEYINPUT20), .B(n717), .Z(n718) );
  NAND2_X1 U796 ( .A1(G2090), .A2(n718), .ZN(n719) );
  XNOR2_X1 U797 ( .A(KEYINPUT21), .B(n719), .ZN(n720) );
  NAND2_X1 U798 ( .A1(n720), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U799 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U800 ( .A1(G69), .A2(G57), .ZN(n721) );
  NOR2_X1 U801 ( .A1(G236), .A2(n721), .ZN(n722) );
  XNOR2_X1 U802 ( .A(KEYINPUT96), .B(n722), .ZN(n723) );
  NAND2_X1 U803 ( .A1(n723), .A2(G108), .ZN(n878) );
  NAND2_X1 U804 ( .A1(n878), .A2(G567), .ZN(n731) );
  XOR2_X1 U805 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n725) );
  NAND2_X1 U806 ( .A1(G132), .A2(G82), .ZN(n724) );
  XNOR2_X1 U807 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U808 ( .A1(n726), .A2(G218), .ZN(n727) );
  XOR2_X1 U809 ( .A(KEYINPUT94), .B(n727), .Z(n728) );
  NOR2_X1 U810 ( .A1(G221), .A2(n728), .ZN(n729) );
  XNOR2_X1 U811 ( .A(KEYINPUT95), .B(n729), .ZN(n879) );
  NAND2_X1 U812 ( .A1(n879), .A2(G2106), .ZN(n730) );
  NAND2_X1 U813 ( .A1(n731), .A2(n730), .ZN(n949) );
  NAND2_X1 U814 ( .A1(G483), .A2(G661), .ZN(n732) );
  NOR2_X1 U815 ( .A1(n949), .A2(n732), .ZN(n877) );
  NAND2_X1 U816 ( .A1(n877), .A2(G36), .ZN(G176) );
  NAND2_X1 U817 ( .A1(G160), .A2(G40), .ZN(n737) );
  INV_X1 U818 ( .A(n737), .ZN(n734) );
  INV_X1 U819 ( .A(n830), .ZN(n738) );
  XNOR2_X1 U820 ( .A(G1996), .B(KEYINPUT103), .ZN(n981) );
  XNOR2_X1 U821 ( .A(n736), .B(KEYINPUT66), .ZN(n743) );
  NAND2_X1 U822 ( .A1(n743), .A2(n1012), .ZN(n742) );
  NOR2_X1 U823 ( .A1(n759), .A2(G1348), .ZN(n740) );
  NOR2_X1 U824 ( .A1(G2067), .A2(n771), .ZN(n739) );
  NOR2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U826 ( .A1(n742), .A2(n741), .ZN(n747) );
  INV_X1 U827 ( .A(n743), .ZN(n745) );
  INV_X1 U828 ( .A(n1012), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U830 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U831 ( .A1(n759), .A2(G2072), .ZN(n749) );
  XNOR2_X1 U832 ( .A(n749), .B(KEYINPUT27), .ZN(n751) );
  XOR2_X1 U833 ( .A(G1956), .B(KEYINPUT102), .Z(n1033) );
  NOR2_X1 U834 ( .A1(n759), .A2(n1033), .ZN(n750) );
  NOR2_X1 U835 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n754), .A2(n1002), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n753), .A2(n752), .ZN(n757) );
  NOR2_X1 U838 ( .A1(n754), .A2(n1002), .ZN(n755) );
  XOR2_X1 U839 ( .A(n755), .B(KEYINPUT28), .Z(n756) );
  XNOR2_X1 U840 ( .A(G2078), .B(KEYINPUT25), .ZN(n982) );
  NAND2_X1 U841 ( .A1(n759), .A2(n982), .ZN(n758) );
  XNOR2_X1 U842 ( .A(n758), .B(KEYINPUT101), .ZN(n761) );
  NOR2_X1 U843 ( .A1(n759), .A2(G1961), .ZN(n760) );
  NOR2_X1 U844 ( .A1(n761), .A2(n760), .ZN(n765) );
  NAND2_X1 U845 ( .A1(n771), .A2(G8), .ZN(n809) );
  NOR2_X1 U846 ( .A1(G1966), .A2(n809), .ZN(n782) );
  NOR2_X1 U847 ( .A1(n771), .A2(G2084), .ZN(n779) );
  NOR2_X1 U848 ( .A1(n782), .A2(n779), .ZN(n762) );
  NAND2_X1 U849 ( .A1(G8), .A2(n762), .ZN(n763) );
  XNOR2_X1 U850 ( .A(KEYINPUT30), .B(n763), .ZN(n764) );
  NOR2_X1 U851 ( .A1(G168), .A2(n764), .ZN(n767) );
  AND2_X1 U852 ( .A1(G301), .A2(n765), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U854 ( .A(n769), .B(KEYINPUT105), .ZN(n780) );
  NAND2_X1 U855 ( .A1(n780), .A2(G286), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT106), .ZN(n776) );
  NOR2_X1 U857 ( .A1(G1971), .A2(n809), .ZN(n773) );
  NOR2_X1 U858 ( .A1(G2090), .A2(n771), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n774), .A2(G303), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U862 ( .A1(n777), .A2(G8), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT32), .ZN(n786) );
  NAND2_X1 U864 ( .A1(G8), .A2(n779), .ZN(n784) );
  INV_X1 U865 ( .A(n780), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U867 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U868 ( .A1(n786), .A2(n785), .ZN(n788) );
  INV_X1 U869 ( .A(KEYINPUT107), .ZN(n787) );
  XNOR2_X1 U870 ( .A(n788), .B(n787), .ZN(n805) );
  NOR2_X1 U871 ( .A1(G1976), .A2(G288), .ZN(n794) );
  NOR2_X1 U872 ( .A1(G303), .A2(G1971), .ZN(n789) );
  NOR2_X1 U873 ( .A1(n794), .A2(n789), .ZN(n1007) );
  NAND2_X1 U874 ( .A1(n805), .A2(n1007), .ZN(n791) );
  INV_X1 U875 ( .A(n809), .ZN(n803) );
  NAND2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  AND2_X1 U877 ( .A1(n803), .A2(n1001), .ZN(n790) );
  XNOR2_X1 U878 ( .A(n792), .B(KEYINPUT64), .ZN(n793) );
  NOR2_X1 U879 ( .A1(n793), .A2(KEYINPUT33), .ZN(n801) );
  INV_X1 U880 ( .A(KEYINPUT33), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n803), .A2(n794), .ZN(n795) );
  NOR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U883 ( .A(n797), .B(KEYINPUT108), .Z(n799) );
  XNOR2_X1 U884 ( .A(G1981), .B(G305), .ZN(n1021) );
  INV_X1 U885 ( .A(n1021), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U887 ( .A1(G1981), .A2(G305), .ZN(n802) );
  XNOR2_X1 U888 ( .A(KEYINPUT24), .B(n802), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n804), .A2(n803), .ZN(n811) );
  NOR2_X1 U890 ( .A1(G2090), .A2(G303), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G8), .A2(n806), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n805), .A2(n807), .ZN(n808) );
  NAND2_X1 U893 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n811), .A2(n810), .ZN(n853) );
  NAND2_X1 U895 ( .A1(G141), .A2(n930), .ZN(n812) );
  XNOR2_X1 U896 ( .A(n812), .B(KEYINPUT100), .ZN(n819) );
  NAND2_X1 U897 ( .A1(G129), .A2(n657), .ZN(n814) );
  NAND2_X1 U898 ( .A1(G117), .A2(n933), .ZN(n813) );
  NAND2_X1 U899 ( .A1(n814), .A2(n813), .ZN(n817) );
  NAND2_X1 U900 ( .A1(n929), .A2(G105), .ZN(n815) );
  XOR2_X1 U901 ( .A(KEYINPUT38), .B(n815), .Z(n816) );
  NOR2_X1 U902 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n819), .A2(n818), .ZN(n920) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n920), .ZN(n820) );
  XOR2_X1 U905 ( .A(KEYINPUT109), .B(n820), .Z(n958) );
  NAND2_X1 U906 ( .A1(G95), .A2(n929), .ZN(n822) );
  NAND2_X1 U907 ( .A1(G131), .A2(n930), .ZN(n821) );
  NAND2_X1 U908 ( .A1(n822), .A2(n821), .ZN(n826) );
  NAND2_X1 U909 ( .A1(G119), .A2(n657), .ZN(n824) );
  NAND2_X1 U910 ( .A1(G107), .A2(n933), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U912 ( .A1(n826), .A2(n825), .ZN(n919) );
  INV_X1 U913 ( .A(G1991), .ZN(n976) );
  NOR2_X1 U914 ( .A1(n919), .A2(n976), .ZN(n828) );
  AND2_X1 U915 ( .A1(n920), .A2(G1996), .ZN(n827) );
  NOR2_X1 U916 ( .A1(n828), .A2(n827), .ZN(n956) );
  NOR2_X1 U917 ( .A1(n830), .A2(n829), .ZN(n854) );
  INV_X1 U918 ( .A(n854), .ZN(n831) );
  NOR2_X1 U919 ( .A1(n956), .A2(n831), .ZN(n855) );
  AND2_X1 U920 ( .A1(n976), .A2(n919), .ZN(n951) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n832) );
  NOR2_X1 U922 ( .A1(n951), .A2(n832), .ZN(n833) );
  NOR2_X1 U923 ( .A1(n855), .A2(n833), .ZN(n834) );
  NOR2_X1 U924 ( .A1(n958), .A2(n834), .ZN(n835) );
  XNOR2_X1 U925 ( .A(n835), .B(KEYINPUT39), .ZN(n847) );
  XNOR2_X1 U926 ( .A(G2067), .B(KEYINPUT37), .ZN(n836) );
  XNOR2_X1 U927 ( .A(n836), .B(KEYINPUT98), .ZN(n848) );
  NAND2_X1 U928 ( .A1(n930), .A2(G140), .ZN(n837) );
  XOR2_X1 U929 ( .A(KEYINPUT99), .B(n837), .Z(n839) );
  NAND2_X1 U930 ( .A1(n929), .A2(G104), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U932 ( .A(KEYINPUT34), .B(n840), .ZN(n845) );
  NAND2_X1 U933 ( .A1(G128), .A2(n657), .ZN(n842) );
  NAND2_X1 U934 ( .A1(G116), .A2(n933), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U936 ( .A(KEYINPUT35), .B(n843), .Z(n844) );
  NOR2_X1 U937 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U938 ( .A(KEYINPUT36), .B(n846), .ZN(n924) );
  NOR2_X1 U939 ( .A1(n848), .A2(n924), .ZN(n960) );
  NAND2_X1 U940 ( .A1(n854), .A2(n960), .ZN(n857) );
  NAND2_X1 U941 ( .A1(n847), .A2(n857), .ZN(n849) );
  NAND2_X1 U942 ( .A1(n848), .A2(n924), .ZN(n962) );
  NAND2_X1 U943 ( .A1(n849), .A2(n962), .ZN(n850) );
  XNOR2_X1 U944 ( .A(KEYINPUT110), .B(n850), .ZN(n851) );
  NAND2_X1 U945 ( .A1(n851), .A2(n854), .ZN(n861) );
  INV_X1 U946 ( .A(n861), .ZN(n852) );
  XNOR2_X1 U947 ( .A(G1986), .B(G290), .ZN(n1009) );
  AND2_X1 U948 ( .A1(n1009), .A2(n854), .ZN(n859) );
  INV_X1 U949 ( .A(n855), .ZN(n856) );
  NAND2_X1 U950 ( .A1(n857), .A2(n856), .ZN(n858) );
  OR2_X1 U951 ( .A1(n859), .A2(n858), .ZN(n860) );
  AND2_X1 U952 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U953 ( .A(G1348), .B(G2454), .ZN(n863) );
  XNOR2_X1 U954 ( .A(n863), .B(G2430), .ZN(n864) );
  XNOR2_X1 U955 ( .A(n864), .B(G1341), .ZN(n870) );
  XOR2_X1 U956 ( .A(G2443), .B(G2427), .Z(n866) );
  XNOR2_X1 U957 ( .A(G2438), .B(G2446), .ZN(n865) );
  XNOR2_X1 U958 ( .A(n866), .B(n865), .ZN(n868) );
  XOR2_X1 U959 ( .A(G2451), .B(G2435), .Z(n867) );
  XNOR2_X1 U960 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U961 ( .A(n870), .B(n869), .ZN(n871) );
  NAND2_X1 U962 ( .A1(n871), .A2(G14), .ZN(n945) );
  XNOR2_X1 U963 ( .A(KEYINPUT111), .B(n945), .ZN(G401) );
  NAND2_X1 U964 ( .A1(n872), .A2(G2106), .ZN(n873) );
  XNOR2_X1 U965 ( .A(n873), .B(KEYINPUT112), .ZN(G217) );
  AND2_X1 U966 ( .A1(G15), .A2(G2), .ZN(n874) );
  NAND2_X1 U967 ( .A1(G661), .A2(n874), .ZN(G259) );
  NAND2_X1 U968 ( .A1(G3), .A2(G1), .ZN(n875) );
  XOR2_X1 U969 ( .A(KEYINPUT113), .B(n875), .Z(n876) );
  NAND2_X1 U970 ( .A1(n877), .A2(n876), .ZN(G188) );
  XOR2_X1 U971 ( .A(G69), .B(KEYINPUT114), .Z(G235) );
  INV_X1 U973 ( .A(G132), .ZN(G219) );
  INV_X1 U974 ( .A(G108), .ZN(G238) );
  INV_X1 U975 ( .A(G82), .ZN(G220) );
  INV_X1 U976 ( .A(G57), .ZN(G237) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(G325) );
  INV_X1 U978 ( .A(G325), .ZN(G261) );
  XOR2_X1 U979 ( .A(n880), .B(G286), .Z(n882) );
  XNOR2_X1 U980 ( .A(G171), .B(n1012), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U982 ( .A1(G37), .A2(n883), .ZN(G397) );
  XOR2_X1 U983 ( .A(G1981), .B(G1961), .Z(n885) );
  XNOR2_X1 U984 ( .A(G1986), .B(G1966), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U986 ( .A(n886), .B(G2474), .Z(n888) );
  XNOR2_X1 U987 ( .A(G1996), .B(G1991), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT41), .B(G1976), .Z(n890) );
  XNOR2_X1 U990 ( .A(G1956), .B(G1971), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(G229) );
  XOR2_X1 U993 ( .A(KEYINPUT42), .B(G2072), .Z(n894) );
  XNOR2_X1 U994 ( .A(G2067), .B(G2078), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U996 ( .A(n895), .B(G2100), .Z(n897) );
  XNOR2_X1 U997 ( .A(G2090), .B(G2084), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n901) );
  XOR2_X1 U999 ( .A(G2096), .B(KEYINPUT43), .Z(n899) );
  XNOR2_X1 U1000 ( .A(G2678), .B(KEYINPUT115), .ZN(n898) );
  XNOR2_X1 U1001 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U1002 ( .A(n901), .B(n900), .Z(G227) );
  NAND2_X1 U1003 ( .A1(n657), .A2(G124), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n902), .B(KEYINPUT44), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(G136), .A2(n930), .ZN(n903) );
  NAND2_X1 U1006 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(KEYINPUT116), .B(n905), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(G100), .A2(n929), .ZN(n907) );
  NAND2_X1 U1009 ( .A1(G112), .A2(n933), .ZN(n906) );
  NAND2_X1 U1010 ( .A1(n907), .A2(n906), .ZN(n908) );
  NOR2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(G162) );
  NAND2_X1 U1012 ( .A1(G130), .A2(n657), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(G118), .A2(n933), .ZN(n910) );
  NAND2_X1 U1014 ( .A1(n911), .A2(n910), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(G106), .A2(n929), .ZN(n913) );
  NAND2_X1 U1016 ( .A1(G142), .A2(n930), .ZN(n912) );
  NAND2_X1 U1017 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1018 ( .A(KEYINPUT117), .B(n914), .ZN(n915) );
  XNOR2_X1 U1019 ( .A(KEYINPUT45), .B(n915), .ZN(n916) );
  NOR2_X1 U1020 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1021 ( .A(n950), .B(n918), .ZN(n928) );
  XOR2_X1 U1022 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n922) );
  XOR2_X1 U1023 ( .A(n920), .B(n919), .Z(n921) );
  XNOR2_X1 U1024 ( .A(n922), .B(n921), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(n924), .B(n923), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(G164), .B(G160), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(n926), .B(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(n928), .B(n927), .ZN(n941) );
  NAND2_X1 U1029 ( .A1(G103), .A2(n929), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(G139), .A2(n930), .ZN(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n939) );
  NAND2_X1 U1032 ( .A1(n933), .A2(G115), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT118), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(G127), .A2(n657), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1036 ( .A(KEYINPUT47), .B(n937), .Z(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n963) );
  XOR2_X1 U1038 ( .A(n963), .B(G162), .Z(n940) );
  XNOR2_X1 U1039 ( .A(n941), .B(n940), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(G37), .A2(n942), .ZN(G395) );
  NOR2_X1 U1041 ( .A1(G229), .A2(G227), .ZN(n943) );
  XOR2_X1 U1042 ( .A(KEYINPUT49), .B(n943), .Z(n944) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(G397), .A2(n946), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(G395), .A2(n949), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(G225) );
  INV_X1 U1047 ( .A(G225), .ZN(G308) );
  INV_X1 U1048 ( .A(n949), .ZN(G319) );
  XNOR2_X1 U1049 ( .A(G160), .B(G2084), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(n954), .B(KEYINPUT119), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n972) );
  XOR2_X1 U1054 ( .A(G2090), .B(G162), .Z(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1056 ( .A(KEYINPUT51), .B(n959), .Z(n970) );
  INV_X1 U1057 ( .A(n960), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n968) );
  XOR2_X1 U1059 ( .A(G2072), .B(n963), .Z(n965) );
  XOR2_X1 U1060 ( .A(G164), .B(G2078), .Z(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1062 ( .A(KEYINPUT50), .B(n966), .Z(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT52), .B(n973), .ZN(n974) );
  INV_X1 U1067 ( .A(KEYINPUT55), .ZN(n996) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n996), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(G29), .ZN(n1059) );
  XNOR2_X1 U1070 ( .A(G2090), .B(G35), .ZN(n991) );
  XNOR2_X1 U1071 ( .A(G25), .B(n976), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n977), .A2(G28), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G2067), .B(G26), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(G2072), .B(G33), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(KEYINPUT120), .B(n980), .ZN(n986) );
  XOR2_X1 U1077 ( .A(n981), .B(G32), .Z(n984) );
  XOR2_X1 U1078 ( .A(n982), .B(G27), .Z(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT53), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n994) );
  XOR2_X1 U1084 ( .A(G2084), .B(KEYINPUT54), .Z(n992) );
  XNOR2_X1 U1085 ( .A(G34), .B(n992), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n996), .B(n995), .ZN(n998) );
  INV_X1 U1088 ( .A(G29), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(G11), .A2(n999), .ZN(n1057) );
  XNOR2_X1 U1091 ( .A(G16), .B(KEYINPUT56), .ZN(n1026) );
  NAND2_X1 U1092 ( .A1(G303), .A2(G1971), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(n1002), .B(G1956), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(G171), .B(G1961), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1005), .B(KEYINPUT122), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G1348), .B(n1012), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT121), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(G1341), .B(n1016), .Z(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT123), .B(n1019), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(G1966), .B(G168), .Z(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT57), .B(n1022), .Z(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1055) );
  INV_X1 U1112 ( .A(G16), .ZN(n1053) );
  XOR2_X1 U1113 ( .A(G1986), .B(G24), .Z(n1030) );
  XNOR2_X1 U1114 ( .A(G1971), .B(G22), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(G23), .B(G1976), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1032) );
  XOR2_X1 U1118 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n1031) );
  XNOR2_X1 U1119 ( .A(n1032), .B(n1031), .ZN(n1049) );
  XNOR2_X1 U1120 ( .A(G1961), .B(G5), .ZN(n1047) );
  XNOR2_X1 U1121 ( .A(G1966), .B(G21), .ZN(n1044) );
  XOR2_X1 U1122 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n1042) );
  XNOR2_X1 U1123 ( .A(n1033), .B(G20), .ZN(n1037) );
  XNOR2_X1 U1124 ( .A(G1341), .B(G19), .ZN(n1035) );
  XNOR2_X1 U1125 ( .A(G6), .B(G1981), .ZN(n1034) );
  NOR2_X1 U1126 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1127 ( .A1(n1037), .A2(n1036), .ZN(n1040) );
  XOR2_X1 U1128 ( .A(KEYINPUT59), .B(G1348), .Z(n1038) );
  XNOR2_X1 U1129 ( .A(G4), .B(n1038), .ZN(n1039) );
  NOR2_X1 U1130 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1131 ( .A(n1042), .B(n1041), .ZN(n1043) );
  NOR2_X1 U1132 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1133 ( .A(KEYINPUT125), .B(n1045), .ZN(n1046) );
  NOR2_X1 U1134 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NAND2_X1 U1135 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XNOR2_X1 U1136 ( .A(n1050), .B(KEYINPUT61), .ZN(n1051) );
  XNOR2_X1 U1137 ( .A(KEYINPUT127), .B(n1051), .ZN(n1052) );
  NAND2_X1 U1138 ( .A1(n1053), .A2(n1052), .ZN(n1054) );
  NAND2_X1 U1139 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  NOR2_X1 U1140 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
  NAND2_X1 U1141 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
  XOR2_X1 U1142 ( .A(KEYINPUT62), .B(n1060), .Z(G311) );
  INV_X1 U1143 ( .A(G311), .ZN(G150) );
endmodule

