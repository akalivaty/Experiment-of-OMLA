//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139, new_n1140, new_n1141;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n465), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n470), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G137), .A3(new_n462), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n467), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(new_n479), .ZN(G160));
  INV_X1    g055(.A(new_n475), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n462), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n481), .A2(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(G136), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT69), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(new_n493), .A3(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT70), .B1(new_n462), .B2(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n465), .A2(new_n471), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n500), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n507), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OAI221_X1 g092(.A(new_n509), .B1(new_n514), .B2(new_n515), .C1(new_n516), .C2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  XOR2_X1   g094(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n511), .A2(new_n512), .B1(new_n506), .B2(new_n507), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G89), .B1(new_n508), .B2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT72), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n522), .A2(new_n528), .A3(new_n525), .A4(new_n523), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(G168));
  AOI22_X1  g105(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n517), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n508), .A2(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n514), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  XNOR2_X1  g111(.A(KEYINPUT73), .B(G43), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n524), .A2(G81), .B1(new_n508), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n517), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT74), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g118(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n544));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(new_n513), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT78), .B(G65), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n514), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n508), .A2(G53), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT77), .B1(new_n556), .B2(KEYINPUT76), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(KEYINPUT77), .B2(new_n556), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n524), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n508), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  INV_X1    g144(.A(G61), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n511), .B2(new_n512), .ZN(new_n571));
  AND2_X1   g146(.A1(G73), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(KEYINPUT79), .B(G651), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n524), .A2(G86), .B1(new_n508), .B2(G48), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(G72), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G60), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n549), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n517), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n582), .B2(new_n581), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT81), .B(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n524), .A2(new_n585), .B1(new_n508), .B2(G47), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n524), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  AOI22_X1  g165(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n517), .B1(new_n591), .B2(KEYINPUT82), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(KEYINPUT82), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n508), .A2(G54), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G284));
  XOR2_X1   g172(.A(G284), .B(KEYINPUT83), .Z(G321));
  OAI21_X1  g173(.A(KEYINPUT84), .B1(new_n562), .B2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  MUX2_X1   g175(.A(KEYINPUT84), .B(new_n599), .S(new_n600), .Z(G297));
  XOR2_X1   g176(.A(G297), .B(KEYINPUT85), .Z(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n596), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g183(.A1(new_n465), .A2(new_n471), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n477), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  INV_X1    g187(.A(G2100), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  AOI22_X1  g190(.A1(G123), .A2(new_n482), .B1(new_n487), .B2(G135), .ZN(new_n616));
  NOR3_X1   g191(.A1(new_n462), .A2(KEYINPUT86), .A3(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT86), .B1(new_n462), .B2(G111), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n616), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n614), .A2(new_n615), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n633), .A2(new_n636), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(G401));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(new_n613), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n644), .B2(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(new_n621), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n657), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  AOI211_X1 g236(.A(new_n659), .B(new_n661), .C1(new_n654), .C2(new_n658), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  XOR2_X1   g238(.A(G1981), .B(G1986), .Z(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n663), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NOR2_X1   g246(.A1(G171), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(G5), .B2(new_n671), .ZN(new_n673));
  INV_X1    g248(.A(G1961), .ZN(new_n674));
  INV_X1    g249(.A(G29), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G32), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n482), .A2(G129), .ZN(new_n677));
  NAND3_X1  g252(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT26), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n487), .A2(G141), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n477), .A2(G105), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n676), .B1(new_n684), .B2(new_n675), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT27), .B(G1996), .Z(new_n686));
  AOI22_X1  g261(.A1(new_n673), .A2(new_n674), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n675), .A2(KEYINPUT89), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n675), .A2(KEYINPUT89), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT24), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n691), .A2(G34), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(G34), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G160), .B2(G29), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n687), .B1(G2084), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT100), .ZN(new_n697));
  INV_X1    g272(.A(new_n690), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G26), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n487), .A2(G140), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n482), .A2(G128), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g279(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n705));
  OAI221_X1 g280(.A(G2104), .B1(G116), .B2(new_n462), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n701), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(new_n675), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n700), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G2067), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G4), .A2(G16), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n595), .B2(new_n671), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT95), .B(G1348), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n690), .A2(G35), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G162), .B2(new_n690), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT29), .B(G2090), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n697), .A2(new_n713), .A3(new_n719), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n671), .A2(G20), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT23), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n562), .B2(new_n671), .ZN(new_n727));
  INV_X1    g302(.A(G1956), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n671), .A2(G21), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G168), .B2(new_n671), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n731), .A2(G1966), .B1(G2084), .B2(new_n695), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n729), .B(new_n732), .C1(G1966), .C2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n671), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n541), .B2(new_n671), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1341), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n685), .A2(new_n686), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n698), .A2(G27), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT101), .Z(new_n739));
  INV_X1    g314(.A(G164), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n690), .ZN(new_n741));
  INV_X1    g316(.A(G2078), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  OR2_X1    g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n744), .A2(new_n675), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n747), .B1(new_n620), .B2(new_n698), .C1(new_n673), .C2(new_n674), .ZN(new_n748));
  OR4_X1    g323(.A1(new_n736), .A2(new_n737), .A3(new_n743), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n675), .A2(G33), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT25), .ZN(new_n751));
  NAND2_X1  g326(.A1(G103), .A2(G2104), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(G2105), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n487), .A2(G139), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n609), .A2(G127), .ZN(new_n756));
  NAND2_X1  g331(.A1(G115), .A2(G2104), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n462), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n750), .B1(new_n761), .B2(new_n675), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT99), .B(G2072), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n724), .A2(new_n733), .A3(new_n749), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G305), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G6), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT32), .B(G1981), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n671), .A2(G22), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT93), .Z(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n671), .ZN(new_n774));
  INV_X1    g349(.A(G1971), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n768), .A2(new_n770), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G23), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT92), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G288), .B2(new_n671), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT33), .B(G1976), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n771), .A2(new_n776), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  MUX2_X1   g361(.A(G24), .B(G290), .S(G16), .Z(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G1986), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(G1986), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n690), .A2(G25), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n487), .A2(G131), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n482), .A2(G119), .ZN(new_n792));
  OR2_X1    g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n690), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT35), .B(G1991), .Z(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT90), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n797), .B(new_n799), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n788), .A2(new_n789), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n785), .A2(new_n786), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT36), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n765), .A2(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  AOI22_X1  g380(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n517), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n508), .A2(G55), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT102), .B(G93), .Z(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n514), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G860), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT37), .ZN(new_n814));
  MUX2_X1   g389(.A(new_n541), .B(new_n540), .S(new_n811), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT38), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n595), .A2(new_n603), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT103), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n814), .B1(new_n821), .B2(new_n822), .ZN(G145));
  XNOR2_X1  g398(.A(new_n761), .B(new_n684), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n611), .B(new_n795), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT105), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n498), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n496), .A2(KEYINPUT105), .A3(new_n497), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(new_n500), .B2(new_n503), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n707), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n482), .A2(G130), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT106), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n487), .A2(G142), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n462), .A2(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n831), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n826), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(G160), .B(KEYINPUT104), .Z(new_n840));
  XNOR2_X1  g415(.A(G162), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n620), .ZN(new_n842));
  AOI21_X1  g417(.A(G37), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n839), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g420(.A(G290), .B(G305), .ZN(new_n846));
  XNOR2_X1  g421(.A(G303), .B(G288), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT42), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n815), .B(new_n605), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n595), .A2(KEYINPUT107), .A3(new_n562), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n562), .B2(new_n595), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT107), .B1(new_n595), .B2(new_n562), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT41), .B1(new_n853), .B2(new_n854), .ZN(new_n857));
  OR3_X1    g432(.A1(new_n853), .A2(KEYINPUT41), .A3(new_n854), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n851), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n850), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n849), .A2(new_n856), .A3(new_n859), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(G868), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(G868), .B2(new_n811), .ZN(G295));
  XNOR2_X1  g441(.A(G295), .B(KEYINPUT108), .ZN(G331));
  XNOR2_X1  g442(.A(G168), .B(G301), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n815), .B(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n855), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n858), .A3(new_n857), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n848), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n848), .A3(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT44), .ZN(G397));
  INV_X1    g454(.A(KEYINPUT126), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n684), .B(G1996), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n707), .B(G2067), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n795), .B(new_n798), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n503), .A2(new_n500), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n496), .A2(KEYINPUT105), .A3(new_n497), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT105), .B1(new_n496), .B2(new_n497), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G1384), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n472), .A2(new_n473), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G2105), .ZN(new_n895));
  INV_X1    g470(.A(new_n479), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(G40), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n885), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  XOR2_X1   g475(.A(G290), .B(G1986), .Z(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT109), .Z(new_n903));
  INV_X1    g478(.A(KEYINPUT49), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n575), .A2(KEYINPUT111), .A3(new_n576), .ZN(new_n905));
  NAND3_X1  g480(.A1(G305), .A2(new_n905), .A3(G1981), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G305), .B1(G1981), .B2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(G1981), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n766), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT49), .A3(new_n906), .ZN(new_n912));
  OAI21_X1  g487(.A(G8), .B1(new_n891), .B2(new_n897), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G288), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n916), .A2(G1976), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT52), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT52), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n916), .B2(G1976), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n913), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G8), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n924));
  NAND3_X1  g499(.A1(G303), .A2(G8), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g501(.A1(G303), .A2(G8), .B1(KEYINPUT110), .B2(KEYINPUT55), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n892), .A2(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n889), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n892), .B1(G164), .B2(G1384), .ZN(new_n931));
  INV_X1    g506(.A(G40), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n474), .A2(new_n479), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n775), .ZN(new_n935));
  INV_X1    g510(.A(G2090), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT50), .B1(new_n889), .B2(new_n890), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT50), .ZN(new_n938));
  NOR3_X1   g513(.A1(G164), .A2(new_n938), .A3(G1384), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n936), .B(new_n933), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  AOI211_X1 g515(.A(new_n923), .B(new_n928), .C1(new_n935), .C2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n922), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n937), .A2(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(G2084), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n933), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT112), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n740), .A2(new_n929), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n828), .A2(new_n829), .ZN(new_n948));
  AOI21_X1  g523(.A(G1384), .B1(new_n948), .B2(new_n886), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n933), .B(new_n947), .C1(new_n949), .C2(KEYINPUT45), .ZN(new_n950));
  INV_X1    g525(.A(G1966), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n496), .A2(new_n497), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n886), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n957));
  INV_X1    g532(.A(new_n945), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n946), .A2(new_n952), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n960), .A2(G8), .A3(G168), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT63), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n935), .A2(new_n940), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(G8), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n964), .B2(new_n928), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n942), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n928), .ZN(new_n967));
  AOI211_X1 g542(.A(KEYINPUT50), .B(G1384), .C1(new_n886), .C2(new_n953), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n897), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n891), .A2(KEYINPUT50), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n970), .A3(new_n936), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n935), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n967), .B1(new_n972), .B2(G8), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n942), .A2(new_n961), .A3(KEYINPUT113), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n962), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n922), .A2(new_n941), .A3(new_n973), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT113), .B1(new_n977), .B2(new_n961), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n966), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(G305), .A2(G1981), .ZN(new_n980));
  NOR2_X1   g555(.A1(G288), .A2(G1976), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n915), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n922), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n983), .A2(new_n914), .B1(new_n984), .B2(new_n941), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT57), .B1(new_n554), .B2(new_n561), .ZN(new_n988));
  INV_X1    g563(.A(new_n561), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n551), .A2(G651), .B1(G91), .B2(new_n524), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n954), .A2(new_n938), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n933), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n938), .B1(new_n889), .B2(new_n890), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n728), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT56), .B(G2072), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n930), .A2(new_n931), .A3(new_n933), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n993), .B1(new_n997), .B2(new_n999), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n718), .B1(new_n956), .B2(new_n933), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n891), .A2(new_n897), .A3(G2067), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n596), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT114), .B(new_n596), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1001), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n988), .A2(new_n992), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1956), .B1(new_n969), .B2(new_n970), .ZN(new_n1011));
  INV_X1    g586(.A(new_n999), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(KEYINPUT61), .A3(new_n1000), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT117), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1013), .A2(new_n1000), .A3(new_n1016), .A4(KEYINPUT61), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(KEYINPUT116), .A3(new_n1000), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT61), .B1(new_n1002), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1015), .A2(new_n1017), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n933), .B1(new_n937), .B2(new_n939), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1004), .B1(new_n1022), .B2(new_n717), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1023), .A2(KEYINPUT60), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n949), .A2(new_n712), .A3(new_n933), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n938), .B1(new_n830), .B2(G1384), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n897), .B1(new_n1026), .B2(new_n955), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT60), .B(new_n1025), .C1(new_n1027), .C2(new_n718), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n596), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(KEYINPUT60), .A3(new_n595), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1996), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n930), .A2(new_n931), .A3(new_n1032), .A4(new_n933), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT58), .B(G1341), .Z(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n891), .B2(new_n897), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n541), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT59), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n541), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1024), .A2(new_n1031), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n987), .B(new_n1009), .C1(new_n1021), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1020), .A2(new_n1018), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1031), .A2(new_n1024), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1009), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT118), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT121), .B(G1961), .Z(new_n1053));
  NAND2_X1  g628(.A1(new_n1022), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(G2078), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n893), .A2(new_n933), .A3(new_n947), .A4(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n930), .A2(new_n931), .A3(new_n742), .A4(new_n933), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1055), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1054), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G171), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n893), .A2(new_n933), .A3(new_n930), .A4(new_n1056), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1054), .A2(new_n1059), .A3(new_n1065), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1066), .A2(G171), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT123), .B1(new_n1060), .B2(G171), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1022), .A2(new_n1053), .B1(new_n1058), .B2(new_n1055), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(G301), .A4(new_n1057), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1069), .B1(new_n1066), .B2(G171), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1075), .A2(KEYINPUT124), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT124), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n977), .B(new_n1070), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n527), .A2(new_n529), .A3(G8), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n945), .B1(new_n1026), .B2(new_n955), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1081), .A2(new_n957), .B1(new_n950), .B2(new_n951), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n1082), .B2(new_n946), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n923), .B1(new_n1082), .B2(new_n946), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1080), .B(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT51), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1084), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1087), .A2(new_n1088), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT120), .B(KEYINPUT51), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1079), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n986), .B1(new_n1052), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1086), .B1(new_n960), .B2(G8), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1088), .B1(new_n1097), .B2(new_n1090), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1093), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1083), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(new_n1104), .A3(new_n1101), .ZN(new_n1105));
  INV_X1    g680(.A(new_n977), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n903), .B1(new_n1096), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n898), .A2(new_n1032), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT46), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n882), .A2(new_n684), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n900), .B2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(new_n1113), .B(KEYINPUT47), .Z(new_n1114));
  OR3_X1    g689(.A1(new_n900), .A2(G1986), .A3(G290), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1117), .A2(new_n899), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n883), .A2(new_n796), .A3(new_n798), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n707), .A2(new_n712), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n900), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1114), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n880), .B1(new_n1109), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n986), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1051), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1049), .A2(KEYINPUT118), .A3(new_n1050), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1106), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1102), .B(new_n1130), .C1(new_n1078), .C2(new_n1077), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1126), .B(new_n1108), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n903), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(KEYINPUT126), .A3(new_n1123), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1125), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g711(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1138));
  OAI21_X1  g712(.A(new_n669), .B1(KEYINPUT127), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g713(.A(new_n1139), .B1(KEYINPUT127), .B2(new_n1138), .ZN(new_n1140));
  NAND2_X1  g714(.A1(new_n1140), .A2(new_n844), .ZN(new_n1141));
  NOR2_X1   g715(.A1(new_n878), .A2(new_n1141), .ZN(G308));
  INV_X1    g716(.A(G308), .ZN(G225));
endmodule


