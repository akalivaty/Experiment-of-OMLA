

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U560 ( .A(n533), .B(KEYINPUT17), .ZN(n586) );
  NOR2_X2 U561 ( .A1(n592), .A2(n591), .ZN(G164) );
  BUF_X1 U562 ( .A(n586), .Z(n580) );
  BUF_X2 U563 ( .A(n576), .Z(n892) );
  INV_X1 U564 ( .A(KEYINPUT93), .ZN(n720) );
  XNOR2_X1 U565 ( .A(n774), .B(n773), .ZN(n775) );
  XOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .Z(n662) );
  AND2_X1 U567 ( .A1(n708), .A2(KEYINPUT91), .ZN(n527) );
  INV_X1 U568 ( .A(KEYINPUT92), .ZN(n711) );
  NAND2_X1 U569 ( .A1(n756), .A2(n755), .ZN(n757) );
  INV_X1 U570 ( .A(KEYINPUT100), .ZN(n773) );
  NOR2_X1 U571 ( .A1(G651), .A2(n662), .ZN(n664) );
  INV_X1 U572 ( .A(G2104), .ZN(n528) );
  NOR2_X1 U573 ( .A1(G2105), .A2(n528), .ZN(n572) );
  NAND2_X1 U574 ( .A1(G101), .A2(n572), .ZN(n529) );
  XOR2_X1 U575 ( .A(n529), .B(KEYINPUT23), .Z(n532) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n534), .ZN(n576) );
  NAND2_X1 U577 ( .A1(G125), .A2(n576), .ZN(n530) );
  XNOR2_X1 U578 ( .A(KEYINPUT64), .B(n530), .ZN(n531) );
  NAND2_X1 U579 ( .A1(n532), .A2(n531), .ZN(n539) );
  OR2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n586), .A2(G137), .ZN(n537) );
  INV_X1 U582 ( .A(G2105), .ZN(n534) );
  NOR2_X1 U583 ( .A1(n528), .A2(n534), .ZN(n571) );
  NAND2_X1 U584 ( .A1(G113), .A2(n571), .ZN(n535) );
  XOR2_X1 U585 ( .A(n535), .B(KEYINPUT65), .Z(n536) );
  NAND2_X1 U586 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X2 U587 ( .A1(n539), .A2(n538), .ZN(G160) );
  NOR2_X1 U588 ( .A1(G543), .A2(G651), .ZN(n653) );
  NAND2_X1 U589 ( .A1(G89), .A2(n653), .ZN(n540) );
  XOR2_X1 U590 ( .A(KEYINPUT4), .B(n540), .Z(n541) );
  XNOR2_X1 U591 ( .A(n541), .B(KEYINPUT69), .ZN(n544) );
  INV_X1 U592 ( .A(G651), .ZN(n546) );
  OR2_X1 U593 ( .A1(n546), .A2(n662), .ZN(n542) );
  XOR2_X2 U594 ( .A(KEYINPUT66), .B(n542), .Z(n656) );
  NAND2_X1 U595 ( .A1(G76), .A2(n656), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U597 ( .A(n545), .B(KEYINPUT5), .ZN(n552) );
  NAND2_X1 U598 ( .A1(G51), .A2(n664), .ZN(n549) );
  NOR2_X1 U599 ( .A1(G543), .A2(n546), .ZN(n547) );
  XOR2_X1 U600 ( .A(KEYINPUT1), .B(n547), .Z(n668) );
  NAND2_X1 U601 ( .A1(G63), .A2(n668), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n550), .Z(n551) );
  NAND2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U605 ( .A(n553), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U607 ( .A1(G77), .A2(n656), .ZN(n554) );
  XOR2_X1 U608 ( .A(KEYINPUT67), .B(n554), .Z(n556) );
  NAND2_X1 U609 ( .A1(n653), .A2(G90), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U611 ( .A(KEYINPUT9), .B(n557), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G52), .A2(n664), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G64), .A2(n668), .ZN(n558) );
  AND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(G301) );
  INV_X1 U616 ( .A(G301), .ZN(G171) );
  XOR2_X1 U617 ( .A(G2443), .B(G2446), .Z(n563) );
  XNOR2_X1 U618 ( .A(G2427), .B(G2451), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n563), .B(n562), .ZN(n569) );
  XOR2_X1 U620 ( .A(G2430), .B(G2454), .Z(n565) );
  XNOR2_X1 U621 ( .A(G1348), .B(G1341), .ZN(n564) );
  XNOR2_X1 U622 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U623 ( .A(G2435), .B(G2438), .Z(n566) );
  XNOR2_X1 U624 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U625 ( .A(n569), .B(n568), .Z(n570) );
  AND2_X1 U626 ( .A1(G14), .A2(n570), .ZN(G401) );
  AND2_X1 U627 ( .A1(G452), .A2(G94), .ZN(G173) );
  BUF_X1 U628 ( .A(n571), .Z(n910) );
  NAND2_X1 U629 ( .A1(G111), .A2(n910), .ZN(n574) );
  BUF_X1 U630 ( .A(n572), .Z(n913) );
  NAND2_X1 U631 ( .A1(G99), .A2(n913), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U633 ( .A(KEYINPUT70), .B(n575), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n892), .A2(G123), .ZN(n577) );
  XOR2_X1 U635 ( .A(KEYINPUT18), .B(n577), .Z(n578) );
  NOR2_X1 U636 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U637 ( .A1(n580), .A2(G135), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n582), .A2(n581), .ZN(n1011) );
  XNOR2_X1 U639 ( .A(G2096), .B(n1011), .ZN(n583) );
  OR2_X1 U640 ( .A1(G2100), .A2(n583), .ZN(G156) );
  INV_X1 U641 ( .A(G132), .ZN(G219) );
  INV_X1 U642 ( .A(G82), .ZN(G220) );
  INV_X1 U643 ( .A(G57), .ZN(G237) );
  NAND2_X1 U644 ( .A1(G114), .A2(n910), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G102), .A2(n913), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(n592) );
  NAND2_X1 U647 ( .A1(G138), .A2(n586), .ZN(n587) );
  XNOR2_X1 U648 ( .A(n587), .B(KEYINPUT84), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G126), .A2(n892), .ZN(n588) );
  XOR2_X1 U650 ( .A(KEYINPUT83), .B(n588), .Z(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n593) );
  XNOR2_X1 U653 ( .A(n593), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G223), .ZN(n850) );
  NAND2_X1 U655 ( .A1(n850), .A2(G567), .ZN(n594) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n594), .Z(G234) );
  NAND2_X1 U657 ( .A1(G56), .A2(n668), .ZN(n595) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n595), .Z(n601) );
  NAND2_X1 U659 ( .A1(n653), .A2(G81), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(KEYINPUT12), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G68), .A2(n656), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U663 ( .A(KEYINPUT13), .B(n599), .Z(n600) );
  NOR2_X1 U664 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U665 ( .A1(n664), .A2(G43), .ZN(n602) );
  NAND2_X1 U666 ( .A1(n603), .A2(n602), .ZN(n985) );
  INV_X1 U667 ( .A(G860), .ZN(n623) );
  OR2_X1 U668 ( .A1(n985), .A2(n623), .ZN(n604) );
  XNOR2_X1 U669 ( .A(KEYINPUT68), .B(n604), .ZN(G153) );
  NAND2_X1 U670 ( .A1(G868), .A2(G301), .ZN(n613) );
  NAND2_X1 U671 ( .A1(G92), .A2(n653), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G79), .A2(n656), .ZN(n605) );
  NAND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U674 ( .A1(G54), .A2(n664), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G66), .A2(n668), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U677 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U678 ( .A(KEYINPUT15), .B(n611), .Z(n987) );
  OR2_X1 U679 ( .A1(n987), .A2(G868), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(G284) );
  NAND2_X1 U681 ( .A1(G53), .A2(n664), .ZN(n615) );
  NAND2_X1 U682 ( .A1(G65), .A2(n668), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U684 ( .A1(G91), .A2(n653), .ZN(n617) );
  NAND2_X1 U685 ( .A1(G78), .A2(n656), .ZN(n616) );
  NAND2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n996) );
  INV_X1 U688 ( .A(n996), .ZN(G299) );
  INV_X1 U689 ( .A(G868), .ZN(n620) );
  NOR2_X1 U690 ( .A1(G286), .A2(n620), .ZN(n622) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n621) );
  NOR2_X1 U692 ( .A1(n622), .A2(n621), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n623), .A2(G559), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n624), .A2(n987), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U696 ( .A1(G868), .A2(n985), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n987), .A2(G868), .ZN(n626) );
  NOR2_X1 U698 ( .A1(G559), .A2(n626), .ZN(n627) );
  NOR2_X1 U699 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U700 ( .A1(G55), .A2(n664), .ZN(n630) );
  NAND2_X1 U701 ( .A1(G67), .A2(n668), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U703 ( .A1(G93), .A2(n653), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G80), .A2(n656), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n676) );
  NAND2_X1 U707 ( .A1(n987), .A2(G559), .ZN(n681) );
  XNOR2_X1 U708 ( .A(n985), .B(n681), .ZN(n635) );
  NOR2_X1 U709 ( .A1(G860), .A2(n635), .ZN(n636) );
  XOR2_X1 U710 ( .A(KEYINPUT71), .B(n636), .Z(n637) );
  XNOR2_X1 U711 ( .A(n676), .B(n637), .ZN(G145) );
  AND2_X1 U712 ( .A1(G72), .A2(n656), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G85), .A2(n653), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G47), .A2(n664), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n668), .A2(G60), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(G290) );
  NAND2_X1 U719 ( .A1(G88), .A2(n653), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G75), .A2(n656), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U722 ( .A(KEYINPUT76), .B(n646), .ZN(n649) );
  NAND2_X1 U723 ( .A1(G62), .A2(n668), .ZN(n647) );
  XNOR2_X1 U724 ( .A(KEYINPUT75), .B(n647), .ZN(n648) );
  NOR2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n664), .A2(G50), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(G303) );
  INV_X1 U728 ( .A(G303), .ZN(G166) );
  NAND2_X1 U729 ( .A1(G61), .A2(n668), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n652), .B(KEYINPUT74), .ZN(n661) );
  NAND2_X1 U731 ( .A1(G86), .A2(n653), .ZN(n655) );
  NAND2_X1 U732 ( .A1(G48), .A2(n664), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n656), .A2(G73), .ZN(n657) );
  XOR2_X1 U735 ( .A(KEYINPUT2), .B(n657), .Z(n658) );
  NOR2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(G305) );
  NAND2_X1 U738 ( .A1(G87), .A2(n662), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(KEYINPUT72), .ZN(n670) );
  NAND2_X1 U740 ( .A1(G49), .A2(n664), .ZN(n666) );
  NAND2_X1 U741 ( .A1(G74), .A2(G651), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U743 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U745 ( .A(KEYINPUT73), .B(n671), .Z(G288) );
  NOR2_X1 U746 ( .A1(G868), .A2(n676), .ZN(n672) );
  XOR2_X1 U747 ( .A(n672), .B(KEYINPUT78), .Z(n684) );
  XNOR2_X1 U748 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n674) );
  XNOR2_X1 U749 ( .A(G290), .B(n996), .ZN(n673) );
  XNOR2_X1 U750 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U751 ( .A(n676), .B(n675), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n985), .B(G166), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U754 ( .A(n679), .B(G305), .ZN(n680) );
  XNOR2_X1 U755 ( .A(n680), .B(G288), .ZN(n858) );
  XOR2_X1 U756 ( .A(n858), .B(n681), .Z(n682) );
  NAND2_X1 U757 ( .A1(G868), .A2(n682), .ZN(n683) );
  NAND2_X1 U758 ( .A1(n684), .A2(n683), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2084), .A2(G2078), .ZN(n685) );
  XNOR2_X1 U760 ( .A(n685), .B(KEYINPUT79), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n686), .B(KEYINPUT20), .ZN(n687) );
  NAND2_X1 U762 ( .A1(n687), .A2(G2090), .ZN(n688) );
  XNOR2_X1 U763 ( .A(n688), .B(KEYINPUT80), .ZN(n689) );
  XNOR2_X1 U764 ( .A(n689), .B(KEYINPUT21), .ZN(n690) );
  NAND2_X1 U765 ( .A1(n690), .A2(G2072), .ZN(n691) );
  XOR2_X1 U766 ( .A(KEYINPUT81), .B(n691), .Z(G158) );
  XNOR2_X1 U767 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U768 ( .A1(G69), .A2(G120), .ZN(n692) );
  NOR2_X1 U769 ( .A1(G237), .A2(n692), .ZN(n693) );
  NAND2_X1 U770 ( .A1(G108), .A2(n693), .ZN(n856) );
  NAND2_X1 U771 ( .A1(n856), .A2(G567), .ZN(n699) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n694) );
  XNOR2_X1 U773 ( .A(KEYINPUT22), .B(n694), .ZN(n695) );
  NAND2_X1 U774 ( .A1(n695), .A2(G96), .ZN(n696) );
  NOR2_X1 U775 ( .A1(G218), .A2(n696), .ZN(n697) );
  XOR2_X1 U776 ( .A(KEYINPUT82), .B(n697), .Z(n857) );
  NAND2_X1 U777 ( .A1(G2106), .A2(n857), .ZN(n698) );
  NAND2_X1 U778 ( .A1(n699), .A2(n698), .ZN(n931) );
  NAND2_X1 U779 ( .A1(G661), .A2(G483), .ZN(n700) );
  NOR2_X1 U780 ( .A1(n931), .A2(n700), .ZN(n855) );
  NAND2_X1 U781 ( .A1(n855), .A2(G36), .ZN(G176) );
  NAND2_X1 U782 ( .A1(G40), .A2(G160), .ZN(n701) );
  XOR2_X1 U783 ( .A(KEYINPUT85), .B(n701), .Z(n780) );
  INV_X1 U784 ( .A(n780), .ZN(n702) );
  NOR2_X1 U785 ( .A1(G164), .A2(G1384), .ZN(n781) );
  NAND2_X2 U786 ( .A1(n702), .A2(n781), .ZN(n750) );
  NAND2_X1 U787 ( .A1(G8), .A2(n750), .ZN(n838) );
  INV_X2 U788 ( .A(n750), .ZN(n733) );
  NAND2_X1 U789 ( .A1(G1996), .A2(n733), .ZN(n703) );
  XNOR2_X1 U790 ( .A(KEYINPUT26), .B(n703), .ZN(n705) );
  INV_X1 U791 ( .A(G1341), .ZN(n935) );
  NOR2_X1 U792 ( .A1(n733), .A2(n935), .ZN(n704) );
  NAND2_X1 U793 ( .A1(KEYINPUT26), .A2(n704), .ZN(n708) );
  NAND2_X1 U794 ( .A1(n705), .A2(n708), .ZN(n707) );
  INV_X1 U795 ( .A(KEYINPUT91), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U797 ( .A1(n985), .A2(n527), .ZN(n709) );
  AND2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n713) );
  NOR2_X1 U799 ( .A1(n713), .A2(n987), .ZN(n712) );
  XNOR2_X1 U800 ( .A(n712), .B(n711), .ZN(n719) );
  NAND2_X1 U801 ( .A1(n713), .A2(n987), .ZN(n717) );
  NOR2_X1 U802 ( .A1(n733), .A2(G1348), .ZN(n715) );
  NOR2_X1 U803 ( .A1(G2067), .A2(n750), .ZN(n714) );
  NOR2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U806 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U807 ( .A(n721), .B(n720), .ZN(n726) );
  NAND2_X1 U808 ( .A1(n733), .A2(G2072), .ZN(n722) );
  XNOR2_X1 U809 ( .A(n722), .B(KEYINPUT27), .ZN(n724) );
  AND2_X1 U810 ( .A1(G1956), .A2(n750), .ZN(n723) );
  NOR2_X1 U811 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U812 ( .A1(n727), .A2(n996), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U814 ( .A1(n727), .A2(n996), .ZN(n728) );
  XOR2_X1 U815 ( .A(n728), .B(KEYINPUT28), .Z(n729) );
  NAND2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n732) );
  XOR2_X1 U817 ( .A(KEYINPUT94), .B(KEYINPUT29), .Z(n731) );
  XNOR2_X1 U818 ( .A(n732), .B(n731), .ZN(n738) );
  OR2_X1 U819 ( .A1(n733), .A2(G1961), .ZN(n735) );
  XNOR2_X1 U820 ( .A(G2078), .B(KEYINPUT25), .ZN(n961) );
  NAND2_X1 U821 ( .A1(n733), .A2(n961), .ZN(n734) );
  NAND2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n739) );
  AND2_X1 U823 ( .A1(n739), .A2(G171), .ZN(n736) );
  XOR2_X1 U824 ( .A(KEYINPUT90), .B(n736), .Z(n737) );
  NAND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n749) );
  NOR2_X1 U826 ( .A1(G171), .A2(n739), .ZN(n745) );
  NOR2_X1 U827 ( .A1(G1966), .A2(n838), .ZN(n764) );
  NOR2_X1 U828 ( .A1(G2084), .A2(n750), .ZN(n761) );
  NOR2_X1 U829 ( .A1(n764), .A2(n761), .ZN(n740) );
  XOR2_X1 U830 ( .A(KEYINPUT95), .B(n740), .Z(n741) );
  NAND2_X1 U831 ( .A1(G8), .A2(n741), .ZN(n742) );
  XNOR2_X1 U832 ( .A(KEYINPUT30), .B(n742), .ZN(n743) );
  NOR2_X1 U833 ( .A1(G168), .A2(n743), .ZN(n744) );
  NOR2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n747) );
  XOR2_X1 U835 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n746) );
  XNOR2_X1 U836 ( .A(n747), .B(n746), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n762) );
  NAND2_X1 U838 ( .A1(n762), .A2(G286), .ZN(n756) );
  NOR2_X1 U839 ( .A1(G2090), .A2(n750), .ZN(n751) );
  XOR2_X1 U840 ( .A(KEYINPUT97), .B(n751), .Z(n753) );
  NOR2_X1 U841 ( .A1(G1971), .A2(n838), .ZN(n752) );
  NOR2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n754), .A2(G303), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n757), .B(KEYINPUT98), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n758), .A2(G8), .ZN(n760) );
  XOR2_X1 U846 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n759) );
  XNOR2_X1 U847 ( .A(n760), .B(n759), .ZN(n829) );
  NAND2_X1 U848 ( .A1(G8), .A2(n761), .ZN(n766) );
  INV_X1 U849 ( .A(n762), .ZN(n763) );
  NOR2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n830) );
  NAND2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n991) );
  AND2_X1 U853 ( .A1(n830), .A2(n991), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n829), .A2(n767), .ZN(n772) );
  INV_X1 U855 ( .A(n991), .ZN(n770) );
  NOR2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n990) );
  NOR2_X1 U857 ( .A1(G1971), .A2(G303), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n990), .A2(n768), .ZN(n769) );
  OR2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n774) );
  NOR2_X1 U861 ( .A1(n838), .A2(n775), .ZN(n776) );
  NOR2_X1 U862 ( .A1(KEYINPUT33), .A2(n776), .ZN(n779) );
  NAND2_X1 U863 ( .A1(n990), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U864 ( .A1(n777), .A2(n838), .ZN(n778) );
  NOR2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n827) );
  XOR2_X1 U866 ( .A(G1981), .B(G305), .Z(n980) );
  NOR2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n823) );
  NAND2_X1 U868 ( .A1(G104), .A2(n913), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G140), .A2(n580), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n784), .ZN(n789) );
  NAND2_X1 U872 ( .A1(G116), .A2(n910), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G128), .A2(n892), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U875 ( .A(KEYINPUT35), .B(n787), .Z(n788) );
  NOR2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U877 ( .A(KEYINPUT36), .B(n790), .ZN(n904) );
  XNOR2_X1 U878 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NOR2_X1 U879 ( .A1(n904), .A2(n811), .ZN(n1019) );
  NAND2_X1 U880 ( .A1(n823), .A2(n1019), .ZN(n819) );
  INV_X1 U881 ( .A(n823), .ZN(n809) );
  NAND2_X1 U882 ( .A1(G107), .A2(n910), .ZN(n792) );
  NAND2_X1 U883 ( .A1(G95), .A2(n913), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G119), .A2(n892), .ZN(n794) );
  NAND2_X1 U886 ( .A1(G131), .A2(n580), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n901) );
  NAND2_X1 U889 ( .A1(G1991), .A2(n901), .ZN(n807) );
  NAND2_X1 U890 ( .A1(G117), .A2(n910), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G129), .A2(n892), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n803) );
  XOR2_X1 U893 ( .A(KEYINPUT38), .B(KEYINPUT87), .Z(n800) );
  NAND2_X1 U894 ( .A1(G105), .A2(n913), .ZN(n799) );
  XNOR2_X1 U895 ( .A(n800), .B(n799), .ZN(n801) );
  XOR2_X1 U896 ( .A(KEYINPUT86), .B(n801), .Z(n802) );
  NOR2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n580), .A2(G141), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n906) );
  NAND2_X1 U900 ( .A1(G1996), .A2(n906), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U902 ( .A(KEYINPUT88), .B(n808), .Z(n1017) );
  NOR2_X1 U903 ( .A1(n809), .A2(n1017), .ZN(n814) );
  INV_X1 U904 ( .A(n814), .ZN(n810) );
  AND2_X1 U905 ( .A1(n819), .A2(n810), .ZN(n842) );
  AND2_X1 U906 ( .A1(n980), .A2(n842), .ZN(n825) );
  NAND2_X1 U907 ( .A1(n904), .A2(n811), .ZN(n1018) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n906), .ZN(n1026) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n901), .ZN(n1014) );
  NOR2_X1 U911 ( .A1(n812), .A2(n1014), .ZN(n813) );
  NOR2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U913 ( .A(KEYINPUT101), .B(n815), .Z(n816) );
  NOR2_X1 U914 ( .A1(n1026), .A2(n816), .ZN(n817) );
  XNOR2_X1 U915 ( .A(KEYINPUT102), .B(n817), .ZN(n818) );
  XNOR2_X1 U916 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n1018), .A2(n821), .ZN(n822) );
  AND2_X1 U919 ( .A1(n822), .A2(n823), .ZN(n843) );
  XNOR2_X1 U920 ( .A(G1986), .B(G290), .ZN(n1000) );
  NAND2_X1 U921 ( .A1(n1000), .A2(n823), .ZN(n824) );
  OR2_X1 U922 ( .A1(n843), .A2(n824), .ZN(n828) );
  AND2_X1 U923 ( .A1(n825), .A2(n828), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n848) );
  INV_X1 U925 ( .A(n828), .ZN(n846) );
  NAND2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n833) );
  NOR2_X1 U927 ( .A1(G2090), .A2(G303), .ZN(n831) );
  NAND2_X1 U928 ( .A1(G8), .A2(n831), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n834), .A2(n838), .ZN(n840) );
  NOR2_X1 U931 ( .A1(G1981), .A2(G305), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n835), .B(KEYINPUT24), .ZN(n836) );
  XNOR2_X1 U933 ( .A(KEYINPUT89), .B(n836), .ZN(n837) );
  OR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n841) );
  AND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(n844) );
  NOR2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n845) );
  OR2_X1 U938 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U939 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U940 ( .A(n849), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U941 ( .A1(G2106), .A2(n850), .ZN(G217) );
  NAND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n852) );
  INV_X1 U943 ( .A(G661), .ZN(n851) );
  NOR2_X1 U944 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U945 ( .A(n853), .B(KEYINPUT103), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U947 ( .A1(n855), .A2(n854), .ZN(G188) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  INV_X1 U951 ( .A(G69), .ZN(G235) );
  NOR2_X1 U952 ( .A1(n857), .A2(n856), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U954 ( .A(n987), .B(G286), .ZN(n859) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n860), .B(G171), .ZN(n861) );
  NOR2_X1 U957 ( .A1(G37), .A2(n861), .ZN(G397) );
  XOR2_X1 U958 ( .A(G2100), .B(G2096), .Z(n863) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(G2678), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(G2090), .Z(n865) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U964 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U965 ( .A(G2084), .B(G2078), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(G227) );
  XOR2_X1 U967 ( .A(KEYINPUT41), .B(KEYINPUT105), .Z(n871) );
  XNOR2_X1 U968 ( .A(KEYINPUT104), .B(G2474), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U970 ( .A(n872), .B(KEYINPUT107), .Z(n874) );
  XNOR2_X1 U971 ( .A(G1971), .B(G1976), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n882) );
  XOR2_X1 U973 ( .A(G1981), .B(G1956), .Z(n876) );
  XNOR2_X1 U974 ( .A(G1986), .B(G1966), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n880) );
  XOR2_X1 U976 ( .A(KEYINPUT106), .B(G1961), .Z(n878) );
  XNOR2_X1 U977 ( .A(G1996), .B(G1991), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(n880), .B(n879), .Z(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(G229) );
  NAND2_X1 U981 ( .A1(n892), .A2(G124), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n883), .B(KEYINPUT44), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G136), .A2(n580), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(KEYINPUT108), .B(n886), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G112), .A2(n910), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G100), .A2(n913), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U989 ( .A1(n890), .A2(n889), .ZN(G162) );
  XNOR2_X1 U990 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n903) );
  NAND2_X1 U991 ( .A1(n580), .A2(G139), .ZN(n891) );
  XNOR2_X1 U992 ( .A(KEYINPUT109), .B(n891), .ZN(n900) );
  NAND2_X1 U993 ( .A1(G115), .A2(n910), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G127), .A2(n892), .ZN(n893) );
  NAND2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n895), .B(KEYINPUT47), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n896), .B(KEYINPUT110), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n913), .A2(G103), .ZN(n897) );
  NAND2_X1 U999 ( .A1(n898), .A2(n897), .ZN(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n1021) );
  XNOR2_X1 U1001 ( .A(n901), .B(n1021), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(G164), .B(G162), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n922) );
  NAND2_X1 U1007 ( .A1(G118), .A2(n910), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(G130), .A2(n892), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n918) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n913), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(G142), .A2(n580), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1013 ( .A(n916), .B(KEYINPUT45), .Z(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n919), .B(n1011), .ZN(n920) );
  XOR2_X1 U1016 ( .A(G160), .B(n920), .Z(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n923), .ZN(G395) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n931), .ZN(n928) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n924) );
  XOR2_X1 U1021 ( .A(KEYINPUT49), .B(n924), .Z(n925) );
  XNOR2_X1 U1022 ( .A(n925), .B(KEYINPUT111), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G397), .A2(n926), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(n929), .A2(G395), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(n930), .B(KEYINPUT112), .ZN(G308) );
  INV_X1 U1027 ( .A(G308), .ZN(G225) );
  INV_X1 U1028 ( .A(n931), .ZN(G319) );
  INV_X1 U1029 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1030 ( .A(KEYINPUT125), .B(G1966), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(G21), .ZN(n951) );
  XOR2_X1 U1032 ( .A(G4), .B(KEYINPUT124), .Z(n934) );
  XNOR2_X1 U1033 ( .A(G1348), .B(KEYINPUT59), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(n934), .B(n933), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(G19), .B(n935), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G1956), .B(G20), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(G6), .B(G1981), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT60), .B(n942), .Z(n949) );
  XNOR2_X1 U1042 ( .A(G1971), .B(G22), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(G23), .B(G1976), .ZN(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n946) );
  XOR2_X1 U1045 ( .A(G1986), .B(G24), .Z(n945) );
  NAND2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(KEYINPUT58), .B(n947), .ZN(n948) );
  NOR2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1050 ( .A(KEYINPUT123), .B(G1961), .Z(n952) );
  XNOR2_X1 U1051 ( .A(G5), .B(n952), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1053 ( .A(n955), .B(KEYINPUT61), .Z(n956) );
  XNOR2_X1 U1054 ( .A(KEYINPUT126), .B(n956), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(G16), .A2(n957), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(n958), .B(KEYINPUT127), .ZN(n979) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(G1996), .B(G32), .ZN(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n965) );
  XOR2_X1 U1060 ( .A(n961), .B(G27), .Z(n963) );
  XNOR2_X1 U1061 ( .A(G33), .B(G2072), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(KEYINPUT117), .B(n966), .ZN(n967) );
  NAND2_X1 U1065 ( .A1(n967), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G25), .B(G1991), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(KEYINPUT116), .B(n968), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n972) );
  XOR2_X1 U1069 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n971) );
  XOR2_X1 U1070 ( .A(n972), .B(n971), .Z(n974) );
  XNOR2_X1 U1071 ( .A(G2090), .B(G35), .ZN(n973) );
  NOR2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1073 ( .A(G2084), .B(KEYINPUT54), .Z(n975) );
  XNOR2_X1 U1074 ( .A(G34), .B(n975), .ZN(n976) );
  NAND2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n1042) );
  INV_X1 U1076 ( .A(KEYINPUT55), .ZN(n1036) );
  OR2_X1 U1077 ( .A1(n1042), .A2(n1036), .ZN(n978) );
  NAND2_X1 U1078 ( .A1(n979), .A2(n978), .ZN(n1009) );
  XOR2_X1 U1079 ( .A(KEYINPUT56), .B(G16), .Z(n1007) );
  XNOR2_X1 U1080 ( .A(G171), .B(G1961), .ZN(n984) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1082 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1083 ( .A(n982), .B(KEYINPUT57), .ZN(n983) );
  NAND2_X1 U1084 ( .A1(n984), .A2(n983), .ZN(n1005) );
  XNOR2_X1 U1085 ( .A(G1341), .B(KEYINPUT122), .ZN(n986) );
  XNOR2_X1 U1086 ( .A(n986), .B(n985), .ZN(n989) );
  XOR2_X1 U1087 ( .A(G1348), .B(n987), .Z(n988) );
  NOR2_X1 U1088 ( .A1(n989), .A2(n988), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(KEYINPUT119), .B(n990), .ZN(n992) );
  NAND2_X1 U1090 ( .A1(n992), .A2(n991), .ZN(n994) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G303), .ZN(n993) );
  NOR2_X1 U1092 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1093 ( .A(KEYINPUT120), .B(n995), .ZN(n998) );
  XNOR2_X1 U1094 ( .A(n996), .B(G1956), .ZN(n997) );
  NAND2_X1 U1095 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1096 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1097 ( .A(KEYINPUT121), .B(n1001), .Z(n1002) );
  NAND2_X1 U1098 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1040) );
  XOR2_X1 U1102 ( .A(G160), .B(G2084), .Z(n1010) );
  XNOR2_X1 U1103 ( .A(KEYINPUT113), .B(n1010), .ZN(n1012) );
  NAND2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(n1015), .B(KEYINPUT114), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1034) );
  INV_X1 U1108 ( .A(n1018), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1032) );
  XOR2_X1 U1110 ( .A(G2072), .B(n1021), .Z(n1023) );
  XOR2_X1 U1111 ( .A(G164), .B(G2078), .Z(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1113 ( .A(KEYINPUT50), .B(n1024), .Z(n1030) );
  XOR2_X1 U1114 ( .A(G2090), .B(G162), .Z(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1116 ( .A(KEYINPUT115), .B(n1027), .Z(n1028) );
  XNOR2_X1 U1117 ( .A(KEYINPUT51), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1121 ( .A(KEYINPUT52), .B(n1035), .ZN(n1037) );
  NAND2_X1 U1122 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(G29), .ZN(n1039) );
  NAND2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1045) );
  NOR2_X1 U1125 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1041) );
  NAND2_X1 U1126 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NAND2_X1 U1127 ( .A1(G11), .A2(n1043), .ZN(n1044) );
  NOR2_X1 U1128 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  XNOR2_X1 U1129 ( .A(n1046), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

