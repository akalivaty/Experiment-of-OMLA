//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT28), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT27), .B(G183gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n206), .B(new_n207), .C1(new_n205), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT27), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n204), .A2(new_n213), .A3(new_n207), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n211), .B1(new_n214), .B2(KEYINPUT28), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT69), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n221), .A2(new_n216), .A3(new_n217), .A4(KEYINPUT69), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n209), .A2(new_n215), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT70), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n209), .A2(new_n215), .A3(new_n226), .A4(new_n223), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT71), .ZN(new_n229));
  INV_X1    g028(.A(G127gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G134gat), .ZN(new_n231));
  INV_X1    g030(.A(G134gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G127gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT71), .B1(new_n230), .B2(G134gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT72), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n235), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n237), .B(new_n238), .C1(new_n239), .C2(new_n229), .ZN(new_n240));
  NAND2_X1  g039(.A1(G113gat), .A2(G120gat), .ZN(new_n241));
  INV_X1    g040(.A(G113gat), .ZN(new_n242));
  INV_X1    g041(.A(G120gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT1), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n236), .A2(new_n240), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT73), .B(G113gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(new_n243), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n247), .A2(new_n239), .A3(new_n244), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT23), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n220), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n250), .B(new_n220), .C1(KEYINPUT66), .C2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT24), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n210), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n212), .A2(new_n207), .ZN(new_n261));
  OAI211_X1 g060(.A(G183gat), .B(G190gat), .C1(KEYINPUT67), .C2(KEYINPUT24), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n253), .A2(new_n255), .A3(new_n257), .A4(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n250), .A2(new_n255), .A3(new_n220), .ZN(new_n265));
  NAND3_X1  g064(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(new_n212), .A3(new_n207), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n270), .A2(new_n271), .B1(new_n259), .B2(new_n210), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n265), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n264), .B1(new_n273), .B2(KEYINPUT25), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n228), .A2(new_n249), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT74), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n228), .A2(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(new_n249), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n265), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n270), .A2(new_n271), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n210), .A2(new_n259), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n266), .B(KEYINPUT64), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n256), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n225), .A2(new_n227), .B1(new_n286), .B2(new_n264), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(new_n288), .A3(new_n249), .ZN(new_n289));
  NAND2_X1  g088(.A1(G227gat), .A2(G233gat), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n276), .A2(new_n279), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n291), .A2(KEYINPUT34), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(KEYINPUT34), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT32), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n279), .A3(new_n289), .ZN(new_n296));
  INV_X1    g095(.A(new_n290), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT33), .B1(new_n296), .B2(new_n297), .ZN(new_n299));
  XNOR2_X1  g098(.A(G15gat), .B(G43gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G71gat), .ZN(new_n301));
  INV_X1    g100(.A(G99gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n298), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  AOI221_X4 g104(.A(new_n295), .B1(KEYINPUT33), .B2(new_n303), .C1(new_n296), .C2(new_n297), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n294), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n296), .A2(new_n297), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT33), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n304), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n298), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n306), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n291), .A2(KEYINPUT34), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n291), .A2(KEYINPUT34), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT36), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT77), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n314), .B2(new_n315), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n292), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(new_n326), .C1(new_n305), .C2(new_n306), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT36), .A3(new_n317), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n327), .A2(KEYINPUT76), .A3(KEYINPUT36), .A4(new_n317), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n321), .A2(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n274), .A2(new_n224), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(new_n333), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT78), .B(G218gat), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT22), .B1(new_n338), .B2(G211gat), .ZN(new_n339));
  XOR2_X1   g138(.A(G197gat), .B(G204gat), .Z(new_n340));
  OAI21_X1  g139(.A(G211gat), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G218gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT78), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G218gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(G211gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT22), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n340), .ZN(new_n349));
  INV_X1    g148(.A(G211gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n341), .A2(G218gat), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(G218gat), .B1(new_n341), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n274), .A2(new_n224), .ZN(new_n355));
  INV_X1    g154(.A(new_n333), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT79), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n334), .A2(new_n337), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT80), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n277), .A2(new_n356), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n333), .B1(new_n336), .B2(KEYINPUT29), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n361), .B1(new_n364), .B2(KEYINPUT80), .ZN(new_n365));
  OAI211_X1 g164(.A(KEYINPUT37), .B(new_n358), .C1(new_n365), .C2(new_n354), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT37), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n333), .B1(new_n228), .B2(new_n274), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT80), .B1(new_n368), .B2(new_n360), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n354), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n358), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(G64gat), .ZN(new_n376));
  INV_X1    g175(.A(G92gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n366), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n372), .B2(new_n373), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(KEYINPUT81), .B(new_n380), .C1(new_n372), .C2(new_n373), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n379), .A2(KEYINPUT38), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G57gat), .B(G85gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G141gat), .B(G148gat), .Z(new_n394));
  INV_X1    g193(.A(KEYINPUT2), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n395), .B2(new_n398), .ZN(new_n401));
  XNOR2_X1  g200(.A(G141gat), .B(G148gat), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n401), .A2(KEYINPUT82), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n395), .ZN(new_n405));
  NAND2_X1  g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n407), .B2(new_n394), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n400), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n409), .A2(new_n245), .A3(new_n248), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT82), .B1(new_n401), .B2(new_n402), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n394), .A3(new_n404), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n411), .A2(new_n412), .B1(new_n396), .B2(new_n399), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n236), .A2(new_n240), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n244), .A2(new_n241), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n247), .A2(new_n239), .A3(new_n244), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n393), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT5), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n417), .A3(new_n413), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(KEYINPUT4), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(KEYINPUT4), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n249), .A2(KEYINPUT84), .A3(new_n425), .A4(new_n413), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n412), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(new_n400), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n430), .B1(new_n413), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n393), .B1(new_n432), .B2(new_n278), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n420), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n430), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n400), .A3(new_n431), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n278), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n393), .A2(KEYINPUT5), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n249), .A2(new_n425), .A3(new_n413), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n425), .B1(new_n249), .B2(new_n413), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n437), .B(new_n438), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n391), .B1(new_n434), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n427), .A2(new_n433), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n390), .B(new_n442), .C1(new_n445), .C2(new_n420), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(KEYINPUT6), .B(new_n391), .C1(new_n434), .C2(new_n443), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n365), .A2(new_n354), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n334), .A2(new_n337), .A3(new_n357), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n451), .B(KEYINPUT37), .C1(new_n354), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT38), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n378), .A4(new_n374), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n385), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n410), .A2(new_n418), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(new_n393), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT90), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(new_n393), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n459), .B(KEYINPUT39), .C1(new_n462), .C2(new_n458), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n424), .A2(new_n439), .B1(new_n432), .B2(new_n278), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n392), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n391), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(KEYINPUT91), .A2(KEYINPUT40), .ZN(new_n468));
  NOR2_X1   g267(.A1(KEYINPUT91), .A2(KEYINPUT40), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n461), .A2(new_n393), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n390), .B1(new_n472), .B2(KEYINPUT39), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT90), .B1(new_n464), .B2(new_n392), .ZN(new_n474));
  INV_X1    g273(.A(new_n458), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n473), .B1(new_n476), .B2(new_n459), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n444), .A2(new_n468), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT30), .B1(new_n383), .B2(new_n384), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT30), .B(new_n380), .C1(new_n372), .C2(new_n373), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n358), .B(new_n378), .C1(new_n365), .C2(new_n354), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n479), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n409), .A2(new_n359), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n352), .B2(new_n353), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n339), .A2(G211gat), .A3(new_n340), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n350), .B1(new_n348), .B2(new_n349), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n342), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n341), .A2(G218gat), .A3(new_n351), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n490), .A2(new_n359), .A3(new_n436), .A4(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n431), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n487), .A2(new_n492), .B1(new_n409), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n485), .B1(new_n494), .B2(KEYINPUT86), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n487), .A2(new_n492), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n435), .ZN(new_n497));
  INV_X1    g296(.A(new_n485), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n409), .A2(new_n493), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n495), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G22gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n495), .B(G22gat), .C1(new_n499), .C2(new_n502), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT87), .A3(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(KEYINPUT87), .ZN(new_n508));
  XOR2_X1   g307(.A(G78gat), .B(G106gat), .Z(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT31), .ZN(new_n510));
  INV_X1    g309(.A(G50gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n503), .A2(new_n515), .A3(new_n504), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n503), .B2(new_n504), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n506), .B(KEYINPUT88), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n456), .A2(new_n484), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n505), .A2(KEYINPUT89), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n515), .A3(new_n504), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n506), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(new_n503), .B2(new_n504), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n512), .B1(new_n528), .B2(new_n506), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n524), .A2(new_n526), .B1(new_n529), .B2(new_n508), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n383), .A2(new_n384), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n483), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n448), .A2(new_n449), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n332), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n305), .A2(new_n306), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n325), .A2(new_n326), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n317), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n523), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(new_n526), .A3(new_n512), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n514), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n450), .A2(new_n480), .A3(new_n483), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n530), .A2(new_n318), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n480), .A2(new_n483), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n535), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n547), .A2(KEYINPUT35), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n202), .B1(new_n539), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n521), .A2(new_n537), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n328), .A2(new_n329), .ZN(new_n557));
  INV_X1    g356(.A(new_n331), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n322), .B1(new_n318), .B2(new_n319), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT77), .B(KEYINPUT36), .C1(new_n307), .C2(new_n317), .ZN(new_n560));
  OAI22_X1  g359(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n318), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n546), .A2(new_n520), .A3(new_n563), .A4(new_n551), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n530), .A2(new_n536), .A3(new_n542), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(KEYINPUT93), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n555), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G8gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT94), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(G1gat), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n570), .B1(new_n574), .B2(KEYINPUT95), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n572), .A2(G1gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n576), .B(new_n574), .C1(KEYINPUT95), .C2(new_n570), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G43gat), .B(G50gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(G29gat), .A2(G36gat), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n583), .A2(KEYINPUT14), .ZN(new_n584));
  INV_X1    g383(.A(new_n583), .ZN(new_n585));
  INV_X1    g384(.A(G29gat), .ZN(new_n586));
  INV_X1    g385(.A(G36gat), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT14), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n584), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n589), .A2(KEYINPUT15), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(KEYINPUT15), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n582), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(KEYINPUT15), .ZN(new_n593));
  INV_X1    g392(.A(new_n582), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT17), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n592), .A2(new_n595), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT17), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n580), .A2(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT96), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n580), .B(new_n598), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n604), .B(KEYINPUT97), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT13), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n601), .A2(KEYINPUT18), .A3(new_n602), .A4(new_n605), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G113gat), .B(G141gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G197gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT11), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n216), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n608), .A2(new_n621), .A3(new_n612), .A4(new_n613), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G57gat), .B(G64gat), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G71gat), .B(G78gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT21), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n581), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G127gat), .B(G155gat), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n580), .A2(new_n631), .A3(new_n630), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n633), .B2(new_n636), .ZN(new_n639));
  OAI211_X1 g438(.A(G231gat), .B(G233gat), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n633), .A2(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n634), .ZN(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n637), .ZN(new_n644));
  XOR2_X1   g443(.A(G183gat), .B(G211gat), .Z(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT99), .B(KEYINPUT20), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n640), .A2(new_n644), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n640), .B2(new_n644), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G85gat), .A2(G92gat), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT7), .B1(new_n653), .B2(KEYINPUT100), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(KEYINPUT100), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(G106gat), .ZN(new_n657));
  OR3_X1    g456(.A1(new_n302), .A2(new_n657), .A3(KEYINPUT101), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT101), .B1(new_n302), .B2(new_n657), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(KEYINPUT8), .A3(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n656), .B(new_n660), .C1(G85gat), .C2(G92gat), .ZN(new_n661));
  XOR2_X1   g460(.A(G99gat), .B(G106gat), .Z(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n600), .A2(new_n597), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n665), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n663), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n598), .ZN(new_n670));
  NAND3_X1  g469(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G190gat), .B(G218gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n667), .A2(new_n670), .A3(new_n673), .A4(new_n671), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT103), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n675), .A2(new_n676), .A3(new_n680), .A4(new_n677), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G134gat), .ZN(new_n684));
  INV_X1    g483(.A(G162gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n675), .A2(new_n677), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(KEYINPUT102), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n679), .A3(new_n681), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n652), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT104), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n217), .ZN(new_n697));
  INV_X1    g496(.A(G204gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n630), .B1(new_n668), .B2(new_n663), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n664), .A2(new_n628), .A3(new_n665), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT10), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n669), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(G230gat), .A2(G233gat), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n705), .A2(KEYINPUT105), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT105), .B1(new_n705), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n701), .ZN(new_n710));
  INV_X1    g509(.A(new_n706), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n699), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n705), .A2(new_n706), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n712), .A3(new_n699), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n694), .A2(KEYINPUT106), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n650), .A2(new_n651), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n719), .A2(new_n717), .A3(new_n692), .A4(new_n691), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n569), .A2(new_n623), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n535), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g525(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n573), .A2(new_n570), .ZN(new_n728));
  NOR4_X1   g527(.A1(new_n724), .A2(new_n549), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n724), .A2(new_n549), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n729), .A2(KEYINPUT42), .B1(new_n730), .B2(G8gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n724), .A2(new_n549), .ZN(new_n732));
  INV_X1    g531(.A(new_n727), .ZN(new_n733));
  INV_X1    g532(.A(new_n728), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT107), .B1(new_n729), .B2(KEYINPUT42), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n731), .A2(new_n738), .A3(new_n739), .ZN(G1325gat));
  INV_X1    g539(.A(G15gat), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n724), .A2(new_n741), .A3(new_n561), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n724), .B2(new_n318), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(G1326gat));
  NOR2_X1   g546(.A1(new_n724), .A2(new_n520), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT43), .B(G22gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1327gat));
  AOI21_X1  g549(.A(new_n566), .B1(new_n545), .B2(new_n546), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n520), .A2(new_n563), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n552), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT109), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n755), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n562), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n693), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n555), .A2(new_n568), .A3(KEYINPUT44), .A4(new_n693), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n717), .ZN(new_n763));
  INV_X1    g562(.A(new_n623), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n719), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n762), .A2(new_n450), .A3(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n555), .A2(new_n568), .A3(new_n693), .A4(new_n765), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n586), .A3(new_n450), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(KEYINPUT45), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(KEYINPUT45), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n766), .A2(new_n586), .B1(new_n770), .B2(new_n771), .ZN(G1328gat));
  INV_X1    g571(.A(new_n549), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n768), .A2(new_n587), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n762), .A2(new_n773), .A3(new_n765), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n587), .ZN(G1329gat));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n332), .A3(new_n761), .A4(new_n765), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G43gat), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n767), .A2(G43gat), .A3(new_n318), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1330gat));
  INV_X1    g583(.A(KEYINPUT48), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n768), .A2(KEYINPUT111), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n520), .B1(new_n767), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n511), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n760), .A2(new_n530), .A3(new_n761), .A4(new_n765), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G50gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n785), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n785), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n767), .A2(new_n787), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n530), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n511), .B1(new_n767), .B2(new_n787), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n786), .A2(new_n788), .A3(new_n793), .A4(new_n511), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n790), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT110), .B1(new_n790), .B2(G50gat), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n792), .B1(new_n800), .B2(new_n803), .ZN(G1331gat));
  AND2_X1   g603(.A1(new_n757), .A2(new_n764), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n652), .A2(new_n693), .A3(new_n717), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n450), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n549), .ZN(new_n811));
  NOR2_X1   g610(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n812));
  AND2_X1   g611(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n811), .B2(new_n812), .ZN(G1333gat));
  NOR2_X1   g614(.A1(new_n807), .A2(new_n318), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n332), .A2(G71gat), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n816), .A2(G71gat), .B1(new_n807), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g618(.A1(new_n808), .A2(new_n530), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g620(.A1(new_n719), .A2(new_n623), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n760), .A2(new_n763), .A3(new_n761), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G85gat), .B1(new_n823), .B2(new_n535), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n757), .A2(new_n693), .A3(new_n822), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n757), .A2(KEYINPUT51), .A3(new_n693), .A4(new_n822), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n717), .A2(G85gat), .A3(new_n535), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT113), .Z(new_n832));
  OAI21_X1  g631(.A(new_n824), .B1(new_n830), .B2(new_n832), .ZN(G1336gat));
  OAI21_X1  g632(.A(G92gat), .B1(new_n823), .B2(new_n549), .ZN(new_n834));
  XNOR2_X1  g633(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n829), .A2(new_n377), .A3(new_n773), .A4(new_n763), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n834), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(G1337gat));
  OAI21_X1  g638(.A(G99gat), .B1(new_n823), .B2(new_n561), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n829), .A2(new_n302), .A3(new_n563), .A4(new_n763), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1338gat));
  OAI21_X1  g641(.A(G106gat), .B1(new_n823), .B2(new_n520), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n829), .A2(new_n657), .A3(new_n530), .A4(new_n763), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n847), .A3(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1339gat));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n707), .B2(new_n708), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n703), .A2(new_n711), .A3(new_n704), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n714), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n699), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n851), .A2(new_n853), .A3(KEYINPUT55), .A4(new_n854), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n857), .A2(new_n623), .A3(new_n715), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n609), .A2(new_n611), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n605), .B1(new_n601), .B2(new_n602), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n618), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n622), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n713), .B2(new_n716), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n693), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n689), .A2(new_n679), .A3(new_n681), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n688), .A2(KEYINPUT102), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n679), .A2(new_n681), .B1(new_n867), .B2(new_n686), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n857), .A2(new_n715), .A3(new_n858), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n652), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n694), .A2(new_n764), .A3(new_n717), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n773), .A2(new_n535), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n530), .A3(new_n542), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n246), .A3(new_n623), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n876), .A2(new_n752), .A3(new_n764), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n242), .ZN(G1340gat));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n243), .A3(new_n763), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n876), .A2(new_n752), .A3(new_n717), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n243), .ZN(G1341gat));
  AOI21_X1  g682(.A(G127gat), .B1(new_n877), .B2(new_n719), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n876), .A2(new_n752), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n652), .A2(new_n230), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(G1342gat));
  NAND3_X1  g686(.A1(new_n877), .A2(new_n232), .A3(new_n693), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n888), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT115), .B1(new_n888), .B2(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n892));
  INV_X1    g691(.A(new_n693), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n548), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G134gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n891), .A2(new_n892), .A3(new_n896), .ZN(G1343gat));
  NAND2_X1  g696(.A1(new_n874), .A2(new_n530), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n561), .A2(new_n875), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(G141gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n623), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  XOR2_X1   g702(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n904));
  NAND2_X1  g703(.A1(new_n855), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n905), .A2(new_n623), .A3(new_n715), .A4(new_n858), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n693), .B1(new_n906), .B2(new_n864), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n652), .B1(new_n907), .B2(new_n871), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT117), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n910), .B(new_n652), .C1(new_n907), .C2(new_n871), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n873), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n903), .B1(new_n912), .B2(new_n530), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT57), .B(new_n520), .C1(new_n872), .C2(new_n873), .ZN(new_n914));
  NOR4_X1   g713(.A1(new_n913), .A2(new_n764), .A3(new_n899), .A4(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n902), .B1(new_n915), .B2(new_n901), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT58), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n902), .B(new_n918), .C1(new_n915), .C2(new_n901), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(G148gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n900), .A2(new_n921), .A3(new_n763), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n913), .A2(new_n899), .A3(new_n914), .ZN(new_n923));
  AOI211_X1 g722(.A(KEYINPUT59), .B(new_n921), .C1(new_n923), .C2(new_n763), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n623), .B1(new_n718), .B2(new_n722), .ZN(new_n926));
  INV_X1    g725(.A(new_n907), .ZN(new_n927));
  INV_X1    g726(.A(new_n871), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n719), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT118), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n720), .A2(new_n721), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n720), .A2(new_n721), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n764), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n908), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n930), .A2(new_n935), .A3(new_n903), .A4(new_n530), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n898), .A2(KEYINPUT57), .ZN(new_n937));
  INV_X1    g736(.A(new_n899), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n936), .A2(new_n763), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n925), .B1(new_n939), .B2(G148gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n940), .ZN(G1345gat));
  AOI21_X1  g740(.A(G155gat), .B1(new_n900), .B2(new_n719), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n719), .A2(G155gat), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT119), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n923), .B2(new_n944), .ZN(G1346gat));
  NOR2_X1   g744(.A1(new_n332), .A2(new_n520), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n894), .A2(new_n685), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n923), .A2(new_n693), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n685), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n549), .A2(new_n450), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n951), .B1(new_n872), .B2(new_n873), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n545), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT120), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n216), .A3(new_n623), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n950), .B(KEYINPUT121), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n874), .A2(new_n548), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(G169gat), .B1(new_n957), .B2(new_n764), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n955), .A2(new_n958), .ZN(G1348gat));
  NOR3_X1   g758(.A1(new_n957), .A2(new_n217), .A3(new_n717), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n954), .A2(new_n763), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n217), .ZN(G1349gat));
  OR3_X1    g761(.A1(new_n957), .A2(KEYINPUT122), .A3(new_n652), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT122), .B1(new_n957), .B2(new_n652), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(G183gat), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n953), .A2(new_n208), .A3(new_n719), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT60), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT124), .Z(new_n970));
  XNOR2_X1  g769(.A(new_n967), .B(new_n970), .ZN(G1350gat));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n207), .A3(new_n693), .ZN(new_n972));
  OAI21_X1  g771(.A(G190gat), .B1(new_n957), .B2(new_n893), .ZN(new_n973));
  XOR2_X1   g772(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n972), .A2(new_n975), .ZN(G1351gat));
  NAND2_X1  g775(.A1(new_n956), .A2(new_n561), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n936), .A2(new_n937), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n764), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n952), .A2(new_n946), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n764), .A2(G197gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(G1352gat));
  NAND4_X1  g782(.A1(new_n936), .A2(new_n763), .A3(new_n937), .A4(new_n978), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n952), .A2(new_n698), .A3(new_n763), .A4(new_n946), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT62), .Z(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n985), .A2(KEYINPUT127), .A3(new_n987), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1353gat));
  NAND4_X1  g791(.A1(new_n936), .A2(new_n719), .A3(new_n937), .A4(new_n978), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n993), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n994));
  AOI21_X1  g793(.A(KEYINPUT63), .B1(new_n993), .B2(G211gat), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n719), .A2(new_n350), .ZN(new_n996));
  OAI22_X1  g795(.A1(new_n994), .A2(new_n995), .B1(new_n981), .B2(new_n996), .ZN(G1354gat));
  INV_X1    g796(.A(new_n338), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n979), .A2(new_n998), .A3(new_n893), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n952), .A2(new_n693), .A3(new_n946), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n999), .B1(new_n342), .B2(new_n1000), .ZN(G1355gat));
endmodule


