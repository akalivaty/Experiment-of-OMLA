

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X4 U555 ( .A1(G651), .A2(G543), .ZN(n587) );
  INV_X1 U556 ( .A(KEYINPUT93), .ZN(n709) );
  AND2_X1 U557 ( .A1(n775), .A2(n755), .ZN(n759) );
  XNOR2_X1 U558 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U559 ( .A1(G8), .A2(n728), .ZN(n780) );
  INV_X1 U560 ( .A(KEYINPUT70), .ZN(n599) );
  NOR2_X2 U561 ( .A1(n660), .A2(n525), .ZN(n590) );
  OR2_X1 U562 ( .A1(n759), .A2(n758), .ZN(n519) );
  AND2_X1 U563 ( .A1(n829), .A2(n986), .ZN(n520) );
  INV_X1 U564 ( .A(KEYINPUT27), .ZN(n692) );
  XNOR2_X1 U565 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U566 ( .A1(n703), .A2(n702), .ZN(n711) );
  NOR2_X1 U567 ( .A1(n752), .A2(n749), .ZN(n729) );
  XNOR2_X1 U568 ( .A(n730), .B(KEYINPUT30), .ZN(n731) );
  XNOR2_X1 U569 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n734) );
  INV_X1 U570 ( .A(KEYINPUT95), .ZN(n738) );
  OR2_X1 U571 ( .A1(n737), .A2(n736), .ZN(n750) );
  INV_X1 U572 ( .A(n780), .ZN(n760) );
  INV_X1 U573 ( .A(n992), .ZN(n765) );
  XNOR2_X1 U574 ( .A(n588), .B(KEYINPUT12), .ZN(n589) );
  AND2_X1 U575 ( .A1(n691), .A2(n796), .ZN(n721) );
  NAND2_X1 U576 ( .A1(n659), .A2(G56), .ZN(n586) );
  NOR2_X1 U577 ( .A1(n798), .A2(n520), .ZN(n815) );
  AND2_X1 U578 ( .A1(n815), .A2(n818), .ZN(n816) );
  INV_X1 U579 ( .A(KEYINPUT1), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n817), .A2(n816), .ZN(n832) );
  NOR2_X1 U581 ( .A1(G651), .A2(n660), .ZN(n655) );
  XNOR2_X1 U582 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n536) );
  XNOR2_X1 U583 ( .A(n537), .B(n536), .ZN(n546) );
  AND2_X1 U584 ( .A1(n546), .A2(n545), .ZN(G160) );
  NAND2_X1 U585 ( .A1(n587), .A2(G89), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(KEYINPUT4), .ZN(n523) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n660) );
  NAND2_X1 U588 ( .A1(G76), .A2(n590), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT5), .ZN(n533) );
  XNOR2_X1 U591 ( .A(KEYINPUT6), .B(KEYINPUT73), .ZN(n531) );
  INV_X1 U592 ( .A(G651), .ZN(n525) );
  NOR2_X1 U593 ( .A1(n525), .A2(G543), .ZN(n527) );
  XNOR2_X2 U594 ( .A(n527), .B(n526), .ZN(n659) );
  NAND2_X1 U595 ( .A1(G63), .A2(n659), .ZN(n529) );
  NAND2_X1 U596 ( .A1(G51), .A2(n655), .ZN(n528) );
  NAND2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(KEYINPUT7), .B(n534), .ZN(G168) );
  INV_X1 U601 ( .A(G2104), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n539), .A2(G2105), .ZN(n535) );
  XNOR2_X2 U603 ( .A(n535), .B(KEYINPUT64), .ZN(n902) );
  NAND2_X1 U604 ( .A1(n902), .A2(G101), .ZN(n537) );
  NOR2_X1 U605 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  XOR2_X1 U606 ( .A(KEYINPUT17), .B(n538), .Z(n622) );
  NAND2_X1 U607 ( .A1(G137), .A2(n622), .ZN(n544) );
  AND2_X1 U608 ( .A1(n539), .A2(G2105), .ZN(n898) );
  NAND2_X1 U609 ( .A1(n898), .A2(G125), .ZN(n542) );
  NAND2_X1 U610 ( .A1(G2105), .A2(G2104), .ZN(n540) );
  XOR2_X1 U611 ( .A(KEYINPUT66), .B(n540), .Z(n551) );
  NAND2_X1 U612 ( .A1(G113), .A2(n551), .ZN(n541) );
  AND2_X1 U613 ( .A1(n542), .A2(n541), .ZN(n543) );
  AND2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U615 ( .A1(G102), .A2(n902), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n622), .A2(G138), .ZN(n547) );
  NAND2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n550) );
  INV_X1 U618 ( .A(KEYINPUT83), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n898), .A2(G126), .ZN(n553) );
  BUF_X1 U621 ( .A(n551), .Z(n899) );
  NAND2_X1 U622 ( .A1(G114), .A2(n899), .ZN(n552) );
  NAND2_X1 U623 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U624 ( .A1(n555), .A2(n554), .ZN(G164) );
  NAND2_X1 U625 ( .A1(G85), .A2(n587), .ZN(n557) );
  NAND2_X1 U626 ( .A1(G60), .A2(n659), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U628 ( .A1(G72), .A2(n590), .ZN(n559) );
  NAND2_X1 U629 ( .A1(G47), .A2(n655), .ZN(n558) );
  NAND2_X1 U630 ( .A1(n559), .A2(n558), .ZN(n560) );
  OR2_X1 U631 ( .A1(n561), .A2(n560), .ZN(G290) );
  XOR2_X1 U632 ( .A(G2443), .B(G2446), .Z(n563) );
  XNOR2_X1 U633 ( .A(G2427), .B(G2451), .ZN(n562) );
  XNOR2_X1 U634 ( .A(n563), .B(n562), .ZN(n569) );
  XOR2_X1 U635 ( .A(G2430), .B(G2454), .Z(n565) );
  XNOR2_X1 U636 ( .A(G1348), .B(G1341), .ZN(n564) );
  XNOR2_X1 U637 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U638 ( .A(G2435), .B(G2438), .Z(n566) );
  XNOR2_X1 U639 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U640 ( .A(n569), .B(n568), .Z(n570) );
  AND2_X1 U641 ( .A1(G14), .A2(n570), .ZN(G401) );
  NAND2_X1 U642 ( .A1(G64), .A2(n659), .ZN(n572) );
  NAND2_X1 U643 ( .A1(G52), .A2(n655), .ZN(n571) );
  NAND2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G90), .A2(n587), .ZN(n574) );
  NAND2_X1 U646 ( .A1(G77), .A2(n590), .ZN(n573) );
  NAND2_X1 U647 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U648 ( .A(KEYINPUT9), .B(n575), .Z(n576) );
  NOR2_X1 U649 ( .A1(n577), .A2(n576), .ZN(G171) );
  AND2_X1 U650 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U651 ( .A1(G65), .A2(n659), .ZN(n579) );
  NAND2_X1 U652 ( .A1(G53), .A2(n655), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U654 ( .A1(G91), .A2(n587), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G78), .A2(n590), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U657 ( .A1(n583), .A2(n582), .ZN(n715) );
  INV_X1 U658 ( .A(n715), .ZN(G299) );
  NAND2_X1 U659 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U660 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U661 ( .A(G223), .ZN(n835) );
  NAND2_X1 U662 ( .A1(n835), .A2(G567), .ZN(n585) );
  XOR2_X1 U663 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  XNOR2_X1 U664 ( .A(n586), .B(KEYINPUT14), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G81), .A2(n587), .ZN(n588) );
  XNOR2_X1 U666 ( .A(n589), .B(KEYINPUT68), .ZN(n592) );
  NAND2_X1 U667 ( .A1(G68), .A2(n590), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U669 ( .A(KEYINPUT13), .B(n593), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n596), .B(KEYINPUT69), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G43), .A2(n655), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X2 U674 ( .A(n600), .B(n599), .ZN(n978) );
  NAND2_X1 U675 ( .A1(G860), .A2(n978), .ZN(G153) );
  XNOR2_X1 U676 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U677 ( .A1(G868), .A2(G301), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G92), .A2(n587), .ZN(n602) );
  NAND2_X1 U679 ( .A1(G66), .A2(n659), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U681 ( .A(KEYINPUT72), .B(n603), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G79), .A2(n590), .ZN(n605) );
  NAND2_X1 U683 ( .A1(G54), .A2(n655), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U686 ( .A(KEYINPUT15), .B(n608), .Z(n975) );
  OR2_X1 U687 ( .A1(n975), .A2(G868), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(G284) );
  XOR2_X1 U689 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n612) );
  INV_X1 U691 ( .A(G868), .ZN(n670) );
  NOR2_X1 U692 ( .A1(G286), .A2(n670), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n612), .A2(n611), .ZN(G297) );
  INV_X1 U694 ( .A(G860), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G559), .A2(n613), .ZN(n614) );
  XNOR2_X1 U696 ( .A(KEYINPUT74), .B(n614), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n615), .A2(n975), .ZN(n616) );
  XNOR2_X1 U698 ( .A(KEYINPUT16), .B(n616), .ZN(G148) );
  NOR2_X1 U699 ( .A1(G559), .A2(n670), .ZN(n617) );
  NAND2_X1 U700 ( .A1(n975), .A2(n617), .ZN(n618) );
  XNOR2_X1 U701 ( .A(n618), .B(KEYINPUT75), .ZN(n620) );
  AND2_X1 U702 ( .A1(n978), .A2(n670), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U704 ( .A1(G123), .A2(n898), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT18), .ZN(n625) );
  INV_X1 U706 ( .A(n622), .ZN(n623) );
  INV_X1 U707 ( .A(n623), .ZN(n904) );
  NAND2_X1 U708 ( .A1(n904), .A2(G135), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G99), .A2(n902), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G111), .A2(n899), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n920) );
  XNOR2_X1 U714 ( .A(n920), .B(G2096), .ZN(n631) );
  INV_X1 U715 ( .A(G2100), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(G156) );
  NAND2_X1 U717 ( .A1(G93), .A2(n587), .ZN(n633) );
  NAND2_X1 U718 ( .A1(G80), .A2(n590), .ZN(n632) );
  NAND2_X1 U719 ( .A1(n633), .A2(n632), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G67), .A2(n659), .ZN(n635) );
  NAND2_X1 U721 ( .A1(G55), .A2(n655), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U723 ( .A(KEYINPUT77), .B(n636), .Z(n637) );
  OR2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n671) );
  NAND2_X1 U725 ( .A1(G559), .A2(n975), .ZN(n639) );
  XOR2_X1 U726 ( .A(n978), .B(n639), .Z(n668) );
  XNOR2_X1 U727 ( .A(KEYINPUT76), .B(n668), .ZN(n640) );
  NOR2_X1 U728 ( .A1(G860), .A2(n640), .ZN(n641) );
  XOR2_X1 U729 ( .A(n671), .B(n641), .Z(G145) );
  NAND2_X1 U730 ( .A1(G88), .A2(n587), .ZN(n643) );
  NAND2_X1 U731 ( .A1(G75), .A2(n590), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U733 ( .A1(G62), .A2(n659), .ZN(n645) );
  NAND2_X1 U734 ( .A1(G50), .A2(n655), .ZN(n644) );
  NAND2_X1 U735 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U736 ( .A1(n647), .A2(n646), .ZN(G166) );
  NAND2_X1 U737 ( .A1(G86), .A2(n587), .ZN(n649) );
  NAND2_X1 U738 ( .A1(G61), .A2(n659), .ZN(n648) );
  NAND2_X1 U739 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U740 ( .A1(n590), .A2(G73), .ZN(n650) );
  XOR2_X1 U741 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U742 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U743 ( .A1(n655), .A2(G48), .ZN(n653) );
  NAND2_X1 U744 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U745 ( .A1(G49), .A2(n655), .ZN(n657) );
  NAND2_X1 U746 ( .A1(G74), .A2(G651), .ZN(n656) );
  NAND2_X1 U747 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U748 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U749 ( .A1(n660), .A2(G87), .ZN(n661) );
  NAND2_X1 U750 ( .A1(n662), .A2(n661), .ZN(G288) );
  XNOR2_X1 U751 ( .A(KEYINPUT19), .B(G290), .ZN(n667) );
  XNOR2_X1 U752 ( .A(n671), .B(n715), .ZN(n663) );
  XNOR2_X1 U753 ( .A(n663), .B(G305), .ZN(n664) );
  XNOR2_X1 U754 ( .A(G166), .B(n664), .ZN(n665) );
  XNOR2_X1 U755 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U756 ( .A(n667), .B(n666), .ZN(n843) );
  XOR2_X1 U757 ( .A(n843), .B(n668), .Z(n669) );
  NOR2_X1 U758 ( .A1(n670), .A2(n669), .ZN(n673) );
  NOR2_X1 U759 ( .A1(G868), .A2(n671), .ZN(n672) );
  NOR2_X1 U760 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2084), .A2(G2078), .ZN(n675) );
  XOR2_X1 U762 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n674) );
  XNOR2_X1 U763 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U764 ( .A1(n676), .A2(G2090), .ZN(n677) );
  XOR2_X1 U765 ( .A(KEYINPUT21), .B(n677), .Z(n678) );
  XNOR2_X1 U766 ( .A(KEYINPUT79), .B(n678), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U768 ( .A(KEYINPUT67), .B(G57), .ZN(G237) );
  XNOR2_X1 U769 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U770 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U771 ( .A1(G237), .A2(n680), .ZN(n681) );
  XNOR2_X1 U772 ( .A(KEYINPUT82), .B(n681), .ZN(n682) );
  NAND2_X1 U773 ( .A1(n682), .A2(G108), .ZN(n841) );
  NAND2_X1 U774 ( .A1(n841), .A2(G567), .ZN(n689) );
  XOR2_X1 U775 ( .A(KEYINPUT80), .B(KEYINPUT22), .Z(n684) );
  NAND2_X1 U776 ( .A1(G132), .A2(G82), .ZN(n683) );
  XNOR2_X1 U777 ( .A(n684), .B(n683), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n685), .A2(G96), .ZN(n686) );
  NOR2_X1 U779 ( .A1(n686), .A2(G218), .ZN(n687) );
  XNOR2_X1 U780 ( .A(n687), .B(KEYINPUT81), .ZN(n840) );
  NAND2_X1 U781 ( .A1(n840), .A2(G2106), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n919) );
  NAND2_X1 U783 ( .A1(G661), .A2(G483), .ZN(n690) );
  NOR2_X1 U784 ( .A1(n919), .A2(n690), .ZN(n839) );
  NAND2_X1 U785 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U786 ( .A(G166), .ZN(G303) );
  INV_X1 U787 ( .A(KEYINPUT90), .ZN(n697) );
  AND2_X1 U788 ( .A1(G160), .A2(G40), .ZN(n691) );
  NOR2_X1 U789 ( .A1(G164), .A2(G1384), .ZN(n796) );
  INV_X1 U790 ( .A(n721), .ZN(n740) );
  NAND2_X1 U791 ( .A1(G1956), .A2(n740), .ZN(n695) );
  NAND2_X1 U792 ( .A1(n721), .A2(G2072), .ZN(n693) );
  NAND2_X1 U793 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U794 ( .A(n697), .B(n696), .ZN(n714) );
  NOR2_X1 U795 ( .A1(n715), .A2(n714), .ZN(n698) );
  XOR2_X1 U796 ( .A(n698), .B(KEYINPUT28), .Z(n719) );
  NAND2_X1 U797 ( .A1(n721), .A2(G1996), .ZN(n699) );
  XNOR2_X1 U798 ( .A(n699), .B(KEYINPUT26), .ZN(n700) );
  NAND2_X1 U799 ( .A1(n700), .A2(n978), .ZN(n703) );
  INV_X1 U800 ( .A(n721), .ZN(n728) );
  NAND2_X1 U801 ( .A1(G1341), .A2(n728), .ZN(n701) );
  XNOR2_X1 U802 ( .A(n701), .B(KEYINPUT91), .ZN(n702) );
  NAND2_X1 U803 ( .A1(n711), .A2(n975), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n740), .A2(G1348), .ZN(n705) );
  NAND2_X1 U805 ( .A1(n721), .A2(G2067), .ZN(n704) );
  NAND2_X1 U806 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U807 ( .A(n706), .B(KEYINPUT92), .ZN(n707) );
  NAND2_X1 U808 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U809 ( .A(n710), .B(n709), .ZN(n713) );
  OR2_X1 U810 ( .A1(n975), .A2(n711), .ZN(n712) );
  NAND2_X1 U811 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U813 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U815 ( .A(n720), .B(KEYINPUT29), .ZN(n725) );
  INV_X1 U816 ( .A(G171), .ZN(n727) );
  XOR2_X1 U817 ( .A(G2078), .B(KEYINPUT25), .Z(n955) );
  NOR2_X1 U818 ( .A1(n955), .A2(n740), .ZN(n723) );
  NOR2_X1 U819 ( .A1(n721), .A2(G1961), .ZN(n722) );
  NOR2_X1 U820 ( .A1(n723), .A2(n722), .ZN(n726) );
  NOR2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n724) );
  NOR2_X1 U822 ( .A1(n725), .A2(n724), .ZN(n737) );
  AND2_X1 U823 ( .A1(n727), .A2(n726), .ZN(n733) );
  NOR2_X1 U824 ( .A1(G1966), .A2(n780), .ZN(n752) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n740), .ZN(n749) );
  NAND2_X1 U826 ( .A1(G8), .A2(n729), .ZN(n730) );
  NOR2_X1 U827 ( .A1(n731), .A2(G168), .ZN(n732) );
  NOR2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U829 ( .A1(n750), .A2(G286), .ZN(n739) );
  XNOR2_X1 U830 ( .A(n739), .B(n738), .ZN(n745) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n780), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U834 ( .A1(G303), .A2(n743), .ZN(n744) );
  NAND2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n746), .A2(G8), .ZN(n748) );
  XNOR2_X1 U837 ( .A(KEYINPUT32), .B(KEYINPUT96), .ZN(n747) );
  XNOR2_X1 U838 ( .A(n748), .B(n747), .ZN(n775) );
  NAND2_X1 U839 ( .A1(n749), .A2(G8), .ZN(n754) );
  INV_X1 U840 ( .A(n750), .ZN(n751) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n776) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n980) );
  AND2_X1 U844 ( .A1(n776), .A2(n980), .ZN(n755) );
  INV_X1 U845 ( .A(n980), .ZN(n757) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U848 ( .A1(n763), .A2(n756), .ZN(n984) );
  NOR2_X1 U849 ( .A1(n757), .A2(n984), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n519), .A2(n760), .ZN(n762) );
  INV_X1 U851 ( .A(KEYINPUT33), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n763), .A2(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U854 ( .A1(n780), .A2(n764), .ZN(n766) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n992) );
  NOR2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U858 ( .A(n769), .B(KEYINPUT97), .ZN(n774) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n770) );
  XNOR2_X1 U860 ( .A(n770), .B(KEYINPUT89), .ZN(n771) );
  XNOR2_X1 U861 ( .A(n771), .B(KEYINPUT24), .ZN(n772) );
  NOR2_X1 U862 ( .A1(n780), .A2(n772), .ZN(n773) );
  NOR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n783) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n779) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n817) );
  XNOR2_X1 U870 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NAND2_X1 U871 ( .A1(n904), .A2(G140), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G104), .A2(n902), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U874 ( .A(KEYINPUT34), .B(n786), .ZN(n792) );
  NAND2_X1 U875 ( .A1(n898), .A2(G128), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G116), .A2(n899), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U878 ( .A(KEYINPUT84), .B(n789), .Z(n790) );
  XNOR2_X1 U879 ( .A(KEYINPUT35), .B(n790), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U881 ( .A(n793), .B(KEYINPUT36), .Z(n794) );
  XNOR2_X1 U882 ( .A(KEYINPUT85), .B(n794), .ZN(n877) );
  NOR2_X1 U883 ( .A1(n826), .A2(n877), .ZN(n928) );
  NAND2_X1 U884 ( .A1(G160), .A2(G40), .ZN(n795) );
  NOR2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n829) );
  NAND2_X1 U886 ( .A1(n928), .A2(n829), .ZN(n797) );
  XNOR2_X1 U887 ( .A(n797), .B(KEYINPUT86), .ZN(n824) );
  INV_X1 U888 ( .A(n824), .ZN(n798) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n986) );
  XOR2_X1 U890 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n800) );
  NAND2_X1 U891 ( .A1(G105), .A2(n902), .ZN(n799) );
  XNOR2_X1 U892 ( .A(n800), .B(n799), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G141), .A2(n904), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G117), .A2(n899), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n898), .A2(G129), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n879) );
  AND2_X1 U899 ( .A1(n879), .A2(G1996), .ZN(n921) );
  NAND2_X1 U900 ( .A1(G107), .A2(n899), .ZN(n809) );
  NAND2_X1 U901 ( .A1(G131), .A2(n904), .ZN(n807) );
  XOR2_X1 U902 ( .A(KEYINPUT87), .B(n807), .Z(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n898), .A2(G119), .ZN(n811) );
  NAND2_X1 U905 ( .A1(G95), .A2(n902), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n876) );
  INV_X1 U908 ( .A(G1991), .ZN(n948) );
  NOR2_X1 U909 ( .A1(n876), .A2(n948), .ZN(n927) );
  OR2_X1 U910 ( .A1(n921), .A2(n927), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n814), .A2(n829), .ZN(n818) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n879), .ZN(n932) );
  INV_X1 U913 ( .A(n818), .ZN(n821) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n819) );
  AND2_X1 U915 ( .A1(n948), .A2(n876), .ZN(n923) );
  NOR2_X1 U916 ( .A1(n819), .A2(n923), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n932), .A2(n822), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n826), .A2(n877), .ZN(n929) );
  NAND2_X1 U922 ( .A1(n827), .A2(n929), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n830), .B(KEYINPUT98), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n834) );
  XOR2_X1 U926 ( .A(KEYINPUT99), .B(KEYINPUT40), .Z(n833) );
  XNOR2_X1 U927 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U928 ( .A1(n835), .A2(G2106), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n836), .B(KEYINPUT100), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U931 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n839), .A2(n838), .ZN(G188) );
  XNOR2_X1 U934 ( .A(G120), .B(KEYINPUT101), .ZN(G236) );
  INV_X1 U936 ( .A(G132), .ZN(G219) );
  INV_X1 U937 ( .A(G108), .ZN(G238) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G82), .ZN(G220) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n842), .B(KEYINPUT102), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  XOR2_X1 U944 ( .A(KEYINPUT111), .B(n843), .Z(n845) );
  XNOR2_X1 U945 ( .A(G171), .B(n975), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n847) );
  XOR2_X1 U947 ( .A(n978), .B(G286), .Z(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  NOR2_X1 U949 ( .A1(G37), .A2(n848), .ZN(G397) );
  XOR2_X1 U950 ( .A(G2100), .B(G2096), .Z(n850) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2678), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(G2072), .Z(n852) );
  XNOR2_X1 U954 ( .A(G2090), .B(G2067), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U957 ( .A(G2084), .B(G2078), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(G227) );
  XOR2_X1 U959 ( .A(G2474), .B(G1991), .Z(n858) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1981), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U962 ( .A(n859), .B(KEYINPUT103), .Z(n861) );
  XNOR2_X1 U963 ( .A(G1971), .B(G1986), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U965 ( .A(G1976), .B(G1956), .Z(n863) );
  XNOR2_X1 U966 ( .A(G1966), .B(G1961), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U968 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U969 ( .A(KEYINPUT41), .B(KEYINPUT104), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U971 ( .A1(n899), .A2(G112), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n904), .A2(G136), .ZN(n869) );
  NAND2_X1 U973 ( .A1(G100), .A2(n902), .ZN(n868) );
  NAND2_X1 U974 ( .A1(n869), .A2(n868), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n898), .A2(G124), .ZN(n870) );
  XOR2_X1 U976 ( .A(KEYINPUT44), .B(n870), .Z(n871) );
  NOR2_X1 U977 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n875), .B(KEYINPUT105), .ZN(G162) );
  XOR2_X1 U980 ( .A(G162), .B(n876), .Z(n878) );
  XNOR2_X1 U981 ( .A(n878), .B(n877), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n882) );
  XNOR2_X1 U983 ( .A(G160), .B(G164), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n882), .B(n881), .ZN(n886) );
  XOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n884) );
  XNOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U988 ( .A(n886), .B(n885), .Z(n897) );
  XNOR2_X1 U989 ( .A(KEYINPUT109), .B(KEYINPUT47), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n898), .A2(G127), .ZN(n888) );
  NAND2_X1 U991 ( .A1(G115), .A2(n899), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n904), .A2(G139), .ZN(n891) );
  XNOR2_X1 U995 ( .A(n891), .B(KEYINPUT108), .ZN(n893) );
  NAND2_X1 U996 ( .A1(G103), .A2(n902), .ZN(n892) );
  NAND2_X1 U997 ( .A1(n893), .A2(n892), .ZN(n894) );
  NOR2_X1 U998 ( .A1(n895), .A2(n894), .ZN(n938) );
  XNOR2_X1 U999 ( .A(n938), .B(n920), .ZN(n896) );
  XNOR2_X1 U1000 ( .A(n897), .B(n896), .ZN(n911) );
  NAND2_X1 U1001 ( .A1(n898), .A2(G130), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(G118), .A2(n899), .ZN(n900) );
  NAND2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(G106), .A2(n902), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n903), .B(KEYINPUT106), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n904), .ZN(n905) );
  NAND2_X1 U1007 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1008 ( .A(n907), .B(KEYINPUT45), .Z(n908) );
  NOR2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1010 ( .A(n911), .B(n910), .Z(n912) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n912), .ZN(G395) );
  NOR2_X1 U1012 ( .A1(G401), .A2(n919), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1015 ( .A1(G397), .A2(n914), .ZN(n915) );
  NAND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n917), .A2(G395), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT112), .ZN(G308) );
  INV_X1 U1019 ( .A(G308), .ZN(G225) );
  INV_X1 U1020 ( .A(n919), .ZN(G319) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n925) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n937) );
  INV_X1 U1026 ( .A(n928), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n935) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n933), .B(KEYINPUT51), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(G2072), .B(n938), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(G164), .B(G2078), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT113), .B(n941), .Z(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT50), .B(n942), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  XOR2_X1 U1040 ( .A(KEYINPUT55), .B(KEYINPUT114), .Z(n968) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n968), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n947), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1043 ( .A(G25), .B(n948), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n949), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G2072), .B(G33), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(n952), .B(KEYINPUT115), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(n955), .B(G27), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n960), .B(KEYINPUT53), .ZN(n967) );
  XNOR2_X1 U1055 ( .A(G2090), .B(G35), .ZN(n965) );
  XOR2_X1 U1056 ( .A(G34), .B(KEYINPUT117), .Z(n962) );
  XNOR2_X1 U1057 ( .A(G2084), .B(KEYINPUT54), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(n962), .B(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n963), .B(KEYINPUT116), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(n969), .B(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT118), .B(n970), .ZN(n972) );
  INV_X1 U1064 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(G11), .ZN(n1030) );
  INV_X1 U1067 ( .A(G16), .ZN(n1026) );
  XNOR2_X1 U1068 ( .A(KEYINPUT56), .B(KEYINPUT119), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n1026), .B(n974), .ZN(n998) );
  XNOR2_X1 U1070 ( .A(G1348), .B(n975), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(G171), .B(G1961), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n990) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n978), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(G1971), .A2(G303), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(G1956), .B(G299), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(KEYINPUT120), .B(n991), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G168), .B(G1966), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(KEYINPUT57), .B(n994), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1028) );
  XNOR2_X1 U1088 ( .A(G1961), .B(KEYINPUT121), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n999), .B(G5), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(G1976), .B(KEYINPUT126), .Z(n1000) );
  XNOR2_X1 U1091 ( .A(G23), .B(n1000), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(G24), .B(G1986), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT58), .B(n1005), .Z(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1023) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1020) );
  XNOR2_X1 U1099 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n1008) );
  XNOR2_X1 U1100 ( .A(n1008), .B(KEYINPUT60), .ZN(n1018) );
  XOR2_X1 U1101 ( .A(G1956), .B(G20), .Z(n1013) );
  XNOR2_X1 U1102 ( .A(G1341), .B(G19), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(G6), .B(G1981), .ZN(n1009) );
  NOR2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1105 ( .A(KEYINPUT122), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1106 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XOR2_X1 U1107 ( .A(KEYINPUT59), .B(G1348), .Z(n1014) );
  XNOR2_X1 U1108 ( .A(G4), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1109 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1110 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NOR2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1112 ( .A(n1021), .B(KEYINPUT125), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

