//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G190gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G190gat), .Z(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(KEYINPUT28), .A3(new_n213), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n211), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OR3_X1    g018(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n220), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(KEYINPUT26), .B2(new_n220), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT24), .B1(new_n209), .B2(new_n210), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G183gat), .B2(new_n215), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n224), .A2(new_n226), .B1(new_n209), .B2(new_n210), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n239), .B2(new_n235), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT73), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244));
  NAND2_X1  g043(.A1(G226gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n223), .A2(new_n246), .A3(new_n241), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n240), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n250), .A2(new_n251), .B1(new_n222), .B2(new_n219), .ZN(new_n252));
  INV_X1    g051(.A(new_n245), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n208), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT74), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n243), .A2(new_n257), .A3(new_n253), .A4(new_n247), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n245), .B1(new_n252), .B2(KEYINPUT29), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n257), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n253), .A3(new_n247), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n208), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n256), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G64gat), .B(G92gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT75), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n251), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT66), .B1(new_n238), .B2(new_n240), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n223), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n253), .B1(new_n273), .B2(new_n244), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n262), .B1(new_n274), .B2(KEYINPUT74), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n264), .B1(new_n275), .B2(new_n258), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(new_n255), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n268), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n270), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n276), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n282), .A2(KEYINPUT30), .A3(new_n256), .A4(new_n268), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n269), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G225gat), .A2(G233gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(KEYINPUT1), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(KEYINPUT1), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n290), .B2(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT77), .B(G155gat), .Z(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT76), .ZN(new_n304));
  XNOR2_X1  g103(.A(G155gat), .B(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(new_n302), .A3(G141gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT2), .B1(new_n301), .B2(new_n303), .ZN(new_n309));
  OAI22_X1  g108(.A1(new_n299), .A2(new_n308), .B1(new_n309), .B2(new_n305), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n296), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT78), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n310), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n310), .A3(KEYINPUT78), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n288), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT83), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT39), .ZN(new_n318));
  OR3_X1    g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n316), .B2(new_n318), .ZN(new_n320));
  INV_X1    g119(.A(new_n310), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n296), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT4), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n321), .A2(KEYINPUT4), .A3(new_n295), .A4(new_n293), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n288), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n319), .A2(new_n320), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(KEYINPUT39), .ZN(new_n332));
  XNOR2_X1  g131(.A(G1gat), .B(G29gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT0), .ZN(new_n334));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(KEYINPUT40), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT84), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n314), .A2(new_n288), .A3(new_n315), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(new_n287), .B1(new_n342), .B2(KEYINPUT5), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n287), .A4(new_n328), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n340), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n346), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(KEYINPUT5), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n344), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n350), .A3(KEYINPUT84), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n351), .A3(new_n337), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n339), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT40), .B1(new_n331), .B2(new_n338), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n286), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT31), .B(G50gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  OAI21_X1  g158(.A(new_n322), .B1(new_n208), .B2(KEYINPUT29), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n310), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n264), .B1(new_n323), .B2(new_n244), .ZN(new_n363));
  OAI21_X1  g162(.A(G22gat), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n362), .A2(new_n363), .A3(G22gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  OR3_X1    g168(.A1(new_n362), .A2(new_n363), .A3(G22gat), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(new_n364), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n359), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(KEYINPUT81), .B(new_n359), .C1(new_n368), .C2(new_n371), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n367), .B1(new_n365), .B2(new_n366), .ZN(new_n377));
  INV_X1    g176(.A(new_n359), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n370), .A2(new_n369), .A3(new_n364), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT82), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n377), .A2(new_n379), .A3(new_n382), .A4(new_n378), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n376), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT38), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n268), .B1(new_n265), .B2(KEYINPUT37), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT37), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n387), .A2(new_n388), .B1(new_n389), .B2(new_n277), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n269), .B1(new_n277), .B2(new_n389), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT85), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n386), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n256), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(new_n278), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n348), .A2(new_n350), .A3(new_n337), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n336), .B1(new_n343), .B2(new_n346), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n401), .B(new_n336), .C1(new_n343), .C2(new_n346), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n352), .A2(new_n400), .A3(new_n397), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n248), .A2(new_n254), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n389), .B1(new_n404), .B2(new_n208), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n263), .B2(new_n208), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n268), .A2(KEYINPUT38), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n406), .B(new_n407), .C1(new_n265), .C2(KEYINPUT37), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n395), .A2(new_n398), .A3(new_n403), .A4(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n356), .B(new_n385), .C1(new_n393), .C2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT69), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n296), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n252), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n296), .B(new_n411), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n273), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT64), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n419), .B(KEYINPUT34), .Z(new_n420));
  XNOR2_X1  g219(.A(G15gat), .B(G43gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n413), .A2(new_n415), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n417), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n418), .B1(new_n413), .B2(new_n415), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT32), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n427), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n425), .B(KEYINPUT32), .C1(new_n426), .C2(new_n423), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n420), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT72), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n434), .A3(new_n420), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT36), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(KEYINPUT72), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n438), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(new_n435), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT36), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n436), .A2(KEYINPUT36), .A3(new_n438), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT71), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n410), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n400), .A2(new_n397), .A3(new_n402), .A4(new_n396), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n452), .A2(new_n398), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n286), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n398), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(new_n281), .A3(new_n285), .A4(KEYINPUT80), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n385), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n444), .A2(new_n385), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n443), .A2(new_n435), .A3(KEYINPUT72), .ZN(new_n463));
  INV_X1    g262(.A(new_n441), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT86), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n439), .A2(new_n466), .A3(new_n441), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n403), .A2(new_n398), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n385), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n286), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n450), .A2(new_n459), .B1(new_n462), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n475));
  XNOR2_X1  g274(.A(G43gat), .B(G50gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  NAND2_X1  g276(.A1(G29gat), .A2(G36gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g280(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n482));
  OAI22_X1  g281(.A1(new_n476), .A2(KEYINPUT15), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  OR3_X1    g285(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n477), .B1(new_n489), .B2(new_n478), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n475), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n480), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n477), .A3(new_n478), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n489), .A2(new_n478), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n496), .B(KEYINPUT89), .C1(new_n497), .C2(new_n477), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n491), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT92), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT90), .ZN(new_n503));
  INV_X1    g302(.A(G1gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT16), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(KEYINPUT90), .A3(G1gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n502), .B2(G1gat), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n508), .A2(new_n507), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(new_n505), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n501), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n496), .B(KEYINPUT17), .C1(new_n497), .C2(new_n477), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n513), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n515), .A3(new_n505), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT92), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n500), .A2(new_n518), .A3(new_n519), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n491), .A2(new_n498), .A3(new_n521), .A4(new_n520), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT18), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n491), .A2(new_n498), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n520), .A2(new_n521), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n525), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(KEYINPUT93), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n524), .B(KEYINPUT13), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n528), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n533), .A2(KEYINPUT94), .A3(new_n536), .A4(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G113gat), .B(G141gat), .Z(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT87), .B(G197gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT11), .B(G169gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT12), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n527), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n527), .B2(new_n540), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n474), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(G85gat), .A3(G92gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  INV_X1    g356(.A(G92gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G99gat), .B(G106gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(new_n559), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n529), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT41), .ZN(new_n569));
  NAND2_X1  g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570));
  OAI22_X1  g369(.A1(new_n568), .A2(KEYINPUT97), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n500), .A2(new_n519), .A3(new_n565), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n569), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n576), .A2(new_n579), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584));
  NAND2_X1  g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G64gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(G57gat), .ZN(new_n590));
  INV_X1    g389(.A(G57gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(G64gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n588), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(new_n586), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n584), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n594), .A2(new_n586), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n591), .A2(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n589), .A2(G57gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G71gat), .B(G78gat), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n597), .A2(new_n600), .A3(new_n601), .A4(new_n588), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G127gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n530), .B1(new_n604), .B2(new_n603), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT96), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G155gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n612), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  XOR2_X1   g419(.A(new_n620), .B(KEYINPUT100), .Z(new_n621));
  INV_X1    g420(.A(G230gat), .ZN(new_n622));
  INV_X1    g421(.A(G233gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n596), .A2(new_n563), .A3(new_n602), .A4(new_n564), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n593), .A2(new_n584), .A3(new_n595), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n598), .A2(new_n599), .B1(new_n594), .B2(new_n586), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n601), .B1(new_n630), .B2(new_n597), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n555), .A2(new_n561), .A3(new_n559), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n561), .B1(new_n555), .B2(new_n559), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n632), .A2(KEYINPUT99), .A3(KEYINPUT10), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n603), .A2(new_n565), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n626), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n624), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n626), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n624), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n621), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(KEYINPUT101), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(KEYINPUT101), .ZN(new_n648));
  INV_X1    g447(.A(new_n620), .ZN(new_n649));
  OR3_X1    g448(.A1(new_n641), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n583), .A2(new_n617), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n550), .A2(new_n453), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n550), .A2(new_n286), .A3(new_n654), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n660), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n658), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(KEYINPUT42), .B2(new_n660), .ZN(G1325gat));
  NAND2_X1  g461(.A1(new_n550), .A2(new_n654), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n449), .A2(KEYINPUT103), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n449), .A2(KEYINPUT103), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n468), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n663), .B2(new_n669), .ZN(G1326gat));
  OAI21_X1  g469(.A(KEYINPUT104), .B1(new_n663), .B2(new_n385), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n550), .A2(new_n672), .A3(new_n458), .A4(new_n654), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n674), .B(new_n676), .ZN(G1327gat));
  NOR3_X1   g476(.A1(new_n583), .A2(new_n617), .A3(new_n651), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n550), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n455), .A2(G29gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT105), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n550), .A2(new_n683), .A3(new_n678), .A4(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n474), .B2(new_n583), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n462), .A2(new_n473), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n459), .A2(new_n410), .A3(new_n449), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(KEYINPUT44), .A3(new_n582), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n617), .A2(new_n549), .A3(new_n651), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G29gat), .B1(new_n696), .B2(new_n455), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n682), .A2(KEYINPUT45), .A3(new_n684), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n687), .A2(new_n697), .A3(new_n698), .ZN(G1328gat));
  INV_X1    g498(.A(new_n286), .ZN(new_n700));
  OAI21_X1  g499(.A(G36gat), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n700), .A2(G36gat), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT46), .B1(new_n679), .B2(new_n702), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n679), .A2(KEYINPUT46), .A3(new_n702), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(G1329gat));
  INV_X1    g504(.A(new_n449), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n689), .A2(new_n693), .A3(new_n706), .A4(new_n695), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G43gat), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n668), .A2(G43gat), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n708), .B(KEYINPUT47), .C1(new_n679), .C2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n679), .A2(new_n709), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n664), .A2(new_n665), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n689), .A2(new_n693), .A3(new_n712), .A4(new_n695), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(G43gat), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n710), .B1(new_n714), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g514(.A1(new_n385), .A2(G50gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n679), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n689), .A2(new_n693), .A3(new_n458), .A4(new_n695), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(G50gat), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n721));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n679), .B2(new_n717), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n550), .A2(new_n723), .A3(new_n678), .A4(new_n716), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(KEYINPUT48), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n719), .A2(G50gat), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n720), .A2(new_n721), .B1(new_n725), .B2(new_n726), .ZN(G1331gat));
  INV_X1    g526(.A(new_n617), .ZN(new_n728));
  INV_X1    g527(.A(new_n548), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n527), .A2(new_n540), .A3(new_n546), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n728), .A2(new_n731), .A3(new_n582), .A4(new_n652), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n692), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n455), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(new_n591), .ZN(G1332gat));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n692), .A2(KEYINPUT108), .A3(new_n732), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n700), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n737), .A2(new_n743), .A3(new_n738), .A4(new_n739), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n742), .B1(new_n741), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1333gat));
  NAND4_X1  g546(.A1(new_n737), .A2(G71gat), .A3(new_n712), .A4(new_n738), .ZN(new_n748));
  INV_X1    g547(.A(G71gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n733), .B2(new_n668), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n458), .A3(new_n738), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g553(.A1(new_n731), .A2(new_n617), .A3(new_n652), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n694), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n455), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n410), .A2(new_n449), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n385), .B1(new_n454), .B2(new_n456), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI22_X1  g559(.A1(KEYINPUT35), .A2(new_n461), .B1(new_n468), .B2(new_n472), .ZN(new_n761));
  OAI211_X1 g560(.A(KEYINPUT110), .B(new_n582), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n731), .A2(new_n617), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT110), .B1(new_n692), .B2(new_n582), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT51), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n474), .B2(new_n583), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n768), .A2(new_n769), .A3(new_n763), .A4(new_n762), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n455), .A2(new_n652), .A3(G85gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n766), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n772), .ZN(G1336gat));
  NOR3_X1   g572(.A1(new_n700), .A2(G92gat), .A3(new_n652), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n769), .A2(KEYINPUT111), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n764), .B2(new_n765), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n768), .A2(new_n763), .A3(new_n762), .A4(new_n776), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n689), .A2(new_n693), .A3(new_n286), .A4(new_n755), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT52), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n770), .A3(new_n774), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n781), .B2(G92gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n756), .B2(new_n666), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n668), .A2(G99gat), .A3(new_n652), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT112), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n766), .A2(new_n790), .A3(new_n770), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(G1338gat));
  NOR3_X1   g591(.A1(new_n385), .A2(new_n652), .A3(G106gat), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n778), .B2(new_n779), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n689), .A2(new_n693), .A3(new_n458), .A4(new_n755), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n766), .A2(new_n770), .A3(new_n793), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n796), .B2(G106gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1339gat));
  NOR2_X1   g601(.A1(new_n653), .A2(new_n731), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n637), .A2(new_n624), .A3(new_n640), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n641), .A3(new_n805), .ZN(new_n806));
  AOI211_X1 g605(.A(KEYINPUT54), .B(new_n624), .C1(new_n637), .C2(new_n640), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT113), .B1(new_n807), .B2(new_n620), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n637), .A2(new_n640), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n805), .A3(new_n644), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n811), .A3(new_n649), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n806), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n650), .B1(new_n813), .B2(KEYINPUT55), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n815), .A3(KEYINPUT55), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n804), .A2(new_n641), .A3(new_n805), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n807), .A2(KEYINPUT113), .A3(new_n620), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n811), .B1(new_n810), .B2(new_n649), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT55), .B(new_n817), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n814), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n536), .B1(new_n533), .B2(new_n534), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n545), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n822), .A2(new_n730), .A3(new_n582), .A4(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n730), .A2(new_n651), .A3(new_n825), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n822), .B2(new_n731), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n828), .B2(new_n582), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n617), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT115), .B(new_n826), .C1(new_n828), .C2(new_n582), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n803), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n458), .A3(new_n668), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n286), .A2(new_n455), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n549), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n833), .A2(new_n455), .ZN(new_n838));
  INV_X1    g637(.A(new_n460), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n286), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n549), .A2(G113gat), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT116), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n837), .B1(new_n841), .B2(new_n843), .ZN(G1340gat));
  INV_X1    g643(.A(new_n841), .ZN(new_n845));
  AOI21_X1  g644(.A(G120gat), .B1(new_n845), .B2(new_n651), .ZN(new_n846));
  INV_X1    g645(.A(G120gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n836), .A2(new_n847), .A3(new_n652), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n848), .ZN(G1341gat));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n608), .A3(new_n617), .ZN(new_n850));
  OAI21_X1  g649(.A(G127gat), .B1(new_n836), .B2(new_n728), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1342gat));
  NOR3_X1   g651(.A1(new_n841), .A2(G134gat), .A3(new_n583), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n836), .B2(new_n583), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(KEYINPUT117), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(KEYINPUT117), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n855), .B(new_n856), .C1(new_n858), .C2(new_n859), .ZN(G1343gat));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n833), .B2(new_n385), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  INV_X1    g662(.A(new_n650), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n815), .B1(new_n813), .B2(KEYINPUT55), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n549), .B1(new_n870), .B2(KEYINPUT118), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n822), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n827), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n826), .B1(new_n874), .B2(new_n582), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n803), .B1(new_n875), .B2(new_n728), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n385), .A2(new_n861), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n863), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n827), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n731), .B1(new_n822), .B2(new_n872), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n870), .A2(KEYINPUT118), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n583), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n617), .B1(new_n884), .B2(new_n826), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT119), .B(new_n877), .C1(new_n885), .C2(new_n803), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n879), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n449), .A2(new_n835), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n731), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G141gat), .ZN(new_n890));
  AND4_X1   g689(.A1(new_n458), .A2(new_n838), .A3(new_n700), .A4(new_n666), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n300), .A3(new_n731), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT58), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n890), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1344gat));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n887), .A2(new_n888), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n898), .B(G148gat), .C1(new_n899), .C2(new_n652), .ZN(new_n900));
  INV_X1    g699(.A(new_n833), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n458), .ZN(new_n902));
  INV_X1    g701(.A(new_n885), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n803), .B(KEYINPUT122), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n385), .A2(KEYINPUT57), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n902), .A2(KEYINPUT57), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n888), .A2(KEYINPUT121), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n888), .A2(KEYINPUT121), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n652), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n302), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n900), .B1(new_n898), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n891), .A2(new_n302), .A3(new_n651), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n891), .A2(KEYINPUT120), .A3(new_n302), .A4(new_n651), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n912), .A2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(new_n298), .B1(new_n899), .B2(new_n728), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n728), .A2(new_n298), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n891), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1346gat));
  OAI21_X1  g721(.A(G162gat), .B1(new_n899), .B2(new_n583), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n583), .A2(G162gat), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n891), .A2(KEYINPUT123), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT123), .B1(new_n891), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n700), .A2(new_n453), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n834), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n229), .A3(new_n549), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT124), .B1(new_n901), .B2(new_n455), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n833), .A2(new_n932), .A3(new_n453), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n839), .A2(new_n700), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(new_n731), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n930), .B1(new_n936), .B2(new_n229), .ZN(G1348gat));
  OAI21_X1  g736(.A(G176gat), .B1(new_n929), .B2(new_n652), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n935), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n651), .A2(new_n230), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(G1349gat));
  NOR2_X1   g740(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n942));
  AND2_X1   g741(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n943));
  OAI21_X1  g742(.A(G183gat), .B1(new_n929), .B2(new_n728), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n728), .A2(new_n214), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n935), .B(new_n945), .C1(new_n931), .C2(new_n933), .ZN(new_n946));
  AOI211_X1 g745(.A(new_n942), .B(new_n943), .C1(new_n944), .C2(new_n946), .ZN(new_n947));
  AND4_X1   g746(.A1(KEYINPUT125), .A2(new_n944), .A3(new_n946), .A4(KEYINPUT60), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(G1350gat));
  NOR2_X1   g748(.A1(new_n668), .A2(new_n458), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n901), .A2(new_n582), .A3(new_n950), .A4(new_n928), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G190gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT126), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n955), .A3(G190gat), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n953), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n582), .A2(new_n217), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n957), .A2(new_n958), .B1(new_n939), .B2(new_n959), .ZN(G1351gat));
  AND2_X1   g759(.A1(new_n666), .A2(new_n928), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n907), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(G197gat), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n962), .A2(new_n963), .A3(new_n549), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n712), .A2(new_n385), .A3(new_n700), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n934), .A2(new_n731), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n964), .B1(new_n963), .B2(new_n966), .ZN(G1352gat));
  NOR2_X1   g766(.A1(new_n652), .A2(G204gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n934), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n934), .A2(new_n971), .A3(new_n965), .A4(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n902), .A2(KEYINPUT57), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n905), .A2(new_n906), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n973), .A2(new_n651), .A3(new_n974), .A4(new_n961), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G204gat), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n970), .B(new_n972), .C1(new_n978), .C2(new_n979), .ZN(G1353gat));
  NAND3_X1  g779(.A1(new_n907), .A2(new_n617), .A3(new_n961), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n934), .A2(new_n965), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n617), .A2(new_n203), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n982), .A2(new_n983), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  OAI21_X1  g785(.A(G218gat), .B1(new_n962), .B2(new_n583), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n582), .A2(new_n204), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n984), .B2(new_n988), .ZN(G1355gat));
endmodule


