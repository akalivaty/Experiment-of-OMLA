//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067;
  XNOR2_X1  g000(.A(KEYINPUT72), .B(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G234), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT73), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT16), .ZN(new_n197));
  OR3_X1    g011(.A1(new_n195), .A2(KEYINPUT16), .A3(G140), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G146), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n196), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT24), .B(G110), .Z(new_n203));
  XNOR2_X1  g017(.A(G119), .B(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(G128), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n212), .A2(G110), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT74), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n205), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OR3_X1    g029(.A1(new_n212), .A2(new_n214), .A3(G110), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n202), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n197), .A2(new_n198), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n200), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n199), .ZN(new_n221));
  AOI22_X1  g035(.A1(G110), .A2(new_n212), .B1(new_n203), .B2(new_n204), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT22), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n226), .B(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n218), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n227), .ZN(new_n229));
  INV_X1    g043(.A(new_n223), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n217), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n188), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n192), .B1(new_n232), .B2(KEYINPUT25), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n228), .A2(new_n234), .A3(new_n188), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n192), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT75), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n228), .A2(new_n239), .A3(new_n231), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n228), .B2(new_n231), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT11), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G137), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(G137), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n246), .A2(new_n248), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT66), .B1(new_n245), .B2(G137), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n250), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n245), .A2(KEYINPUT66), .A3(G137), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n200), .A2(G143), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n210), .B1(new_n256), .B2(KEYINPUT1), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT65), .B1(new_n200), .B2(G143), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G146), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT64), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT64), .A2(G143), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n200), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n257), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT64), .A2(G143), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(G146), .A3(new_n263), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n269), .A2(new_n256), .A3(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n251), .B(new_n255), .C1(new_n267), .C2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n246), .A2(new_n250), .A3(new_n248), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G131), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n251), .ZN(new_n275));
  AND2_X1   g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NOR2_X1   g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G146), .B1(new_n268), .B2(new_n263), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n258), .A2(new_n261), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n269), .A2(new_n256), .A3(new_n276), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n275), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n272), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g100(.A1(KEYINPUT2), .A2(G113), .ZN(new_n287));
  NOR2_X1   g101(.A1(KEYINPUT2), .A2(G113), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G116), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT67), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G116), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n293), .A3(G119), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n290), .A2(G119), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n289), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(new_n289), .A3(new_n296), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n272), .A2(KEYINPUT30), .A3(new_n283), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n286), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n224), .A3(G210), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT27), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n304), .B(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT26), .ZN(new_n307));
  INV_X1    g121(.A(G101), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n299), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(new_n297), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n272), .A2(new_n311), .A3(new_n283), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n302), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT31), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT68), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n316), .A3(KEYINPUT31), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n272), .A2(new_n311), .A3(new_n283), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n311), .B1(new_n272), .B2(new_n283), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT69), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n312), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n309), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n302), .A2(new_n329), .A3(new_n309), .A4(new_n312), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n315), .A2(new_n317), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(G472), .A2(G902), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n331), .A2(KEYINPUT32), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT32), .B1(new_n331), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n302), .A2(new_n312), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n327), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n320), .A2(new_n323), .A3(new_n309), .A4(new_n325), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT70), .B1(new_n339), .B2(new_n338), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n188), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n339), .A2(KEYINPUT70), .A3(new_n338), .ZN(new_n343));
  OAI21_X1  g157(.A(G472), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n243), .B1(new_n335), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n303), .A2(new_n224), .A3(G143), .A4(G214), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT64), .B(G143), .ZN(new_n347));
  INV_X1    g161(.A(G214), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n348), .A2(G237), .A3(G953), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n346), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G131), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT17), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n303), .A2(new_n224), .A3(G214), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n268), .A3(new_n263), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n249), .A3(new_n346), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n350), .A2(KEYINPUT17), .A3(G131), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n356), .A2(new_n220), .A3(new_n199), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(KEYINPUT18), .A2(G131), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n354), .A2(KEYINPUT83), .A3(new_n346), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT83), .B1(new_n354), .B2(new_n346), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n359), .B(new_n346), .C1(new_n347), .C2(new_n349), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT85), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT85), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n354), .A2(new_n366), .A3(new_n359), .A4(new_n346), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n201), .A2(KEYINPUT84), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n194), .A2(new_n196), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G146), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(KEYINPUT84), .A3(G146), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n363), .A2(new_n368), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT88), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n358), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n357), .A2(new_n220), .A3(new_n199), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n365), .A2(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n356), .A2(new_n382), .B1(new_n383), .B2(new_n363), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n378), .B1(new_n384), .B2(KEYINPUT89), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n358), .A2(new_n375), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT89), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n381), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G475), .B1(new_n389), .B2(G902), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n197), .A2(G146), .A3(new_n198), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n351), .B2(new_n355), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT19), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n394), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n396), .A2(new_n370), .A3(new_n397), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n370), .A2(new_n393), .A3(new_n394), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n200), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n383), .A2(new_n363), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n378), .B1(new_n401), .B2(KEYINPUT87), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n400), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n375), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n381), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n407), .A2(KEYINPUT20), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n384), .A2(new_n380), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n375), .A2(KEYINPUT87), .A3(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(new_n378), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n401), .A2(KEYINPUT87), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n411), .B1(new_n417), .B2(new_n408), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n390), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n407), .B2(new_n409), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n411), .A3(new_n408), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT90), .A3(new_n390), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n347), .A2(new_n210), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT13), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n260), .A2(G128), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n245), .B1(new_n426), .B2(new_n427), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OR3_X1    g246(.A1(new_n426), .A2(G134), .A3(new_n428), .ZN(new_n433));
  INV_X1    g247(.A(G107), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n291), .A2(new_n293), .A3(G122), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT91), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n290), .A2(G122), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n435), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n439), .A2(new_n434), .A3(new_n440), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n432), .B(new_n433), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G134), .B1(new_n426), .B2(new_n428), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n433), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT14), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n437), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT92), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n435), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n449), .B1(new_n448), .B2(new_n435), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n441), .B(new_n446), .C1(new_n454), .C2(new_n434), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT9), .B(G234), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n224), .A3(new_n187), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n444), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n444), .B2(new_n455), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n188), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G478), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI221_X1 g280(.A(new_n188), .B1(KEYINPUT15), .B2(new_n464), .C1(new_n461), .C2(new_n462), .ZN(new_n467));
  INV_X1    g281(.A(G952), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n190), .B2(new_n303), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n224), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(G898), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n466), .A2(new_n467), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n421), .A2(new_n425), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G140), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n224), .A2(G227), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n269), .A2(new_n256), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT1), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n347), .B2(new_n200), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n484), .B2(new_n210), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT77), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n269), .A2(new_n486), .A3(new_n256), .A4(new_n270), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n269), .A2(new_n256), .A3(new_n270), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT77), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n491));
  XNOR2_X1  g305(.A(G104), .B(G107), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n491), .B1(new_n492), .B2(new_n308), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n434), .A2(G104), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n377), .A2(G107), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT76), .A3(G101), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n434), .A3(G104), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n498), .A2(new_n500), .A3(new_n308), .A4(new_n495), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n493), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n490), .A2(new_n502), .ZN(new_n503));
  XOR2_X1   g317(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n275), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n498), .A2(new_n500), .A3(new_n495), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(G101), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n281), .A2(new_n509), .A3(new_n282), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(G101), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT10), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n483), .B1(G143), .B2(new_n200), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n279), .A2(new_n280), .B1(new_n210), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n516), .B2(new_n488), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n511), .A2(new_n513), .B1(new_n517), .B2(new_n502), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n505), .A2(new_n506), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n493), .A2(new_n497), .A3(new_n501), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n488), .A3(new_n516), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n503), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT12), .B1(new_n522), .B2(new_n275), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n524));
  AOI211_X1 g338(.A(new_n524), .B(new_n506), .C1(new_n503), .C2(new_n521), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n481), .B(new_n519), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n504), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n490), .B2(new_n502), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT10), .B1(new_n267), .B2(new_n271), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n512), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n530));
  OAI22_X1  g344(.A1(new_n529), .A2(new_n520), .B1(new_n530), .B2(new_n510), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n275), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n519), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n480), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G469), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n188), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n528), .A2(new_n531), .A3(new_n275), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n480), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n532), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n522), .A2(KEYINPUT12), .A3(new_n275), .ZN(new_n541));
  OAI21_X1  g355(.A(G128), .B1(new_n279), .B2(new_n483), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n542), .A2(new_n482), .B1(new_n488), .B2(KEYINPUT77), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n520), .B1(new_n543), .B2(new_n487), .ZN(new_n544));
  INV_X1    g358(.A(new_n521), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n275), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n524), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n538), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n540), .B(G469), .C1(new_n481), .C2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n536), .A2(new_n237), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n537), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G221), .B1(new_n456), .B2(G902), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G214), .B1(G237), .B2(G902), .ZN(new_n555));
  XNOR2_X1  g369(.A(G110), .B(G122), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n509), .B1(new_n310), .B2(new_n297), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(new_n530), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n294), .A2(KEYINPUT5), .A3(new_n296), .ZN(new_n560));
  INV_X1    g374(.A(G113), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT5), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n295), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n564), .A2(new_n520), .A3(new_n310), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n557), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n560), .A2(new_n563), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n502), .A2(new_n299), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n568), .B(new_n556), .C1(new_n530), .C2(new_n558), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(KEYINPUT6), .A3(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n276), .A2(new_n277), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n262), .B2(new_n266), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n269), .A2(new_n256), .A3(new_n276), .ZN(new_n573));
  OAI21_X1  g387(.A(G125), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n516), .A2(new_n195), .A3(new_n488), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT79), .B(G224), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n224), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n576), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT6), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(new_n557), .C1(new_n559), .C2(new_n565), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n570), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n583), .A2(new_n237), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(KEYINPUT7), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT80), .B1(new_n576), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n587));
  INV_X1    g401(.A(new_n585), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n587), .B(new_n588), .C1(new_n574), .C2(new_n575), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n556), .B(KEYINPUT8), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n493), .A2(new_n497), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n592), .A2(new_n501), .B1(new_n567), .B2(new_n299), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n565), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n574), .A2(KEYINPUT7), .A3(new_n575), .A4(new_n578), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT81), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n576), .A2(new_n579), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n520), .B1(new_n564), .B2(new_n310), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n568), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n598), .A2(KEYINPUT7), .B1(new_n600), .B2(new_n591), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n267), .A2(new_n271), .A3(G125), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n195), .B1(new_n281), .B2(new_n282), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n585), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n587), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n576), .A2(KEYINPUT80), .A3(new_n585), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT81), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n601), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n597), .A2(new_n609), .A3(new_n569), .ZN(new_n610));
  OAI21_X1  g424(.A(G210), .B1(G237), .B2(G902), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT82), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n584), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n584), .B2(new_n610), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n555), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n477), .A2(new_n554), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n345), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n461), .B2(new_n462), .ZN(new_n621));
  INV_X1    g435(.A(new_n462), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(KEYINPUT33), .A3(new_n460), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n189), .A2(new_n464), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n463), .A2(new_n464), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n424), .A2(KEYINPUT90), .A3(new_n390), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT90), .B1(new_n424), .B2(new_n390), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n555), .B(new_n475), .C1(new_n614), .C2(new_n615), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT93), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n328), .A2(new_n330), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n313), .A2(new_n316), .A3(KEYINPUT31), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n316), .B1(new_n313), .B2(KEYINPUT31), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n634), .B1(new_n638), .B2(new_n189), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n331), .A2(KEYINPUT93), .A3(new_n188), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(G472), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n332), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n243), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n552), .A2(new_n645), .A3(new_n553), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n641), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n633), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT34), .B(G104), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  AND3_X1   g464(.A1(new_n641), .A2(new_n644), .A3(new_n646), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT94), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n424), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n466), .A2(new_n467), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT94), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n653), .A2(new_n390), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n331), .A2(new_n188), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(new_n634), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n643), .B1(new_n663), .B2(new_n640), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n218), .A2(new_n223), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n229), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n238), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n236), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n664), .A2(new_n617), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT37), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT95), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(G110), .Z(G12));
  NOR2_X1   g487(.A1(new_n554), .A2(new_n616), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT32), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n638), .B2(new_n642), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n331), .A2(KEYINPUT32), .A3(new_n332), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n344), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n470), .B(KEYINPUT96), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n680), .B1(new_n681), .B2(new_n472), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n656), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n674), .A2(new_n678), .A3(new_n683), .A4(new_n669), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XOR2_X1   g499(.A(new_n682), .B(KEYINPUT39), .Z(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n554), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT40), .Z(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n690), .A2(KEYINPUT97), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n584), .A2(new_n610), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n612), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n584), .A2(new_n610), .A3(new_n613), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n693), .A2(KEYINPUT38), .A3(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n555), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n669), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n336), .A2(new_n309), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n318), .A2(new_n319), .ZN(new_n703));
  AOI21_X1  g517(.A(G902), .B1(new_n327), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n661), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n676), .A2(new_n677), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n654), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n421), .B2(new_n425), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n701), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n690), .B2(KEYINPUT97), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n691), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n347), .ZN(G45));
  AND2_X1   g527(.A1(new_n625), .A2(new_n626), .ZN(new_n714));
  AOI211_X1 g528(.A(new_n682), .B(new_n714), .C1(new_n421), .C2(new_n425), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n674), .A3(new_n678), .A4(new_n669), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT98), .B(G146), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G48));
  NAND2_X1  g532(.A1(new_n547), .A2(new_n541), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n539), .A2(new_n719), .B1(new_n533), .B2(new_n480), .ZN(new_n720));
  OAI21_X1  g534(.A(G469), .B1(new_n720), .B2(new_n189), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n537), .A3(new_n553), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n632), .A2(new_n678), .A3(new_n645), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n657), .A2(new_n678), .A3(new_n645), .A4(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT99), .B(G116), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G18));
  INV_X1    g543(.A(new_n477), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n616), .A2(new_n722), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n678), .A2(new_n730), .A3(new_n731), .A4(new_n669), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  NAND2_X1  g547(.A1(new_n421), .A2(new_n425), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n700), .B1(new_n693), .B2(new_n694), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n734), .A2(new_n735), .A3(new_n654), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n328), .A2(new_n314), .A3(new_n330), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n332), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT100), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(new_n740), .A3(new_n332), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n661), .B1(new_n331), .B2(new_n188), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n742), .A2(new_n743), .A3(new_n243), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n722), .A2(new_n474), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n736), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  INV_X1    g561(.A(new_n669), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n742), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n715), .A3(new_n731), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n693), .A2(new_n555), .A3(new_n694), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT101), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n753), .B1(new_n554), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n552), .A2(KEYINPUT101), .A3(new_n553), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n678), .A3(new_n645), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n715), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n752), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n554), .A2(new_n754), .ZN(new_n760));
  INV_X1    g574(.A(new_n753), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n760), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(new_n345), .A3(KEYINPUT42), .A4(new_n715), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n345), .A3(new_n683), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  NAND3_X1  g581(.A1(new_n421), .A2(new_n425), .A3(new_n627), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT43), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n421), .A2(new_n770), .A3(new_n425), .A4(new_n627), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n772), .A2(new_n664), .A3(new_n748), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT44), .Z(new_n774));
  OAI21_X1  g588(.A(new_n540), .B1(new_n481), .B2(new_n548), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n536), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n540), .B(KEYINPUT45), .C1(new_n481), .C2(new_n548), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n550), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n537), .B1(new_n779), .B2(KEYINPUT46), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n548), .A2(new_n481), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n519), .A2(new_n532), .A3(new_n481), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n776), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(G469), .A3(new_n778), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n551), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n553), .B1(new_n780), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n687), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n774), .A2(new_n761), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NAND2_X1  g604(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n784), .A2(new_n551), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n537), .A3(new_n785), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n553), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n678), .A2(new_n645), .A3(new_n753), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n791), .A2(new_n797), .A3(new_n715), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  NAND4_X1  g614(.A1(new_n749), .A2(new_n715), .A3(new_n755), .A4(new_n756), .ZN(new_n801));
  INV_X1    g615(.A(new_n682), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n708), .A2(new_n669), .A3(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n554), .A2(new_n753), .A3(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n653), .A2(new_n390), .A3(new_n655), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n678), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n683), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n801), .B(new_n806), .C1(new_n757), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT103), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT103), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n766), .A2(new_n810), .A3(new_n806), .A4(new_n801), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n748), .B1(new_n335), .B2(new_n344), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n674), .C1(new_n683), .C2(new_n715), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n553), .A2(new_n552), .A3(new_n748), .A4(new_n802), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n707), .A2(new_n815), .A3(new_n735), .A4(new_n709), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(KEYINPUT52), .A3(new_n750), .A4(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n716), .A2(new_n750), .A3(new_n684), .A4(new_n816), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n421), .A2(new_n425), .A3(new_n654), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n631), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n644), .A3(new_n641), .A4(new_n646), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n670), .A2(KEYINPUT102), .A3(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n651), .A2(new_n632), .B1(new_n345), .B2(new_n617), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n670), .A2(new_n825), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT102), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n724), .A2(new_n746), .A3(new_n727), .A4(new_n732), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n828), .A2(new_n764), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n822), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n821), .B2(KEYINPUT104), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n826), .A2(new_n827), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT102), .B1(new_n670), .B2(new_n825), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n839), .A2(new_n840), .A3(new_n832), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n764), .A3(new_n821), .A4(new_n812), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n836), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT54), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n831), .A2(new_n826), .A3(new_n827), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n764), .A2(KEYINPUT53), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n809), .A2(new_n811), .B1(new_n817), .B2(new_n820), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n477), .A2(new_n616), .A3(new_n722), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n662), .A2(G472), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n737), .A2(new_n740), .A3(new_n332), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n740), .B1(new_n737), .B2(new_n332), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n645), .A2(new_n745), .A3(new_n851), .A4(new_n854), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n813), .A2(new_n850), .B1(new_n855), .B2(new_n736), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT105), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n724), .A4(new_n727), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n832), .A2(KEYINPUT105), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n848), .A2(new_n849), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n861), .A2(KEYINPUT106), .B1(new_n842), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT106), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n848), .A2(new_n849), .A3(new_n865), .A4(new_n860), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n744), .A2(new_n680), .A3(new_n769), .A4(new_n771), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n699), .A2(new_n700), .A3(new_n723), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n769), .A2(new_n680), .A3(new_n771), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n555), .B(new_n722), .C1(new_n697), .C2(new_n698), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT50), .A4(new_n744), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n753), .A2(new_n722), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n680), .A2(new_n769), .A3(new_n771), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n243), .A2(new_n470), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n335), .A2(new_n877), .A3(new_n706), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n734), .A2(new_n627), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n878), .A2(new_n749), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n876), .A2(KEYINPUT108), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n721), .A2(new_n537), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n553), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n553), .ZN(new_n887));
  INV_X1    g701(.A(new_n537), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n792), .B2(new_n793), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT47), .B(new_n887), .C1(new_n889), .C2(new_n785), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n796), .B1(new_n795), .B2(new_n553), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT107), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n870), .B2(new_n753), .ZN(new_n894));
  INV_X1    g708(.A(new_n870), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(KEYINPUT107), .A3(new_n761), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n892), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n883), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT108), .B1(new_n876), .B2(new_n882), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n878), .A2(new_n345), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT48), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n731), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n880), .A2(new_n734), .A3(new_n627), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n469), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT111), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n876), .A2(new_n882), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT109), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT109), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n876), .A2(new_n910), .A3(new_n882), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n885), .B1(new_n791), .B2(new_n797), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT110), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n894), .B(new_n896), .C1(new_n913), .C2(KEYINPUT110), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT51), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n907), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n791), .A2(new_n797), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT110), .B1(new_n919), .B2(new_n886), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n896), .A2(new_n894), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n868), .B1(new_n922), .B2(new_n914), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n909), .A2(new_n911), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(KEYINPUT111), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n906), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n845), .B(new_n867), .C1(new_n926), .C2(KEYINPUT112), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n900), .A2(new_n905), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n912), .A2(new_n917), .A3(new_n907), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT111), .B1(new_n923), .B2(new_n924), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT112), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT113), .B1(new_n927), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n867), .A2(new_n845), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n931), .A2(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n926), .A2(KEYINPUT112), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT113), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n468), .A2(new_n224), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n934), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n884), .A2(KEYINPUT49), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n884), .A2(KEYINPUT49), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n553), .A2(new_n555), .ZN(new_n944));
  NOR4_X1   g758(.A1(new_n942), .A2(new_n943), .A3(new_n243), .A4(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n707), .A2(new_n768), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n699), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT114), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n941), .A2(KEYINPUT114), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G75));
  NOR2_X1   g766(.A1(new_n224), .A2(G952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n188), .B1(new_n863), .B2(new_n866), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT56), .B1(new_n955), .B2(new_n612), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n570), .A2(new_n582), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n580), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT55), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n954), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n956), .B2(new_n959), .ZN(G51));
  AND3_X1   g775(.A1(new_n670), .A2(KEYINPUT102), .A3(new_n825), .ZN(new_n962));
  INV_X1    g776(.A(new_n617), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n678), .A2(new_n645), .ZN(new_n964));
  OAI22_X1  g778(.A1(new_n963), .A2(new_n964), .B1(new_n633), .B2(new_n647), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n962), .A2(new_n840), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n862), .B1(new_n759), .B2(new_n763), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n860), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT106), .B1(new_n968), .B2(new_n822), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n862), .B1(new_n822), .B2(new_n834), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n866), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(KEYINPUT54), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n867), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n550), .B(KEYINPUT115), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT57), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT116), .B1(new_n976), .B2(new_n535), .ZN(new_n977));
  INV_X1    g791(.A(new_n784), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n955), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n976), .A2(KEYINPUT116), .A3(new_n535), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n953), .B1(new_n979), .B2(new_n980), .ZN(G54));
  NAND3_X1  g795(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(new_n407), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT117), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n953), .B1(new_n982), .B2(new_n407), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(G60));
  AND2_X1   g802(.A1(new_n621), .A2(new_n623), .ZN(new_n989));
  INV_X1    g803(.A(new_n935), .ZN(new_n990));
  NAND2_X1  g804(.A1(G478), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT59), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n989), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n973), .A2(new_n989), .A3(new_n992), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n993), .A2(new_n953), .A3(new_n994), .ZN(G63));
  NAND2_X1  g809(.A1(G217), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT118), .Z(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT60), .Z(new_n998));
  AND3_X1   g812(.A1(new_n971), .A2(new_n667), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n240), .A2(new_n241), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n971), .B2(new_n998), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n999), .A2(new_n1002), .A3(new_n953), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT120), .B1(new_n1003), .B2(KEYINPUT61), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n971), .A2(new_n667), .A3(new_n998), .ZN(new_n1005));
  INV_X1    g819(.A(new_n998), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n863), .B2(new_n866), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n954), .B(new_n1005), .C1(new_n1007), .C2(new_n1001), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT120), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT61), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n971), .A2(new_n998), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n953), .B1(new_n1012), .B2(new_n1000), .ZN(new_n1013));
  AOI211_X1 g827(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n1013), .C2(new_n1005), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT119), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1016));
  OAI22_X1  g830(.A1(new_n1004), .A2(new_n1011), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT121), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1003), .A2(KEYINPUT120), .A3(KEYINPUT61), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1009), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1022), .B(KEYINPUT121), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1019), .A2(new_n1023), .ZN(G66));
  INV_X1    g838(.A(new_n473), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n224), .B1(new_n1025), .B2(new_n577), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT122), .ZN(new_n1027));
  INV_X1    g841(.A(new_n841), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(new_n224), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n957), .B1(G898), .B2(new_n224), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1029), .B(new_n1030), .Z(G69));
  NAND2_X1  g845(.A1(new_n681), .A2(G953), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT126), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n789), .A2(new_n799), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n788), .A2(new_n345), .A3(new_n736), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1034), .A2(new_n764), .A3(new_n766), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n814), .A2(new_n750), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1037), .B(KEYINPUT124), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1033), .B1(new_n1039), .B2(G953), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n286), .A2(new_n301), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1041), .B(KEYINPUT123), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n398), .A2(new_n399), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1038), .B1(new_n691), .B2(new_n711), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT62), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g862(.A(new_n1048), .B(KEYINPUT125), .Z(new_n1049));
  NAND2_X1  g863(.A1(new_n630), .A2(new_n823), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n345), .A2(new_n688), .A3(new_n761), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1034), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1052), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1053));
  AOI21_X1  g867(.A(G953), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1045), .B1(new_n1054), .B2(new_n1044), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n224), .B1(G227), .B2(G900), .ZN(new_n1056));
  XNOR2_X1  g870(.A(new_n1055), .B(new_n1056), .ZN(G72));
  NAND3_X1  g871(.A1(new_n1049), .A2(new_n841), .A3(new_n1053), .ZN(new_n1058));
  XNOR2_X1  g872(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1059));
  NOR2_X1   g873(.A1(new_n661), .A2(new_n237), .ZN(new_n1060));
  XNOR2_X1  g874(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n702), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n327), .A2(new_n312), .A3(new_n302), .ZN(new_n1063));
  AND4_X1   g877(.A1(new_n702), .A2(new_n844), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g878(.A(new_n1061), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1065), .B1(new_n1039), .B2(new_n841), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n954), .B1(new_n1066), .B2(new_n1063), .ZN(new_n1067));
  NOR3_X1   g881(.A1(new_n1062), .A2(new_n1064), .A3(new_n1067), .ZN(G57));
endmodule


