//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT67), .Z(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT68), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n209), .B(new_n210), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT69), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n208), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  INV_X1    g0034(.A(KEYINPUT0), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(new_n235), .B2(new_n234), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT66), .Z(new_n238));
  NOR3_X1   g0038(.A1(new_n224), .A2(new_n225), .A3(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G68), .ZN(new_n251));
  INV_X1    g0051(.A(G68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G58), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n250), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(KEYINPUT71), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  AND3_X1   g0059(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT8), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(KEYINPUT71), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n229), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n263), .B2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n266), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n259), .A2(new_n252), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n272), .A2(new_n201), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n273), .A2(G20), .B1(G159), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT7), .B1(new_n280), .B2(new_n230), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT80), .ZN(new_n282));
  INV_X1    g0082(.A(new_n279), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(new_n276), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n230), .A2(KEYINPUT7), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n276), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n279), .ZN(new_n291));
  INV_X1    g0091(.A(new_n286), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(KEYINPUT80), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n281), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n275), .B1(new_n294), .B2(new_n252), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT16), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n268), .ZN(new_n298));
  INV_X1    g0098(.A(new_n275), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT79), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n278), .ZN(new_n301));
  NAND2_X1  g0101(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G33), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(G20), .B1(new_n303), .B2(new_n277), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT7), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n252), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n277), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n288), .A2(new_n289), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(G33), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT7), .B1(new_n309), .B2(G20), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n299), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n298), .B1(new_n311), .B2(KEYINPUT16), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n271), .B1(new_n297), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G41), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(G1), .A3(G13), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n229), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(KEYINPUT70), .A3(new_n314), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  MUX2_X1   g0120(.A(G223), .B(G226), .S(G1698), .Z(new_n321));
  NAND2_X1  g0121(.A1(new_n309), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G87), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n315), .ZN(new_n325));
  INV_X1    g0125(.A(G41), .ZN(new_n326));
  INV_X1    g0126(.A(G45), .ZN(new_n327));
  AOI21_X1  g0127(.A(G1), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G232), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n315), .A3(G274), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n324), .B2(new_n332), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT83), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n335), .A2(KEYINPUT83), .A3(new_n337), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n313), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(new_n342), .B(KEYINPUT17), .Z(new_n343));
  INV_X1    g0143(.A(KEYINPUT82), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT81), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n333), .A2(G179), .ZN(new_n347));
  OAI21_X1  g0147(.A(G169), .B1(new_n324), .B2(new_n332), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n346), .B1(new_n313), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n271), .ZN(new_n351));
  INV_X1    g0151(.A(new_n281), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT80), .B1(new_n291), .B2(new_n292), .ZN(new_n353));
  AOI211_X1 g0153(.A(new_n282), .B(new_n286), .C1(new_n290), .C2(new_n279), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G68), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT16), .B1(new_n356), .B2(new_n275), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n306), .A2(new_n310), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n275), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n268), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n351), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n347), .A2(new_n348), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(KEYINPUT18), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n345), .B1(new_n350), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT18), .B1(new_n361), .B2(new_n362), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(KEYINPUT81), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n344), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n313), .A2(new_n346), .A3(new_n349), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT81), .B1(new_n368), .B2(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n350), .A2(new_n345), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(KEYINPUT82), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n343), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n315), .A2(G238), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n331), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n317), .A2(new_n319), .ZN(new_n377));
  INV_X1    g0177(.A(G1698), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n277), .A2(new_n279), .A3(G226), .A4(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n277), .A2(new_n279), .A3(G232), .A4(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G97), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n376), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI211_X1 g0185(.A(KEYINPUT13), .B(new_n376), .C1(new_n377), .C2(new_n382), .ZN(new_n386));
  OAI21_X1  g0186(.A(G169), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT14), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n377), .A2(new_n382), .ZN(new_n389));
  INV_X1    g0189(.A(new_n376), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n383), .A2(new_n384), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(G169), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n391), .A2(new_n398), .A3(KEYINPUT13), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT76), .B1(new_n383), .B2(new_n384), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n393), .A2(KEYINPUT77), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT77), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n386), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(G179), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT78), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n393), .B(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT78), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(G179), .A4(new_n401), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n397), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n274), .A2(G50), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n230), .B2(G68), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n230), .A2(G33), .ZN(new_n413));
  INV_X1    g0213(.A(G77), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n268), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT11), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n420), .A2(new_n422), .B1(new_n269), .B2(G68), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n410), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n407), .A2(G190), .A3(new_n401), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n394), .B2(G200), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n413), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n262), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n274), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n298), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n265), .A2(new_n202), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n270), .B2(new_n202), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(KEYINPUT9), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT74), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n437), .A2(KEYINPUT74), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT10), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n280), .A2(G1698), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G222), .ZN(new_n444));
  INV_X1    g0244(.A(new_n280), .ZN(new_n445));
  INV_X1    g0245(.A(G223), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(G1698), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n444), .B1(new_n414), .B2(new_n445), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n377), .ZN(new_n449));
  INV_X1    g0249(.A(new_n331), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(G226), .B2(new_n329), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(G190), .A3(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n449), .A2(new_n451), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(new_n453), .B2(new_n336), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n442), .B1(new_n454), .B2(KEYINPUT75), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n336), .B1(new_n449), .B2(new_n451), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(G190), .B2(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n436), .A2(KEYINPUT9), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n441), .A2(new_n455), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n440), .C2(new_n439), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT75), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT10), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G179), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n453), .A2(new_n466), .ZN(new_n467));
  OAI221_X1 g0267(.A(new_n467), .B1(G169), .B2(new_n453), .C1(new_n433), .C2(new_n435), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n443), .A2(G232), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n445), .A2(G238), .A3(G1698), .ZN(new_n470));
  INV_X1    g0270(.A(G107), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n469), .B(new_n470), .C1(new_n471), .C2(new_n445), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n377), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n450), .B1(G244), .B2(new_n329), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n334), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n269), .A2(G77), .ZN(new_n477));
  XOR2_X1   g0277(.A(new_n477), .B(KEYINPUT73), .Z(new_n478));
  INV_X1    g0278(.A(new_n261), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n479), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT72), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT15), .B(G87), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n413), .ZN(new_n483));
  INV_X1    g0283(.A(new_n482), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(KEYINPUT72), .A3(new_n430), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(new_n268), .B1(new_n414), .B2(new_n265), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n476), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n475), .A2(G200), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G169), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n475), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n473), .A2(new_n466), .A3(new_n474), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n488), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n429), .A2(new_n465), .A3(new_n468), .A4(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n373), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NOR4_X1   g0301(.A1(new_n280), .A2(KEYINPUT22), .A3(G20), .A4(new_n213), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n303), .A2(new_n230), .A3(G87), .A4(new_n277), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT22), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT90), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(KEYINPUT90), .A3(KEYINPUT22), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G116), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT84), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT84), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G116), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G33), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G20), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT23), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n230), .B2(G107), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n471), .A2(KEYINPUT23), .A3(G20), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n508), .A2(new_n520), .A3(KEYINPUT24), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT24), .ZN(new_n522));
  INV_X1    g0322(.A(new_n502), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n503), .A2(KEYINPUT90), .A3(KEYINPUT22), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT90), .B1(new_n503), .B2(KEYINPUT22), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n522), .B1(new_n526), .B2(new_n519), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n268), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT25), .B1(new_n265), .B2(new_n471), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n265), .A2(KEYINPUT25), .A3(new_n471), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n263), .A2(G33), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n264), .A2(new_n532), .A3(new_n229), .A4(new_n267), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n530), .A2(new_n531), .B1(G107), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT91), .ZN(new_n536));
  INV_X1    g0336(.A(G274), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n318), .B2(new_n314), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n327), .A2(G1), .ZN(new_n539));
  XNOR2_X1  g0339(.A(KEYINPUT5), .B(G41), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n539), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n315), .ZN(new_n543));
  INV_X1    g0343(.A(G264), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G250), .A2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n216), .B2(G1698), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n303), .A3(new_n277), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n320), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n536), .B1(new_n551), .B2(new_n493), .ZN(new_n552));
  OAI211_X1 g0352(.A(KEYINPUT91), .B(G169), .C1(new_n545), .C2(new_n550), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(G179), .B2(new_n551), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n528), .A2(new_n535), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT24), .B1(new_n508), .B2(new_n520), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n526), .A2(new_n522), .A3(new_n519), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n298), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n551), .A2(new_n334), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G200), .B2(new_n551), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n535), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  MUX2_X1   g0365(.A(G238), .B(G244), .S(G1698), .Z(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n303), .A3(new_n277), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n320), .B1(new_n567), .B2(new_n514), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n538), .A2(new_n539), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n315), .B(G250), .C1(G1), .C2(new_n327), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G179), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n572), .B2(new_n493), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n484), .A2(new_n264), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n303), .A2(new_n230), .A3(G68), .A4(new_n277), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT85), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n579));
  AOI21_X1  g0379(.A(G20), .B1(G33), .B2(G97), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT19), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OR3_X1    g0381(.A1(new_n413), .A2(KEYINPUT19), .A3(new_n215), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n576), .A2(new_n577), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n575), .B1(new_n584), .B2(new_n268), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n533), .A2(new_n482), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n586), .B(KEYINPUT86), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n533), .A2(new_n213), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n575), .B(new_n589), .C1(new_n584), .C2(new_n268), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n568), .A2(new_n334), .A3(new_n571), .ZN(new_n591));
  INV_X1    g0391(.A(new_n571), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n567), .A2(new_n514), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n320), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n591), .B1(G200), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n574), .A2(new_n588), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n303), .A2(G244), .A3(new_n378), .A4(new_n277), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT4), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(KEYINPUT4), .A2(G244), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n277), .A2(new_n279), .A3(new_n600), .A4(new_n378), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n277), .A2(new_n279), .A3(G250), .A4(G1698), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G283), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n377), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n543), .A2(new_n216), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n541), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n493), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n320), .B1(new_n599), .B2(new_n604), .ZN(new_n611));
  INV_X1    g0411(.A(new_n541), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n611), .A2(new_n612), .A3(new_n607), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n466), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n355), .A2(G107), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n471), .A2(KEYINPUT6), .A3(G97), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n215), .A2(new_n471), .ZN(new_n617));
  NOR2_X1   g0417(.A1(G97), .A2(G107), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(KEYINPUT6), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(G20), .B1(G77), .B2(new_n274), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n298), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n265), .A2(new_n215), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n533), .B2(new_n215), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n610), .B(new_n614), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n606), .A2(new_n334), .A3(new_n541), .A4(new_n608), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n613), .B2(G200), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n621), .B1(new_n294), .B2(new_n471), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n624), .B1(new_n628), .B2(new_n268), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n596), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT87), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT21), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n533), .A2(new_n509), .B1(new_n264), .B2(new_n513), .ZN(new_n634));
  AOI21_X1  g0434(.A(G20), .B1(G33), .B2(G283), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n276), .A2(G97), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n635), .A2(new_n636), .B1(new_n267), .B2(new_n229), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n510), .A2(new_n512), .A3(G20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n637), .A2(KEYINPUT20), .A3(new_n638), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n634), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT89), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI211_X1 g0445(.A(KEYINPUT89), .B(new_n634), .C1(new_n641), .C2(new_n642), .ZN(new_n646));
  OAI21_X1  g0446(.A(G169), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G270), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n541), .B1(new_n543), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n544), .A2(new_n378), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n303), .A2(new_n277), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT88), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n280), .A2(G303), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT88), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n303), .A2(new_n654), .A3(new_n277), .A4(new_n650), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n303), .A2(G257), .A3(new_n378), .A4(new_n277), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n652), .A2(new_n653), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n657), .B2(new_n377), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n633), .B1(new_n647), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n645), .A2(new_n646), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(G190), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n660), .B(new_n661), .C1(new_n336), .C2(new_n658), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n643), .B(new_n644), .ZN(new_n663));
  INV_X1    g0463(.A(new_n658), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT21), .A4(G169), .ZN(new_n665));
  AOI211_X1 g0465(.A(new_n466), .B(new_n649), .C1(new_n657), .C2(new_n377), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n659), .A2(new_n662), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT87), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n596), .A2(new_n625), .A3(new_n630), .A4(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n565), .A2(new_n632), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n501), .A2(new_n672), .ZN(G372));
  NAND2_X1  g0473(.A1(new_n350), .A2(new_n363), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n427), .A2(new_n428), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n426), .B1(new_n675), .B2(new_n497), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n676), .B2(new_n343), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n465), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n468), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n625), .A2(KEYINPUT92), .ZN(new_n681));
  INV_X1    g0481(.A(new_n629), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT92), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n610), .A4(new_n614), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n684), .A3(new_n596), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n588), .A2(new_n574), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n590), .A2(new_n595), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n690), .A2(new_n625), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n688), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n631), .A2(new_n564), .ZN(new_n696));
  INV_X1    g0496(.A(new_n551), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n552), .B(new_n553), .C1(new_n466), .C2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n559), .B2(new_n563), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n659), .A3(new_n667), .A4(new_n665), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n695), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n680), .B1(new_n501), .B2(new_n703), .ZN(G369));
  NAND3_X1  g0504(.A1(new_n659), .A2(new_n665), .A3(new_n667), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n263), .A2(new_n230), .A3(G13), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G213), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G343), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n660), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n668), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT94), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n716), .B(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n711), .B1(new_n559), .B2(new_n563), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n565), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n699), .B2(new_n712), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n556), .A2(new_n712), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n705), .A2(new_n712), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n565), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n233), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n579), .A2(new_n509), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n728), .A2(new_n263), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n228), .B2(new_n728), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT28), .Z(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n702), .A2(new_n733), .A3(new_n712), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n691), .B1(new_n690), .B2(new_n625), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n685), .B2(new_n686), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n711), .B1(new_n701), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n734), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n556), .A2(new_n668), .A3(new_n564), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(new_n632), .A3(new_n671), .A4(new_n712), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT95), .B1(new_n613), .B2(new_n551), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT95), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n609), .A2(new_n743), .A3(new_n697), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n658), .A2(G179), .A3(new_n572), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT96), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n611), .A2(new_n607), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n749), .A2(new_n551), .A3(new_n572), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n658), .A2(G179), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n551), .A2(new_n572), .A3(new_n751), .ZN(new_n755));
  INV_X1    g0555(.A(new_n748), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n666), .A3(new_n749), .A4(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n746), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n711), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT31), .B1(new_n758), .B2(new_n711), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n739), .B1(new_n741), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n738), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n732), .B1(new_n763), .B2(G1), .ZN(G364));
  INV_X1    g0564(.A(new_n728), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n230), .A2(G13), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n263), .B1(new_n766), .B2(G45), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n229), .B1(G20), .B2(new_n493), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n230), .A2(new_n466), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n772), .A2(new_n334), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n230), .A2(G179), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n336), .A2(G190), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n334), .A2(new_n336), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n777), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G179), .A2(G200), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G20), .A3(new_n334), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(G329), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n230), .B1(new_n785), .B2(G190), .ZN(new_n789));
  INV_X1    g0589(.A(G294), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n781), .A2(new_n771), .ZN(new_n791));
  INV_X1    g0591(.A(G326), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n280), .B1(new_n789), .B2(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n780), .A2(new_n784), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT98), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g0600(.A1(new_n771), .A2(KEYINPUT99), .A3(new_n778), .ZN(new_n801));
  AOI21_X1  g0601(.A(KEYINPUT99), .B1(new_n771), .B2(new_n778), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  OAI221_X1 g0604(.A(new_n794), .B1(new_n795), .B2(new_n800), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n791), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n773), .A2(G58), .B1(new_n806), .B2(G50), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n471), .B2(new_n779), .ZN(new_n808));
  INV_X1    g0608(.A(new_n803), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(G68), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n800), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G77), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n786), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT32), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n782), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n280), .B(new_n816), .C1(G87), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n789), .A2(new_n215), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n815), .B2(new_n814), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n810), .A2(new_n812), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n770), .B1(new_n805), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT97), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n769), .ZN(new_n828));
  INV_X1    g0628(.A(new_n309), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n233), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n327), .B2(new_n228), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n327), .B2(new_n256), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n233), .A2(G355), .A3(new_n445), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(G116), .C2(new_n233), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n768), .B(new_n822), .C1(new_n828), .C2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n715), .B2(new_n826), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n768), .B1(new_n715), .B2(G330), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n718), .B2(new_n837), .ZN(G396));
  OR2_X1    g0638(.A1(new_n496), .A2(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n496), .A2(KEYINPUT102), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n492), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n556), .A2(new_n705), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n528), .A2(new_n535), .A3(new_n561), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n844), .A2(new_n625), .A3(new_n630), .A4(new_n596), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n688), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n692), .B1(new_n685), .B2(new_n686), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n712), .B(new_n842), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT103), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n702), .A2(KEYINPUT103), .A3(new_n712), .A4(new_n842), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n488), .A2(new_n711), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n839), .A2(new_n491), .A3(new_n840), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n497), .A2(new_n711), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n702), .B2(new_n712), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  OR3_X1    g0659(.A1(new_n859), .A2(KEYINPUT104), .A3(new_n762), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT104), .B1(new_n859), .B2(new_n762), .ZN(new_n861));
  INV_X1    g0661(.A(new_n768), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n859), .B2(new_n762), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n770), .A2(new_n824), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n862), .B1(G77), .B2(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n774), .A2(new_n790), .B1(new_n791), .B2(new_n783), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n782), .A2(new_n471), .B1(new_n786), .B2(new_n795), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n280), .B1(new_n779), .B2(new_n213), .ZN(new_n869));
  NOR4_X1   g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n819), .ZN(new_n870));
  INV_X1    g0670(.A(new_n513), .ZN(new_n871));
  XNOR2_X1  g0671(.A(KEYINPUT100), .B(G283), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n870), .B1(new_n871), .B2(new_n800), .C1(new_n803), .C2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n773), .A2(G143), .B1(new_n806), .B2(G137), .ZN(new_n874));
  INV_X1    g0674(.A(G150), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n874), .B1(new_n875), .B2(new_n803), .C1(new_n800), .C2(new_n813), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT34), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n878));
  INV_X1    g0678(.A(new_n779), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G68), .ZN(new_n880));
  INV_X1    g0680(.A(G132), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n880), .B1(new_n202), .B2(new_n782), .C1(new_n881), .C2(new_n786), .ZN(new_n882));
  INV_X1    g0682(.A(new_n789), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n829), .B(new_n882), .C1(G58), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n873), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n866), .B1(new_n887), .B2(new_n769), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n857), .B2(new_n824), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n864), .A2(new_n889), .ZN(G384));
  OR2_X1    g0690(.A1(new_n620), .A2(KEYINPUT35), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n620), .A2(KEYINPUT35), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(G116), .A3(new_n231), .A4(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT36), .Z(new_n894));
  OR3_X1    g0694(.A1(new_n227), .A2(new_n414), .A3(new_n272), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n263), .B(G13), .C1(new_n895), .C2(new_n251), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n766), .A2(new_n263), .ZN(new_n898));
  INV_X1    g0698(.A(new_n709), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n361), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n342), .B(new_n900), .C1(new_n313), .C2(new_n349), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n351), .B1(new_n360), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n362), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n899), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n342), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(KEYINPUT38), .B(new_n909), .C1(new_n372), .C2(new_n906), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n901), .B(KEYINPUT37), .Z(new_n912));
  XNOR2_X1  g0712(.A(new_n342), .B(KEYINPUT17), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n900), .B1(new_n913), .B2(new_n674), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n911), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n367), .A2(new_n371), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n906), .B1(new_n919), .B2(new_n913), .ZN(new_n920));
  INV_X1    g0720(.A(new_n909), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n911), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n923));
  INV_X1    g0723(.A(new_n426), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(new_n711), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n918), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n674), .A2(new_n899), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n425), .A2(new_n712), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT105), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n675), .C1(new_n410), .C2(new_n425), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT105), .B(new_n675), .C1(new_n410), .C2(new_n425), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n410), .A2(new_n928), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n929), .A2(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n841), .A2(new_n712), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n852), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n922), .A2(new_n910), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n927), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n926), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n738), .A2(new_n500), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT106), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n738), .A2(new_n500), .A3(KEYINPUT106), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n679), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n940), .B(new_n945), .Z(new_n946));
  OAI21_X1  g0746(.A(new_n761), .B1(new_n672), .B2(new_n711), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n947), .A2(new_n934), .A3(new_n857), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n916), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n857), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n741), .B2(new_n761), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT107), .B1(new_n951), .B2(new_n934), .ZN(new_n952));
  OR2_X1    g0752(.A1(KEYINPUT107), .A2(KEYINPUT40), .ZN(new_n953));
  AND4_X1   g0753(.A1(new_n947), .A2(new_n934), .A3(new_n857), .A4(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n949), .A2(KEYINPUT40), .B1(new_n938), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n500), .A2(new_n947), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n959), .A2(new_n960), .A3(new_n739), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n898), .B1(new_n946), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT108), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n962), .A2(new_n963), .B1(new_n946), .B2(new_n961), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n897), .B1(new_n964), .B2(new_n965), .ZN(G367));
  OAI21_X1  g0766(.A(new_n828), .B1(new_n233), .B2(new_n482), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n830), .A2(new_n246), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n862), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(G143), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n774), .A2(new_n875), .B1(new_n791), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n789), .A2(new_n252), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n445), .B1(new_n779), .B2(new_n414), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n202), .B2(new_n800), .C1(new_n813), .C2(new_n803), .ZN(new_n975));
  INV_X1    g0775(.A(G137), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n782), .A2(new_n259), .B1(new_n786), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT113), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n795), .B2(new_n791), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(G303), .B2(new_n773), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n790), .B2(new_n803), .C1(new_n800), .C2(new_n872), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n779), .A2(new_n215), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n983), .B(new_n309), .C1(G317), .C2(new_n787), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n871), .A2(new_n782), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(KEYINPUT46), .B2(new_n985), .C1(new_n471), .C2(new_n789), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n975), .A2(new_n978), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n969), .B1(new_n988), .B2(new_n769), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n590), .A2(new_n712), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n695), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n690), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n989), .B1(new_n826), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n767), .B(KEYINPUT111), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n763), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT110), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n722), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n625), .A2(new_n712), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n625), .B(new_n630), .C1(new_n629), .C2(new_n712), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n725), .B2(new_n723), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT44), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT109), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(KEYINPUT109), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n718), .A2(KEYINPUT110), .A3(new_n721), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n725), .A2(new_n723), .A3(new_n1001), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT45), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n998), .A2(new_n1009), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1011), .B(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n997), .B(new_n722), .C1(new_n1008), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n716), .B(KEYINPUT94), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n725), .B1(new_n721), .B2(new_n724), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n996), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n996), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n728), .B(KEYINPUT41), .Z(new_n1023));
  OAI21_X1  g0823(.A(new_n995), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT112), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1001), .A2(new_n565), .A3(new_n724), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT42), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n625), .B1(new_n1000), .B2(new_n699), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1026), .A2(KEYINPUT42), .B1(new_n712), .B2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1027), .A2(new_n1029), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n718), .A2(new_n721), .A3(new_n1001), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1032), .B(new_n1033), .Z(new_n1034));
  AND3_X1   g0834(.A1(new_n1024), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1025), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n993), .B1(new_n1035), .B2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n1021), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n996), .A2(new_n1020), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n728), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n233), .A2(new_n445), .A3(new_n729), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n243), .A2(new_n327), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n830), .ZN(new_n1043));
  AOI211_X1 g0843(.A(G45), .B(new_n729), .C1(G68), .C2(G77), .ZN(new_n1044));
  OR3_X1    g0844(.A1(new_n261), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT50), .B1(new_n261), .B2(G50), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1043), .A2(new_n1047), .B1(new_n471), .B2(new_n727), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n828), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n862), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n773), .A2(G50), .B1(new_n806), .B2(G159), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n875), .B2(new_n786), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n811), .B2(G68), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n782), .A2(new_n414), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n789), .A2(new_n482), .ZN(new_n1055));
  NOR4_X1   g0855(.A1(new_n829), .A2(new_n1054), .A3(new_n983), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n809), .A2(new_n262), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1053), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n782), .A2(new_n790), .B1(new_n789), .B2(new_n872), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n773), .A2(G317), .B1(new_n806), .B2(G322), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n795), .B2(new_n803), .C1(new_n800), .C2(new_n783), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n871), .A2(new_n779), .B1(new_n792), .B2(new_n786), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1067), .A2(new_n309), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1058), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT114), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n770), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1050), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n721), .B2(new_n826), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1040), .B(new_n1075), .C1(new_n1020), .C2(new_n995), .ZN(G393));
  AOI21_X1  g0876(.A(new_n765), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1021), .B2(new_n1017), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n999), .A2(new_n1000), .A3(new_n827), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n828), .B1(new_n215), .B2(new_n233), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n830), .A2(new_n250), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n862), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n811), .A2(G294), .B1(G303), .B2(new_n809), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n773), .A2(G311), .B1(new_n806), .B2(G317), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT52), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n280), .B1(new_n779), .B2(new_n471), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n782), .A2(new_n872), .B1(new_n786), .B2(new_n775), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n513), .C2(new_n883), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1083), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n811), .A2(new_n479), .B1(G50), .B2(new_n809), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT115), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n773), .A2(G159), .B1(new_n806), .B2(G150), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  AOI22_X1  g0893(.A1(G68), .A2(new_n817), .B1(new_n879), .B2(G87), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n970), .B2(new_n786), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n789), .A2(new_n414), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1095), .A2(new_n829), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1091), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1090), .A2(KEYINPUT115), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1089), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1082), .B1(new_n1100), .B2(new_n769), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1017), .A2(new_n994), .B1(new_n1079), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1078), .A2(new_n1102), .ZN(G390));
  INV_X1    g0903(.A(G128), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n791), .A2(new_n1104), .B1(new_n779), .B2(new_n202), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G125), .B2(new_n787), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT117), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1106), .B1(new_n976), .B2(new_n803), .C1(new_n800), .C2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n782), .A2(new_n875), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n280), .B1(new_n773), .B2(G132), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(new_n813), .C2(new_n789), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n445), .B(new_n1096), .C1(G87), .C2(new_n817), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n787), .A2(G294), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n773), .A2(G116), .B1(new_n806), .B2(G283), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1114), .A2(new_n880), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n800), .A2(new_n215), .B1(new_n471), .B2(new_n803), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1109), .A2(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n770), .B1(new_n1119), .B2(KEYINPUT118), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(KEYINPUT118), .B2(new_n1119), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n862), .C1(new_n262), .C2(new_n865), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n918), .A2(new_n923), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n823), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n762), .A2(new_n857), .A3(new_n934), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT116), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1126), .A2(KEYINPUT116), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n925), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n852), .A2(new_n936), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n934), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1129), .A2(new_n1131), .B1(new_n918), .B2(new_n923), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n936), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n737), .B2(new_n842), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1134), .A2(new_n935), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n925), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n916), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1127), .B(new_n1128), .C1(new_n1132), .C2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT39), .B1(new_n910), .B2(new_n915), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1140), .A2(new_n1141), .B1(new_n925), .B2(new_n937), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1142), .A2(KEYINPUT116), .A3(new_n1126), .A4(new_n1137), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1124), .B1(new_n1144), .B2(new_n994), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n947), .A2(G330), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n935), .B1(new_n1146), .B2(new_n950), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n1125), .A3(new_n1134), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1147), .A2(new_n1125), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1133), .B1(new_n850), .B2(new_n851), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n500), .A2(new_n762), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n945), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n728), .B1(new_n1144), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1145), .B1(new_n1155), .B2(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(KEYINPUT120), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n944), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT106), .B1(new_n738), .B2(new_n500), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n680), .B(new_n1152), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n459), .A2(new_n463), .A3(new_n468), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n436), .A2(new_n709), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n956), .B2(new_n739), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1166), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n938), .A2(new_n955), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT40), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n916), .B2(new_n948), .ZN(new_n1171));
  OAI211_X1 g0971(.A(G330), .B(new_n1168), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1167), .A2(new_n940), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n940), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1156), .A2(new_n1161), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1158), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n765), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1161), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1174), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1167), .A2(new_n940), .A3(new_n1172), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1177), .A2(new_n1178), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n309), .A2(G41), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G33), .A2(G41), .ZN(new_n1188));
  OR3_X1    g0988(.A1(new_n1187), .A2(G50), .A3(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1187), .B1(new_n215), .B2(new_n803), .C1(new_n800), .C2(new_n482), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n879), .A2(G58), .B1(new_n787), .B2(G283), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n509), .B2(new_n791), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n774), .A2(new_n471), .B1(new_n414), .B2(new_n782), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1190), .A2(new_n972), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1189), .B1(new_n1194), .B2(KEYINPUT58), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT119), .Z(new_n1196));
  AOI22_X1  g0996(.A1(new_n773), .A2(G128), .B1(new_n806), .B2(G125), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n875), .B2(new_n789), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n811), .B2(G137), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n881), .B2(new_n803), .C1(new_n782), .C2(new_n1108), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  INV_X1    g1001(.A(G124), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1188), .B1(new_n786), .B2(new_n1202), .C1(new_n779), .C2(new_n813), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1200), .B2(KEYINPUT59), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1201), .A2(new_n1204), .B1(KEYINPUT58), .B2(new_n1194), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n770), .B1(new_n1196), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n862), .B1(G50), .B2(new_n865), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n1166), .C2(new_n823), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1184), .B2(new_n994), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1186), .A2(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n1151), .A2(new_n994), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n862), .B1(G68), .B2(new_n865), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n774), .A2(new_n776), .B1(new_n791), .B2(new_n790), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n782), .A2(new_n215), .B1(new_n786), .B2(new_n783), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n280), .B1(new_n779), .B2(new_n414), .ZN(new_n1215));
  OR4_X1    g1015(.A1(new_n1055), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n800), .A2(new_n471), .B1(new_n871), .B2(new_n803), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n806), .A2(G132), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT121), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n803), .B2(new_n1108), .C1(new_n800), .C2(new_n875), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n829), .B1(G50), .B2(new_n883), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n879), .A2(G58), .B1(new_n787), .B2(G128), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n773), .A2(G137), .B1(G159), .B2(new_n817), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n1216), .A2(new_n1217), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1212), .B1(new_n1225), .B2(new_n769), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n934), .B2(new_n824), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1211), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1154), .A2(new_n1023), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1151), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1161), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1229), .B1(new_n1230), .B2(new_n1233), .ZN(G381));
  OR2_X1    g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  OR4_X1    g1035(.A1(G384), .A2(G381), .A3(new_n1235), .A4(G390), .ZN(new_n1236));
  OR4_X1    g1036(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1236), .ZN(G407));
  INV_X1    g1037(.A(G378), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n710), .A2(G213), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G375), .C2(new_n1241), .ZN(G409));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  INV_X1    g1043(.A(G390), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n993), .B(G390), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  XOR2_X1   g1047(.A(G393), .B(G396), .Z(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1248), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1024), .A2(new_n1034), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT112), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1024), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G390), .B1(new_n1254), .B2(new_n993), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1250), .B1(new_n1255), .B2(KEYINPUT125), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G387), .A2(KEYINPUT125), .A3(new_n1244), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1246), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1254), .A2(KEYINPUT126), .A3(new_n993), .A4(G390), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1249), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1186), .A2(G378), .A3(new_n1209), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1209), .B1(new_n1023), .B2(new_n1175), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1238), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1240), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1231), .A2(new_n1161), .A3(KEYINPUT60), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(new_n728), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1232), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1267), .B1(new_n1272), .B2(new_n1228), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1228), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(G384), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(G2897), .A3(new_n1240), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1274), .B(new_n1267), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT123), .ZN(new_n1279));
  INV_X1    g1079(.A(G2897), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1239), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT124), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1283));
  AND4_X1   g1083(.A1(KEYINPUT124), .A2(new_n1273), .A3(new_n1275), .A4(new_n1282), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1277), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1243), .B(new_n1262), .C1(new_n1266), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1240), .B(new_n1276), .C1(new_n1263), .C2(new_n1265), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT63), .B1(new_n1288), .B2(KEYINPUT122), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1266), .A2(new_n1278), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT122), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1287), .A2(new_n1289), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1266), .A2(new_n1295), .A3(new_n1278), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1243), .B1(new_n1266), .B2(new_n1285), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1266), .B2(new_n1278), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1294), .B1(new_n1299), .B2(new_n1262), .ZN(G405));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1238), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1263), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1301), .A2(KEYINPUT127), .A3(new_n1263), .A4(new_n1278), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1262), .ZN(G402));
endmodule


