//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT72), .A3(G128), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT24), .B(G110), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT73), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n193), .B2(G119), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n195), .A2(new_n197), .A3(new_n198), .A4(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n194), .A3(new_n192), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT73), .B1(new_n202), .B2(new_n196), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n191), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n194), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(KEYINPUT23), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n201), .A2(new_n203), .B1(G110), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT74), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT74), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G125), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(G125), .A2(G140), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT16), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n213), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n209), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n216), .A2(G146), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(G146), .B1(new_n216), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n208), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(G146), .A3(new_n219), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT65), .A2(G146), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT65), .A2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n210), .A2(new_n209), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n215), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n207), .A2(G110), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n202), .A2(new_n196), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n223), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n233), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n222), .A2(new_n231), .A3(new_n236), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n188), .A3(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n241), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n238), .A2(new_n188), .A3(new_n239), .A4(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n190), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n239), .ZN(new_n246));
  NOR3_X1   g060(.A1(new_n246), .A2(G902), .A3(new_n189), .ZN(new_n247));
  OR2_X1    g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n249));
  INV_X1    g063(.A(G237), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n234), .A3(G210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n249), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(G116), .B(G119), .Z(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OR2_X1    g072(.A1(KEYINPUT64), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT64), .A2(G143), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(G146), .A3(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(KEYINPUT65), .A2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT65), .A2(G146), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(G143), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n261), .A2(new_n264), .A3(new_n265), .A4(G128), .ZN(new_n266));
  AOI21_X1  g080(.A(G146), .B1(new_n259), .B2(new_n260), .ZN(new_n267));
  AOI21_X1  g081(.A(G143), .B1(new_n262), .B2(new_n263), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n193), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G134), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT66), .B1(new_n272), .B2(G137), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT11), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G134), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT11), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT66), .B(new_n279), .C1(new_n272), .C2(G137), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n274), .A2(new_n275), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n272), .A2(G137), .ZN(new_n282));
  OAI21_X1  g096(.A(G131), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  NOR2_X1   g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n267), .B2(new_n268), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n261), .A2(new_n264), .A3(new_n286), .ZN(new_n290));
  INV_X1    g104(.A(new_n281), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n277), .B1(new_n273), .B2(KEYINPUT11), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n275), .B1(new_n292), .B2(new_n280), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n289), .B(new_n290), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT30), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n285), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n258), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n285), .A2(new_n294), .A3(new_n258), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n285), .A2(new_n294), .A3(new_n302), .A4(new_n258), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n254), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n301), .B2(new_n303), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n300), .A2(new_n308), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n295), .A2(new_n257), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n309), .A2(new_n312), .A3(new_n254), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n188), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n292), .A2(new_n280), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G131), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n281), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n289), .A2(new_n290), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n318), .A2(new_n319), .B1(new_n271), .B2(new_n284), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n302), .B1(new_n320), .B2(new_n258), .ZN(new_n321));
  INV_X1    g135(.A(new_n303), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n301), .A2(KEYINPUT70), .A3(new_n303), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n308), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n254), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT29), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n325), .A2(new_n312), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G472), .B1(new_n314), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n254), .B1(new_n309), .B2(new_n312), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n321), .A2(new_n322), .ZN(new_n331));
  INV_X1    g145(.A(new_n298), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n297), .B1(new_n285), .B2(new_n294), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n257), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n331), .A2(new_n334), .A3(new_n326), .A4(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n299), .A2(new_n304), .A3(new_n254), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT31), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n330), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT32), .ZN(new_n340));
  NOR2_X1   g154(.A1(G472), .A2(G902), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n339), .B2(new_n341), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n329), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT71), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT71), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n329), .B(new_n346), .C1(new_n342), .C2(new_n343), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n248), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G110), .B(G140), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n234), .A2(G227), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n354));
  INV_X1    g168(.A(G107), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n355), .A2(G104), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT3), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n354), .A2(new_n361), .A3(new_n355), .A4(G104), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n353), .B(G101), .C1(new_n360), .C2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n289), .A3(new_n290), .ZN(new_n365));
  INV_X1    g179(.A(G101), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n357), .A2(new_n366), .A3(new_n362), .A4(new_n359), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT4), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n358), .B1(new_n356), .B2(KEYINPUT3), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n369), .B2(new_n362), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n352), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G101), .B1(new_n360), .B2(new_n363), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(new_n319), .A3(KEYINPUT77), .A4(new_n364), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G128), .B1(new_n267), .B2(new_n265), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n261), .A2(new_n264), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n266), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G107), .ZN(new_n382));
  OAI21_X1  g196(.A(G101), .B1(new_n382), .B2(new_n358), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n367), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n265), .B1(new_n226), .B2(G143), .ZN(new_n387));
  OAI22_X1  g201(.A1(new_n387), .A2(new_n193), .B1(new_n267), .B2(new_n268), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(new_n266), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n385), .A2(new_n386), .B1(new_n389), .B2(new_n384), .ZN(new_n390));
  INV_X1    g204(.A(new_n318), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n376), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n376), .B2(new_n390), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n351), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n271), .A2(new_n384), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n367), .A2(new_n383), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n379), .B2(new_n266), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n318), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT12), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(new_n398), .A3(new_n266), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n385), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(KEYINPUT78), .A3(KEYINPUT12), .A4(new_n318), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n401), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n351), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n392), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n395), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G469), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n188), .ZN(new_n412));
  INV_X1    g226(.A(new_n407), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n351), .B1(new_n413), .B2(new_n393), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n392), .A2(new_n408), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n376), .A2(new_n390), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n318), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(G469), .A3(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n411), .A2(new_n188), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n412), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT9), .B(G234), .ZN(new_n423));
  OAI21_X1  g237(.A(G221), .B1(new_n423), .B2(G902), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT13), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n259), .A2(new_n427), .A3(G128), .A4(new_n260), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n193), .A2(G143), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n259), .A2(new_n260), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(new_n193), .ZN(new_n431));
  OAI211_X1 g245(.A(G134), .B(new_n428), .C1(new_n431), .C2(new_n427), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G116), .ZN(new_n434));
  INV_X1    g248(.A(G116), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(G122), .ZN(new_n436));
  OAI21_X1  g250(.A(G107), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(G122), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(G116), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n355), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT82), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n272), .B(new_n429), .C1(new_n430), .C2(new_n193), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n437), .A2(new_n444), .A3(new_n440), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n432), .A2(new_n442), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n431), .A2(G134), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n443), .ZN(new_n448));
  INV_X1    g262(.A(new_n440), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n438), .B1(new_n436), .B2(KEYINPUT14), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT14), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n434), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n438), .B2(KEYINPUT14), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n449), .B1(new_n455), .B2(G107), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n423), .A2(new_n187), .A3(G953), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n446), .A2(new_n457), .A3(new_n459), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(KEYINPUT84), .A3(new_n460), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n188), .A4(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n467), .A2(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n426), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n467), .A2(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n467), .A2(new_n469), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(KEYINPUT86), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n250), .A2(new_n234), .A3(G143), .A4(G214), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n250), .A2(new_n234), .A3(G214), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(new_n430), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT18), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(KEYINPUT80), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(G131), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n275), .B(new_n477), .C1(new_n430), .C2(new_n478), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n485), .B2(new_n481), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT81), .ZN(new_n487));
  INV_X1    g301(.A(new_n215), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n211), .A2(new_n213), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n209), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT81), .B1(new_n214), .B2(new_n215), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(G146), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n228), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n381), .ZN(new_n496));
  INV_X1    g310(.A(new_n221), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n483), .A2(new_n498), .A3(new_n484), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n479), .A2(KEYINPUT17), .A3(G131), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n223), .A4(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n496), .B1(new_n494), .B2(new_n501), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n188), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G475), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT19), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n490), .B2(new_n491), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n227), .A2(KEYINPUT19), .A3(new_n215), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n226), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n485), .A2(new_n223), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n510), .A2(new_n511), .B1(new_n486), .B2(new_n493), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n502), .B1(new_n512), .B2(new_n496), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n506), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n234), .A2(G952), .ZN(new_n520));
  INV_X1    g334(.A(G234), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(new_n521), .B2(new_n250), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n188), .B(new_n234), .C1(G234), .C2(G237), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT21), .B(G898), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n476), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G224), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G953), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n217), .B1(new_n388), .B2(new_n266), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n289), .A2(new_n290), .A3(new_n217), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT7), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n533), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n271), .A2(new_n489), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n364), .B(new_n257), .C1(new_n368), .C2(new_n370), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n255), .A2(new_n256), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT5), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n191), .A3(G116), .ZN(new_n542));
  OAI211_X1 g356(.A(G113), .B(new_n542), .C1(new_n255), .C2(new_n541), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n384), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(G110), .B(G122), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n539), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(KEYINPUT8), .ZN(new_n547));
  AND4_X1   g361(.A1(new_n540), .A2(new_n543), .A3(new_n367), .A4(new_n383), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n543), .A2(new_n540), .B1(new_n367), .B2(new_n383), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n534), .A2(new_n538), .A3(new_n546), .A4(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n551), .A2(new_n188), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n539), .A2(new_n544), .ZN(new_n553));
  INV_X1    g367(.A(new_n545), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n532), .A2(new_n530), .A3(new_n533), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT6), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n553), .A2(new_n560), .A3(new_n554), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n552), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G210), .B1(G237), .B2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n552), .A2(new_n562), .A3(new_n564), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(KEYINPUT79), .A3(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n567), .A2(KEYINPUT79), .ZN(new_n569));
  OAI21_X1  g383(.A(G214), .B1(G237), .B2(G902), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n425), .A2(new_n528), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n348), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT87), .B(G101), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(G3));
  INV_X1    g389(.A(G472), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n339), .B2(new_n188), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n339), .A2(new_n341), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n425), .A2(new_n580), .A3(new_n248), .ZN(new_n581));
  INV_X1    g395(.A(new_n570), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n566), .B2(new_n567), .ZN(new_n583));
  INV_X1    g397(.A(new_n526), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n464), .A2(new_n586), .A3(new_n466), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n461), .A2(KEYINPUT33), .A3(new_n463), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n188), .A2(G478), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n464), .A2(new_n188), .A3(new_n466), .ZN(new_n591));
  OAI22_X1  g405(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(G478), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n519), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n581), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT34), .B(G104), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G6));
  NAND2_X1  g413(.A1(new_n513), .A2(new_n515), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT20), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n601), .A2(new_n516), .B1(G475), .B2(new_n505), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n472), .A2(new_n475), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n603), .A2(KEYINPUT90), .A3(new_n584), .A4(new_n583), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT90), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n472), .A2(new_n475), .A3(new_n602), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n605), .B1(new_n606), .B2(new_n585), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n581), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G107), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  NOR2_X1   g425(.A1(new_n237), .A2(KEYINPUT36), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n232), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n222), .A2(new_n231), .A3(new_n612), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n614), .A2(new_n188), .A3(new_n190), .A4(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT91), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT92), .B1(new_n618), .B2(new_n245), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n242), .A2(new_n244), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n189), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n616), .B(KEYINPUT91), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  OR3_X1    g439(.A1(new_n580), .A2(KEYINPUT93), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT93), .B1(new_n580), .B2(new_n625), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n572), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT37), .B(G110), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  INV_X1    g444(.A(KEYINPUT94), .ZN(new_n631));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n523), .B1(new_n524), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n603), .A2(new_n631), .A3(new_n583), .A4(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n472), .A2(new_n475), .A3(new_n602), .A4(new_n634), .ZN(new_n636));
  INV_X1    g450(.A(new_n583), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT94), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n345), .A2(new_n347), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n422), .A2(new_n424), .A3(new_n619), .A4(new_n624), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  NAND2_X1  g458(.A1(new_n579), .A2(KEYINPUT32), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n331), .A2(new_n334), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n326), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n188), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n311), .A2(new_n323), .A3(new_n254), .A4(new_n324), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT96), .ZN(new_n654));
  INV_X1    g468(.A(new_n568), .ZN(new_n655));
  INV_X1    g469(.A(new_n569), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n476), .A2(new_n602), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n621), .A2(new_n622), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n570), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n654), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n424), .ZN(new_n665));
  AOI21_X1  g479(.A(G902), .B1(new_n395), .B2(new_n409), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n420), .B1(new_n666), .B2(new_n411), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n665), .B1(new_n667), .B2(new_n419), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT97), .B(KEYINPUT39), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n633), .B(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT40), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n430), .ZN(G45));
  NOR3_X1   g488(.A1(new_n637), .A2(new_n593), .A3(new_n633), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n640), .A2(new_n642), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  AOI21_X1  g491(.A(new_n411), .B1(new_n410), .B2(new_n188), .ZN(new_n678));
  AOI211_X1 g492(.A(G469), .B(G902), .C1(new_n395), .C2(new_n409), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n424), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n417), .A2(new_n392), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n351), .A2(new_n683), .B1(new_n415), .B2(new_n407), .ZN(new_n684));
  OAI21_X1  g498(.A(G469), .B1(new_n684), .B2(G902), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n424), .A3(new_n412), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n348), .A2(new_n688), .A3(new_n594), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND3_X1  g505(.A1(new_n348), .A2(new_n688), .A3(new_n608), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NAND4_X1  g507(.A1(new_n476), .A2(new_n527), .A3(new_n619), .A4(new_n624), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n685), .A2(new_n424), .A3(new_n583), .A4(new_n412), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n346), .B1(new_n647), .B2(new_n329), .ZN(new_n697));
  INV_X1    g511(.A(new_n347), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  INV_X1    g514(.A(new_n341), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT99), .B1(new_n325), .B2(new_n312), .ZN(new_n702));
  INV_X1    g516(.A(new_n324), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT70), .B1(new_n301), .B2(new_n303), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT28), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT99), .ZN(new_n706));
  INV_X1    g520(.A(new_n312), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n702), .A2(new_n708), .A3(new_n254), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT31), .B1(new_n648), .B2(new_n254), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n336), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n701), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n713), .A2(new_n248), .A3(new_n577), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n583), .A2(new_n472), .A3(new_n475), .A4(new_n519), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n526), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n714), .A2(new_n687), .A3(new_n682), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  NOR2_X1   g532(.A1(new_n325), .A2(new_n312), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n326), .B1(new_n719), .B2(new_n706), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n711), .B1(new_n720), .B2(new_n702), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n578), .B(new_n661), .C1(new_n721), .C2(new_n701), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n519), .A2(new_n592), .A3(new_n634), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n680), .A2(new_n424), .A3(new_n723), .A4(new_n583), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n210), .ZN(G27));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n647), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n645), .A2(KEYINPUT101), .A3(new_n646), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n329), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n248), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n582), .B1(new_n568), .B2(new_n569), .ZN(new_n732));
  AND4_X1   g546(.A1(new_n424), .A2(new_n732), .A3(new_n422), .A4(new_n723), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n640), .A2(KEYINPUT100), .A3(new_n731), .A4(new_n733), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT100), .B1(new_n348), .B2(new_n733), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(KEYINPUT102), .B(new_n734), .C1(new_n737), .C2(new_n738), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n275), .ZN(G33));
  INV_X1    g558(.A(new_n636), .ZN(new_n745));
  INV_X1    g559(.A(new_n732), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n425), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n348), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND2_X1  g563(.A1(new_n602), .A2(new_n592), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT43), .Z(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT103), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n750), .B(KEYINPUT43), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n662), .B1(new_n578), .B2(new_n579), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n755), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n732), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(KEYINPUT105), .B(new_n732), .C1(new_n760), .C2(new_n761), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n760), .A2(new_n761), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n414), .A2(new_n418), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n414), .A2(KEYINPUT45), .A3(new_n418), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT46), .B1(new_n772), .B2(new_n421), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n679), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n421), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n665), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n670), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n767), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n766), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  NAND3_X1  g594(.A1(new_n732), .A2(new_n723), .A3(new_n248), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n640), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT106), .B(G140), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G42));
  NOR2_X1   g600(.A1(new_n753), .A2(new_n522), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(new_n714), .ZN(new_n788));
  INV_X1    g602(.A(new_n686), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(KEYINPUT112), .A3(new_n582), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n686), .B2(new_n570), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n788), .A2(new_n659), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT50), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n753), .A2(new_n746), .A3(new_n522), .A4(new_n686), .ZN(new_n795));
  INV_X1    g609(.A(new_n722), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n746), .A2(new_n686), .A3(new_n248), .A4(new_n522), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n654), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n519), .A3(new_n592), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n794), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n680), .A2(KEYINPUT111), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n680), .A2(KEYINPUT111), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n665), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n782), .A2(new_n783), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n732), .A3(new_n788), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n730), .A2(new_n731), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n795), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT48), .Z(new_n810));
  OR2_X1    g624(.A1(new_n799), .A2(new_n593), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n788), .A2(new_n583), .A3(new_n789), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n520), .A3(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n807), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n742), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n733), .B(new_n731), .C1(new_n697), .C2(new_n698), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT100), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n736), .A3(new_n735), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT102), .B1(new_n819), .B2(new_n734), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n713), .A2(new_n593), .A3(new_n577), .A4(new_n662), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n473), .A2(new_n474), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n625), .A2(new_n823), .A3(new_n519), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n640), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n747), .A2(new_n634), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n748), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n602), .A2(new_n823), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n526), .B1(new_n828), .B2(new_n593), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n581), .A2(new_n570), .A3(new_n657), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n573), .A2(new_n830), .A3(new_n628), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT107), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n731), .B1(new_n697), .B2(new_n698), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n682), .A2(new_n687), .A3(new_n594), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n699), .B(new_n717), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n348), .A2(new_n608), .A3(new_n688), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n699), .A2(new_n717), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(KEYINPUT107), .A3(new_n689), .A4(new_n692), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n832), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n715), .B1(new_n647), .B2(new_n652), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n661), .A2(new_n633), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT108), .B1(new_n668), .B2(new_n843), .ZN(new_n844));
  AND4_X1   g658(.A1(KEYINPUT108), .A2(new_n422), .A3(new_n843), .A4(new_n424), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n722), .A2(new_n724), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n643), .A2(new_n676), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n641), .B1(new_n345), .B2(new_n347), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n725), .B1(new_n851), .B2(new_n639), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n676), .A4(new_n846), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT109), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT109), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n821), .A2(new_n841), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT53), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n832), .A2(new_n838), .A3(new_n840), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n743), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n854), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n859), .A2(KEYINPUT54), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n838), .A2(new_n840), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n741), .A3(new_n742), .A4(new_n832), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n857), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT110), .B1(new_n836), .B2(new_n837), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT110), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n839), .A2(new_n871), .A3(new_n689), .A4(new_n692), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n827), .A2(new_n831), .A3(new_n862), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n739), .A2(new_n873), .A3(new_n854), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n868), .A2(new_n869), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n788), .A2(new_n732), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n805), .B2(KEYINPUT113), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(KEYINPUT113), .B2(new_n805), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n801), .A3(KEYINPUT51), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n814), .A2(new_n864), .A3(new_n877), .A4(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(G952), .B2(G953), .ZN(new_n883));
  INV_X1    g697(.A(new_n680), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n884), .A2(KEYINPUT49), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(KEYINPUT49), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n731), .A2(new_n424), .A3(new_n570), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n750), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n654), .A3(new_n659), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n883), .A2(new_n889), .ZN(G75));
  AOI21_X1  g704(.A(new_n875), .B1(new_n858), .B2(new_n862), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT114), .B1(new_n891), .B2(new_n188), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT114), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT109), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT109), .B1(new_n850), .B2(new_n853), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT53), .B1(new_n861), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n893), .B(G902), .C1(new_n897), .C2(new_n875), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n565), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n556), .A2(new_n561), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n559), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT116), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(KEYINPUT116), .ZN(new_n904));
  XOR2_X1   g718(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n899), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n234), .A2(G952), .ZN(new_n908));
  OAI211_X1 g722(.A(G210), .B(G902), .C1(new_n897), .C2(new_n875), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n911), .B2(new_n902), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n907), .A2(new_n912), .ZN(G51));
  OAI21_X1  g727(.A(KEYINPUT54), .B1(new_n897), .B2(new_n875), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n877), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n420), .B(KEYINPUT117), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT57), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n410), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n772), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n892), .A2(new_n920), .A3(new_n898), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n908), .B1(new_n919), .B2(new_n921), .ZN(G54));
  AND2_X1   g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n892), .A2(new_n898), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n513), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n908), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n892), .A2(new_n513), .A3(new_n898), .A4(new_n923), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G60));
  XNOR2_X1  g743(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n468), .A2(new_n188), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n930), .B(new_n931), .Z(new_n932));
  AOI21_X1  g746(.A(new_n862), .B1(new_n861), .B2(new_n896), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n854), .A2(new_n862), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n743), .A2(new_n934), .A3(new_n860), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n869), .A3(new_n935), .ZN(new_n936));
  AOI211_X1 g750(.A(KEYINPUT54), .B(new_n875), .C1(new_n858), .C2(new_n862), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n589), .B(KEYINPUT118), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n932), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n864), .B2(new_n877), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT120), .B1(new_n944), .B2(new_n940), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n941), .A2(new_n943), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n908), .B1(new_n915), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n942), .A2(new_n945), .A3(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n891), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n614), .A2(new_n615), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n246), .B1(new_n891), .B2(new_n950), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(new_n927), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n927), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(G66));
  INV_X1    g773(.A(new_n525), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n234), .B1(new_n960), .B2(G224), .ZN(new_n961));
  INV_X1    g775(.A(new_n831), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n865), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n961), .B1(new_n963), .B2(new_n234), .ZN(new_n964));
  INV_X1    g778(.A(G898), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n900), .B1(new_n965), .B2(G953), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G69));
  AND2_X1   g781(.A1(new_n852), .A2(new_n676), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n673), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n828), .A2(new_n593), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n348), .A2(new_n671), .A3(new_n732), .A4(new_n972), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT122), .Z(new_n974));
  NOR2_X1   g788(.A1(new_n784), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n971), .A2(new_n975), .A3(new_n779), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n234), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n332), .A2(new_n333), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n508), .A2(new_n509), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT121), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT123), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n983));
  INV_X1    g797(.A(new_n981), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n983), .B(new_n984), .C1(new_n976), .C2(new_n234), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n777), .B(new_n767), .C1(new_n764), .C2(new_n765), .ZN(new_n987));
  INV_X1    g801(.A(new_n968), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n808), .A2(new_n583), .A3(new_n660), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n748), .B1(new_n777), .B2(new_n990), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n743), .A2(new_n784), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n779), .A2(KEYINPUT124), .A3(new_n968), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n234), .A2(new_n989), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n980), .B1(new_n632), .B2(new_n234), .ZN(new_n995));
  OAI22_X1  g809(.A1(new_n982), .A2(new_n985), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n234), .B1(G227), .B2(G900), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n997), .ZN(new_n999));
  OAI221_X1 g813(.A(new_n999), .B1(new_n994), .B2(new_n995), .C1(new_n982), .C2(new_n985), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(G72));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT125), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n976), .B2(new_n963), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(new_n326), .A3(new_n648), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n648), .A2(new_n326), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1008), .A2(new_n649), .A3(new_n1003), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT127), .Z(new_n1010));
  NAND3_X1  g824(.A1(new_n859), .A2(new_n863), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n963), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n989), .A2(new_n992), .A3(new_n1013), .A4(new_n993), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1008), .B1(new_n1014), .B2(new_n1004), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n1015), .A2(KEYINPUT126), .A3(new_n908), .ZN(new_n1016));
  OAI21_X1  g830(.A(KEYINPUT126), .B1(new_n1015), .B2(new_n908), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(G57));
endmodule


