//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n203), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT73), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT73), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n207), .B2(new_n209), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT74), .B(G141gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n203), .B1(new_n218), .B2(G148gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n207), .B1(new_n206), .B2(new_n209), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n219), .A2(KEYINPUT75), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT75), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT74), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G141gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n225), .A3(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n203), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n211), .B1(new_n210), .B2(KEYINPUT2), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n222), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n215), .B(new_n217), .C1(new_n221), .C2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G197gat), .A2(G204gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G211gat), .ZN(new_n239));
  INV_X1    g038(.A(G218gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G211gat), .A2(G218gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(KEYINPUT71), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n238), .A2(new_n243), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n233), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G228gat), .ZN(new_n248));
  INV_X1    g047(.A(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252));
  AND2_X1   g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(new_n235), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n254), .B2(new_n234), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n241), .A2(new_n242), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT22), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(KEYINPUT82), .C1(new_n235), .C2(new_n253), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n255), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n242), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n252), .B(new_n261), .C1(new_n254), .C2(new_n234), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n232), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n217), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n215), .B1(new_n221), .B2(new_n230), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n262), .A2(new_n232), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n255), .A2(new_n242), .A3(new_n241), .A4(new_n259), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n216), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n208), .A2(new_n212), .A3(new_n214), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT75), .B1(new_n219), .B2(new_n220), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n228), .A2(new_n222), .A3(new_n229), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT83), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n247), .A2(new_n251), .A3(new_n267), .A4(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n246), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n277), .B1(new_n231), .B2(new_n232), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n273), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n232), .B1(new_n244), .B2(new_n245), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n215), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n250), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G78gat), .B(G106gat), .ZN(new_n284));
  INV_X1    g083(.A(G50gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n286), .B(KEYINPUT81), .Z(new_n287));
  AND3_X1   g086(.A1(new_n276), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n276), .B2(new_n283), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n290), .B(G22gat), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT29), .B1(new_n274), .B2(new_n217), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n251), .B1(new_n294), .B2(new_n277), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n267), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n283), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n287), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n276), .A2(new_n283), .A3(new_n287), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n291), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT26), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(new_n303), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G183gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT27), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G183gat), .ZN(new_n315));
  INV_X1    g114(.A(G190gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n318), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT27), .B(G183gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(new_n316), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n311), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n305), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT64), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n307), .B1(new_n303), .B2(KEYINPUT23), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n332), .A2(G169gat), .A3(G176gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT65), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n303), .A2(KEYINPUT23), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n332), .B1(G169gat), .B2(G176gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT65), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n335), .A2(new_n307), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n330), .A2(new_n334), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n307), .A3(new_n336), .ZN(new_n341));
  AND2_X1   g140(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n305), .A2(new_n324), .B1(new_n342), .B2(G190gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT25), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n323), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  OAI22_X1  g144(.A1(KEYINPUT70), .A2(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(KEYINPUT70), .B2(KEYINPUT1), .ZN(new_n347));
  NAND2_X1  g146(.A1(G127gat), .A2(G134gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(G127gat), .A2(G134gat), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT69), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n350), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT69), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n348), .ZN(new_n354));
  AND2_X1   g153(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n356));
  OAI21_X1  g155(.A(G120gat), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n347), .A2(new_n351), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT67), .ZN(new_n359));
  NAND2_X1  g158(.A1(G113gat), .A2(G120gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(G113gat), .A2(G120gat), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT1), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n352), .A2(new_n348), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n359), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n362), .A2(KEYINPUT1), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n360), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n367), .A2(KEYINPUT67), .A3(new_n352), .A4(new_n348), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n358), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n345), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G227gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(new_n249), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n358), .A2(new_n365), .A3(new_n368), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n373), .A2(new_n323), .A3(new_n340), .A4(new_n344), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT32), .ZN(new_n376));
  XOR2_X1   g175(.A(G15gat), .B(G43gat), .Z(new_n377));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT34), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n370), .A2(new_n374), .ZN(new_n384));
  INV_X1    g183(.A(new_n372), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g185(.A(KEYINPUT34), .B(new_n372), .C1(new_n370), .C2(new_n374), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n382), .A2(new_n386), .A3(new_n387), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n376), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n381), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n379), .ZN(new_n393));
  INV_X1    g192(.A(new_n387), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n384), .A2(new_n385), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT34), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n376), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n388), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n302), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT5), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n266), .A2(new_n373), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n274), .A2(new_n369), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n406), .B(KEYINPUT77), .Z(new_n407));
  AOI21_X1  g206(.A(new_n402), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n231), .B(new_n373), .C1(new_n274), .C2(new_n281), .ZN(new_n409));
  INV_X1    g208(.A(new_n407), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n266), .B2(new_n373), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n274), .A2(new_n369), .A3(KEYINPUT4), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n409), .A2(new_n410), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n266), .A2(new_n411), .A3(new_n373), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT4), .B1(new_n274), .B2(new_n369), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n418), .A2(new_n402), .A3(new_n410), .A4(new_n409), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(G1gat), .B(G29gat), .Z(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n415), .A2(new_n419), .A3(new_n425), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n420), .A2(new_n426), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n428), .B2(new_n430), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n427), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G226gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n345), .B2(new_n232), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n317), .A2(new_n318), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n321), .A2(new_n316), .A3(new_n320), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n331), .A2(new_n333), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n325), .A2(new_n326), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n441), .A2(new_n311), .B1(new_n444), .B2(KEYINPUT25), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n436), .B1(new_n445), .B2(new_n340), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n438), .A2(new_n446), .A3(new_n246), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G8gat), .B(G36gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT72), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n345), .A2(new_n232), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n436), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n345), .A2(new_n437), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT29), .B1(new_n445), .B2(new_n340), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n437), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n460), .B2(new_n455), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n448), .B(new_n454), .C1(new_n461), .C2(new_n277), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n455), .B1(new_n438), .B2(new_n446), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT72), .B1(new_n459), .B2(new_n437), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n277), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n452), .B1(new_n465), .B2(new_n447), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n464), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n447), .B1(new_n468), .B2(new_n246), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT30), .B1(new_n469), .B2(new_n451), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n401), .A2(new_n435), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT84), .B1(new_n467), .B2(new_n470), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n448), .B(new_n451), .C1(new_n461), .C2(new_n277), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n453), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n462), .A4(new_n466), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n397), .A2(new_n398), .A3(new_n388), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n398), .B1(new_n397), .B2(new_n388), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n428), .A2(new_n430), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n425), .B(KEYINPUT85), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n415), .B2(new_n419), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n427), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n292), .B1(new_n288), .B2(new_n289), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n299), .A2(new_n291), .A3(new_n300), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n482), .A2(new_n486), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT88), .B1(new_n479), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g291(.A(new_n430), .B(new_n425), .C1(new_n415), .C2(new_n419), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n428), .A2(new_n430), .ZN(new_n494));
  INV_X1    g293(.A(new_n485), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(KEYINPUT35), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n474), .A2(new_n478), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n497), .A2(new_n401), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n473), .A2(new_n492), .A3(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n391), .A2(KEYINPUT36), .A3(new_n399), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT36), .B1(new_n391), .B2(new_n399), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n435), .A2(new_n471), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n302), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n452), .A2(KEYINPUT37), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT38), .B1(new_n466), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n461), .A2(new_n509), .A3(new_n277), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n468), .A2(new_n246), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n460), .A2(new_n246), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT87), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n510), .B(KEYINPUT37), .C1(new_n511), .C2(new_n513), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n508), .A2(new_n514), .B1(new_n451), .B2(new_n469), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n448), .B1(new_n461), .B2(new_n277), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n452), .B1(new_n516), .B2(KEYINPUT37), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT37), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n469), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT38), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n496), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n407), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(KEYINPUT39), .C1(new_n407), .C2(new_n405), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT39), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n525), .A3(new_n407), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n526), .A2(KEYINPUT86), .A3(new_n484), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT86), .B1(new_n526), .B2(new_n484), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT40), .B(new_n524), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n495), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n521), .B(new_n490), .C1(new_n533), .C2(new_n498), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n506), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n501), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G197gat), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT11), .B(G169gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT12), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR3_X1   g341(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(KEYINPUT89), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G29gat), .A2(G36gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n285), .A2(G43gat), .ZN(new_n550));
  INV_X1    g349(.A(G43gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G50gat), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n550), .A2(new_n552), .A3(KEYINPUT15), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(KEYINPUT90), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n545), .A2(new_n546), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n553), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n544), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(new_n543), .ZN(new_n560));
  AOI211_X1 g359(.A(new_n553), .B(new_n560), .C1(G29gat), .C2(G36gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT15), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n550), .B(KEYINPUT91), .Z(new_n563));
  XOR2_X1   g362(.A(KEYINPUT92), .B(G50gat), .Z(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(G43gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n562), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n554), .A2(new_n558), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT16), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(G1gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(G1gat), .B2(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n571), .B(G8gat), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n567), .B2(KEYINPUT17), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n566), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT90), .B1(new_n549), .B2(new_n553), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n556), .A2(new_n555), .A3(new_n557), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n574), .B1(new_n576), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(KEYINPUT13), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n567), .A2(new_n573), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n590), .B2(new_n574), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n585), .B1(new_n583), .B2(new_n586), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n542), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n582), .ZN(new_n595));
  INV_X1    g394(.A(new_n574), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n586), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n584), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(new_n587), .A3(new_n541), .A4(new_n591), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  XOR2_X1   g401(.A(G99gat), .B(G106gat), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n604), .B1(new_n606), .B2(new_n610), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n602), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n606), .A2(new_n610), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n603), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(KEYINPUT98), .A3(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G57gat), .B(G64gat), .Z(new_n620));
  INV_X1    g419(.A(KEYINPUT9), .ZN(new_n621));
  INV_X1    g420(.A(G71gat), .ZN(new_n622));
  INV_X1    g421(.A(G78gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G71gat), .B(G78gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n620), .A2(new_n626), .A3(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(KEYINPUT95), .A3(new_n629), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n634), .A3(KEYINPUT10), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n628), .B(new_n629), .C1(new_n612), .C2(new_n613), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n630), .A2(new_n611), .A3(new_n616), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI211_X1 g440(.A(KEYINPUT100), .B(KEYINPUT10), .C1(new_n637), .C2(new_n638), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n635), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n637), .A2(new_n638), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G120gat), .B(G148gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT101), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n645), .A2(new_n647), .A3(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT94), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  INV_X1    g459(.A(KEYINPUT21), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n632), .B2(new_n633), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT96), .B1(new_n662), .B2(new_n575), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n662), .A2(KEYINPUT96), .A3(new_n575), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n662), .A2(KEYINPUT96), .A3(new_n575), .ZN(new_n667));
  INV_X1    g466(.A(new_n660), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n630), .A2(new_n661), .ZN(new_n671));
  XOR2_X1   g470(.A(G127gat), .B(G155gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(G183gat), .B(G211gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n666), .A2(new_n675), .A3(new_n669), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n567), .A2(KEYINPUT17), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n582), .A2(new_n680), .A3(new_n618), .ZN(new_n681));
  AND2_X1   g480(.A1(G232gat), .A2(G233gat), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n619), .A2(new_n580), .B1(KEYINPUT41), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G190gat), .B(G218gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT99), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n682), .A2(KEYINPUT41), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  XNOR2_X1  g488(.A(G134gat), .B(G162gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n686), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n681), .A2(new_n692), .A3(new_n683), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n687), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n691), .ZN(new_n695));
  INV_X1    g494(.A(new_n693), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n681), .B2(new_n683), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n601), .A2(new_n656), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n536), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n435), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n498), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(KEYINPUT102), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n706), .A2(KEYINPUT102), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT42), .B1(new_n704), .B2(new_n572), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n704), .A2(new_n705), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n707), .B1(new_n708), .B2(new_n711), .ZN(G1325gat));
  INV_X1    g511(.A(new_n504), .ZN(new_n713));
  OAI21_X1  g512(.A(G15gat), .B1(new_n701), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n400), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n701), .B2(new_n715), .ZN(G1326gat));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n490), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT103), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT43), .B(G22gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  NAND2_X1  g519(.A1(new_n698), .A2(new_n694), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n501), .B2(new_n535), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n601), .A2(new_n656), .A3(new_n679), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n435), .ZN(new_n726));
  INV_X1    g525(.A(G29gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n725), .A2(KEYINPUT104), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT104), .B1(new_n725), .B2(new_n728), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n729), .A2(KEYINPUT45), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT45), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n698), .A2(KEYINPUT105), .A3(new_n694), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT105), .B1(new_n698), .B2(new_n694), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(KEYINPUT44), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n536), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT106), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n536), .A2(new_n721), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT44), .ZN(new_n741));
  INV_X1    g540(.A(new_n737), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n501), .B2(new_n535), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n739), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n746), .A2(new_n726), .A3(new_n724), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n733), .B1(new_n727), .B2(new_n747), .ZN(G1328gat));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n479), .A3(new_n724), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n746), .A2(KEYINPUT107), .A3(new_n479), .A4(new_n724), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(G36gat), .A3(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n725), .A2(G36gat), .A3(new_n498), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1329gat));
  NAND4_X1  g555(.A1(new_n746), .A2(G43gat), .A3(new_n504), .A4(new_n724), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n551), .B1(new_n725), .B2(new_n400), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n757), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1330gat));
  NOR2_X1   g562(.A1(new_n490), .A2(new_n564), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n724), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n564), .B1(new_n725), .B2(new_n490), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT48), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT48), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1331gat));
  NOR2_X1   g570(.A1(new_n699), .A2(new_n600), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n656), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n536), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n726), .A2(KEYINPUT109), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n435), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g581(.A1(new_n775), .A2(new_n498), .ZN(new_n783));
  NOR2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  AND2_X1   g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n783), .B2(new_n784), .ZN(G1333gat));
  NOR3_X1   g586(.A1(new_n775), .A2(new_n622), .A3(new_n713), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n400), .B(KEYINPUT110), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n536), .A2(new_n774), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(new_n622), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g591(.A1(new_n775), .A2(new_n490), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(new_n623), .ZN(G1335gat));
  INV_X1    g593(.A(new_n679), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n601), .A2(KEYINPUT111), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n600), .B2(new_n679), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n536), .A2(new_n721), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n796), .B2(new_n798), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n723), .A2(KEYINPUT112), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT112), .B1(new_n723), .B2(new_n803), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n806), .A2(new_n608), .A3(new_n726), .A4(new_n656), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n799), .A2(new_n656), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n740), .A2(KEYINPUT44), .B1(new_n743), .B2(new_n744), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n739), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n726), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n608), .ZN(G1336gat));
  AOI21_X1  g611(.A(new_n609), .B1(new_n810), .B2(new_n479), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n800), .A2(new_n801), .B1(new_n723), .B2(new_n803), .ZN(new_n815));
  INV_X1    g614(.A(new_n656), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n498), .A2(new_n816), .A3(G92gat), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n814), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT51), .B1(new_n723), .B2(new_n799), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n536), .A2(new_n721), .A3(new_n803), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT113), .B(new_n817), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT52), .B1(new_n813), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n808), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n738), .A2(KEYINPUT106), .B1(new_n723), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n743), .A2(new_n744), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n479), .B(new_n826), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G92gat), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n821), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n723), .A2(KEYINPUT112), .A3(new_n803), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n820), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT114), .B1(new_n835), .B2(new_n818), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n806), .A2(new_n837), .A3(new_n817), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n831), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n840), .ZN(G1337gat));
  AND2_X1   g640(.A1(new_n810), .A2(new_n504), .ZN(new_n842));
  INV_X1    g641(.A(G99gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n482), .A2(new_n656), .A3(new_n843), .ZN(new_n844));
  OAI22_X1  g643(.A1(new_n842), .A2(new_n843), .B1(new_n835), .B2(new_n844), .ZN(G1338gat));
  INV_X1    g644(.A(G106gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n810), .B2(new_n302), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n816), .A2(G106gat), .A3(new_n490), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT115), .B1(new_n815), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n851), .B(new_n848), .C1(new_n820), .C2(new_n822), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT53), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n302), .B(new_n826), .C1(new_n828), .C2(new_n829), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(G106gat), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT116), .B1(new_n835), .B2(new_n849), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n806), .A2(new_n858), .A3(new_n848), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n856), .A2(new_n857), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n854), .A2(new_n861), .ZN(G1339gat));
  NOR2_X1   g661(.A1(new_n734), .A2(new_n735), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n639), .A2(new_n640), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT100), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n639), .A2(new_n636), .A3(new_n640), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n646), .A3(new_n635), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n869), .A2(new_n645), .A3(KEYINPUT54), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n653), .B1(new_n645), .B2(KEYINPUT54), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n646), .B1(new_n868), .B2(new_n635), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n652), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n645), .A3(KEYINPUT54), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(KEYINPUT55), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n600), .A2(new_n872), .A3(new_n655), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n583), .A2(new_n586), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n590), .A2(new_n574), .A3(new_n588), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n540), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n599), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n656), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n863), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n882), .A2(new_n872), .A3(new_n655), .A4(new_n877), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n736), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n795), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n699), .A2(new_n600), .A3(new_n656), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n302), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n479), .A2(new_n435), .A3(new_n400), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n600), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G113gat), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n887), .A2(new_n889), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n780), .A2(new_n479), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n401), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n601), .A2(new_n356), .A3(new_n355), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(G1340gat));
  INV_X1    g699(.A(new_n898), .ZN(new_n901));
  AOI21_X1  g700(.A(G120gat), .B1(new_n901), .B2(new_n656), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n656), .A2(G120gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n892), .B2(new_n903), .ZN(G1341gat));
  NOR3_X1   g703(.A1(new_n898), .A2(G127gat), .A3(new_n795), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n906));
  INV_X1    g705(.A(G127gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n892), .B2(new_n679), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n905), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1342gat));
  NOR2_X1   g710(.A1(new_n722), .A2(G134gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n401), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n913), .B2(KEYINPUT56), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n913), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n892), .A2(new_n721), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G134gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n917), .A2(new_n922), .A3(new_n924), .ZN(G1343gat));
  NOR2_X1   g724(.A1(new_n504), .A2(new_n490), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n601), .A2(G141gat), .ZN(new_n927));
  AND4_X1   g726(.A1(new_n895), .A2(new_n896), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n504), .A2(new_n479), .A3(new_n435), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT57), .B1(new_n895), .B2(new_n302), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n302), .A2(KEYINPUT57), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n721), .B1(new_n878), .B2(new_n883), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n795), .B1(new_n886), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n933), .B2(new_n889), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n600), .B(new_n929), .C1(new_n930), .C2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n218), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n928), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n937), .B(new_n939), .ZN(G1344gat));
  AND2_X1   g739(.A1(new_n929), .A2(new_n656), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n877), .A2(new_n655), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT55), .B1(new_n875), .B2(new_n876), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n599), .A2(new_n881), .ZN(new_n944));
  NOR4_X1   g743(.A1(new_n942), .A2(new_n722), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n795), .B1(new_n932), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n947), .B1(new_n772), .B2(new_n816), .ZN(new_n948));
  NOR4_X1   g747(.A1(new_n699), .A2(new_n600), .A3(KEYINPUT121), .A4(new_n656), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT57), .B1(new_n951), .B2(new_n302), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n931), .B1(new_n887), .B2(new_n889), .ZN(new_n953));
  OAI211_X1 g752(.A(KEYINPUT122), .B(new_n941), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G148gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n878), .A2(new_n883), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n736), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n943), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n863), .A3(new_n882), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n679), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(new_n888), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n490), .B1(new_n946), .B2(new_n950), .ZN(new_n962));
  OAI22_X1  g761(.A1(new_n961), .A2(new_n931), .B1(new_n962), .B2(KEYINPUT57), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT122), .B1(new_n963), .B2(new_n941), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT59), .B1(new_n955), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n204), .A2(KEYINPUT59), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n929), .B1(new_n930), .B2(new_n934), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n816), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n897), .A2(new_n926), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n204), .A3(new_n656), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1345gat));
  OAI21_X1  g771(.A(G155gat), .B1(new_n967), .B2(new_n795), .ZN(new_n973));
  INV_X1    g772(.A(G155gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n974), .A3(new_n679), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1346gat));
  NAND2_X1  g775(.A1(new_n863), .A2(G162gat), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n967), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(G162gat), .B1(new_n970), .B2(new_n721), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(G1347gat));
  AOI211_X1 g780(.A(new_n726), .B(new_n498), .C1(new_n887), .C2(new_n889), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(new_n401), .ZN(new_n983));
  INV_X1    g782(.A(G169gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n983), .A2(new_n984), .A3(new_n600), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT123), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n780), .A2(new_n479), .A3(new_n789), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n890), .A2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(new_n600), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n986), .B1(new_n990), .B2(G169gat), .ZN(new_n991));
  AOI211_X1 g790(.A(KEYINPUT123), .B(new_n984), .C1(new_n989), .C2(new_n600), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n985), .B1(new_n991), .B2(new_n992), .ZN(G1348gat));
  INV_X1    g792(.A(G176gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n983), .A2(new_n994), .A3(new_n656), .ZN(new_n995));
  OAI21_X1  g794(.A(G176gat), .B1(new_n988), .B2(new_n816), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1349gat));
  OAI21_X1  g796(.A(KEYINPUT124), .B1(new_n988), .B2(new_n795), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n890), .A2(new_n999), .A3(new_n679), .A4(new_n987), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n998), .A2(G183gat), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n321), .A3(new_n679), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT60), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT60), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1350gat));
  NAND3_X1  g806(.A1(new_n983), .A2(new_n316), .A3(new_n863), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n989), .A2(new_n721), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1009), .B1(new_n1010), .B2(G190gat), .ZN(new_n1011));
  AOI211_X1 g810(.A(KEYINPUT61), .B(new_n316), .C1(new_n989), .C2(new_n721), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(G1351gat));
  AND2_X1   g812(.A1(new_n982), .A2(new_n926), .ZN(new_n1014));
  AOI21_X1  g813(.A(G197gat), .B1(new_n1014), .B2(new_n600), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n779), .A2(new_n498), .A3(new_n504), .ZN(new_n1016));
  XNOR2_X1  g815(.A(new_n1016), .B(KEYINPUT125), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n963), .A2(new_n1017), .ZN(new_n1018));
  AND2_X1   g817(.A1(new_n600), .A2(G197gat), .ZN(new_n1019));
  AOI21_X1  g818(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(G1352gat));
  INV_X1    g819(.A(G204gat), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n963), .A2(new_n1017), .A3(new_n656), .ZN(new_n1022));
  AOI21_X1  g821(.A(new_n1021), .B1(new_n1022), .B2(KEYINPUT126), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1023), .B1(KEYINPUT126), .B2(new_n1022), .ZN(new_n1024));
  NAND4_X1  g823(.A1(new_n982), .A2(new_n1021), .A3(new_n656), .A4(new_n926), .ZN(new_n1025));
  XOR2_X1   g824(.A(new_n1025), .B(KEYINPUT62), .Z(new_n1026));
  NAND2_X1  g825(.A1(new_n1024), .A2(new_n1026), .ZN(G1353gat));
  NAND3_X1  g826(.A1(new_n1014), .A2(new_n239), .A3(new_n679), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n963), .A2(new_n1016), .A3(new_n679), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n1029), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1030));
  AOI21_X1  g829(.A(KEYINPUT63), .B1(new_n1029), .B2(G211gat), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(G1354gat));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n963), .A2(new_n1017), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n1034), .A2(new_n721), .ZN(new_n1035));
  AOI21_X1  g834(.A(new_n1033), .B1(new_n963), .B2(new_n1017), .ZN(new_n1036));
  OAI21_X1  g835(.A(G218gat), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g836(.A1(new_n1014), .A2(new_n240), .A3(new_n863), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1037), .A2(new_n1038), .ZN(G1355gat));
endmodule


