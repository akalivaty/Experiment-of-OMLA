

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599;

  NOR2_X1 U325 ( .A1(n596), .A2(n465), .ZN(n466) );
  XOR2_X1 U326 ( .A(n489), .B(KEYINPUT28), .Z(n544) );
  XNOR2_X1 U327 ( .A(n426), .B(n425), .ZN(n533) );
  XOR2_X1 U328 ( .A(n316), .B(n446), .Z(n293) );
  NOR2_X1 U329 ( .A1(n438), .A2(n484), .ZN(n427) );
  XNOR2_X1 U330 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n473) );
  XNOR2_X1 U331 ( .A(n474), .B(n473), .ZN(n481) );
  XNOR2_X1 U332 ( .A(n362), .B(n361), .ZN(n371) );
  XNOR2_X1 U333 ( .A(n485), .B(KEYINPUT54), .ZN(n486) );
  XNOR2_X1 U334 ( .A(n384), .B(KEYINPUT22), .ZN(n385) );
  XNOR2_X1 U335 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U336 ( .A(n293), .B(n320), .ZN(n321) );
  XNOR2_X1 U337 ( .A(n386), .B(n385), .ZN(n391) );
  XNOR2_X1 U338 ( .A(n322), .B(n321), .ZN(n323) );
  INV_X1 U339 ( .A(KEYINPUT58), .ZN(n493) );
  XOR2_X1 U340 ( .A(KEYINPUT38), .B(n467), .Z(n516) );
  XNOR2_X1 U341 ( .A(n493), .B(G190GAT), .ZN(n494) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n468) );
  XNOR2_X1 U343 ( .A(n495), .B(n494), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n469), .B(n468), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(G176GAT), .B(G64GAT), .Z(n416) );
  XOR2_X1 U346 ( .A(G85GAT), .B(G92GAT), .Z(n331) );
  XNOR2_X1 U347 ( .A(n416), .B(n331), .ZN(n308) );
  XOR2_X1 U348 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n295) );
  NAND2_X1 U349 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n297) );
  INV_X1 U351 ( .A(KEYINPUT32), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U353 ( .A(G78GAT), .B(G106GAT), .Z(n299) );
  XNOR2_X1 U354 ( .A(G148GAT), .B(G204GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n381) );
  XNOR2_X1 U356 ( .A(G120GAT), .B(G99GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n300), .B(G71GAT), .ZN(n407) );
  XNOR2_X1 U358 ( .A(n381), .B(n407), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n304) );
  INV_X1 U360 ( .A(KEYINPUT31), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U362 ( .A(G57GAT), .B(KEYINPUT13), .Z(n445) );
  XNOR2_X1 U363 ( .A(n445), .B(KEYINPUT71), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n586) );
  XOR2_X1 U366 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n310) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(KEYINPUT70), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n324) );
  XOR2_X1 U369 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n312) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(KEYINPUT68), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n334) );
  XOR2_X1 U372 ( .A(n334), .B(G141GAT), .Z(n314) );
  NAND2_X1 U373 ( .A1(G229GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n322) );
  XNOR2_X1 U375 ( .A(G50GAT), .B(G43GAT), .ZN(n316) );
  XNOR2_X1 U376 ( .A(G1GAT), .B(G15GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n315), .B(KEYINPUT69), .ZN(n446) );
  XOR2_X1 U378 ( .A(G36GAT), .B(G8GAT), .Z(n417) );
  XOR2_X1 U379 ( .A(KEYINPUT29), .B(G22GAT), .Z(n318) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(G169GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n417), .B(n319), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n580) );
  NOR2_X1 U384 ( .A1(n586), .A2(n580), .ZN(n504) );
  XOR2_X1 U385 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n326) );
  XNOR2_X1 U386 ( .A(G190GAT), .B(G99GAT), .ZN(n325) );
  XNOR2_X1 U387 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U388 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n328) );
  XNOR2_X1 U389 ( .A(KEYINPUT74), .B(G106GAT), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n342) );
  XOR2_X1 U392 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n333) );
  XOR2_X1 U393 ( .A(G162GAT), .B(G50GAT), .Z(n372) );
  XNOR2_X1 U394 ( .A(n372), .B(n331), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U396 ( .A(G134GAT), .B(G43GAT), .Z(n400) );
  XNOR2_X1 U397 ( .A(n400), .B(n334), .ZN(n336) );
  AND2_X1 U398 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U400 ( .A(n338), .B(n337), .Z(n340) );
  XNOR2_X1 U401 ( .A(G218GAT), .B(G36GAT), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n555) );
  XOR2_X1 U404 ( .A(n555), .B(KEYINPUT36), .Z(n596) );
  NAND2_X1 U405 ( .A1(G225GAT), .A2(G233GAT), .ZN(n348) );
  XOR2_X1 U406 ( .A(G148GAT), .B(KEYINPUT74), .Z(n344) );
  XNOR2_X1 U407 ( .A(G162GAT), .B(G85GAT), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U409 ( .A(G134GAT), .B(G29GAT), .Z(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n370) );
  XOR2_X1 U412 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n350) );
  XNOR2_X1 U413 ( .A(KEYINPUT6), .B(KEYINPUT93), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n368) );
  XOR2_X1 U415 ( .A(G155GAT), .B(G57GAT), .Z(n352) );
  XNOR2_X1 U416 ( .A(G1GAT), .B(G120GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U418 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n354) );
  XNOR2_X1 U419 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U421 ( .A(n356), .B(n355), .Z(n366) );
  INV_X1 U422 ( .A(KEYINPUT90), .ZN(n357) );
  NAND2_X1 U423 ( .A1(n357), .A2(KEYINPUT2), .ZN(n360) );
  INV_X1 U424 ( .A(KEYINPUT2), .ZN(n358) );
  NAND2_X1 U425 ( .A1(n358), .A2(KEYINPUT90), .ZN(n359) );
  NAND2_X1 U426 ( .A1(n360), .A2(n359), .ZN(n362) );
  XNOR2_X1 U427 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n361) );
  XOR2_X1 U428 ( .A(KEYINPUT79), .B(KEYINPUT0), .Z(n364) );
  XNOR2_X1 U429 ( .A(G113GAT), .B(G127GAT), .ZN(n363) );
  XNOR2_X1 U430 ( .A(n364), .B(n363), .ZN(n408) );
  XNOR2_X1 U431 ( .A(n371), .B(n408), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U433 ( .A(n368), .B(n367), .Z(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n531) );
  XOR2_X1 U435 ( .A(KEYINPUT100), .B(KEYINPUT25), .Z(n431) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n376) );
  INV_X1 U437 ( .A(n376), .ZN(n374) );
  AND2_X1 U438 ( .A1(G228GAT), .A2(G233GAT), .ZN(n375) );
  INV_X1 U439 ( .A(n375), .ZN(n373) );
  NAND2_X1 U440 ( .A1(n374), .A2(n373), .ZN(n378) );
  NAND2_X1 U441 ( .A1(n376), .A2(n375), .ZN(n377) );
  NAND2_X1 U442 ( .A1(n378), .A2(n377), .ZN(n380) );
  INV_X1 U443 ( .A(KEYINPUT23), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n381), .B(KEYINPUT91), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n386) );
  XOR2_X1 U447 ( .A(G155GAT), .B(G22GAT), .Z(n457) );
  XNOR2_X1 U448 ( .A(n457), .B(KEYINPUT24), .ZN(n384) );
  XNOR2_X1 U449 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n387), .B(KEYINPUT88), .ZN(n388) );
  XOR2_X1 U451 ( .A(n388), .B(G197GAT), .Z(n390) );
  XNOR2_X1 U452 ( .A(KEYINPUT89), .B(G218GAT), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n425) );
  XNOR2_X1 U454 ( .A(n391), .B(n425), .ZN(n489) );
  INV_X1 U455 ( .A(n489), .ZN(n429) );
  XOR2_X1 U456 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n393) );
  XNOR2_X1 U457 ( .A(G183GAT), .B(KEYINPUT85), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U459 ( .A(n394), .B(G169GAT), .Z(n396) );
  XNOR2_X1 U460 ( .A(KEYINPUT19), .B(G190GAT), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n424) );
  XOR2_X1 U462 ( .A(KEYINPUT83), .B(KEYINPUT86), .Z(n398) );
  XNOR2_X1 U463 ( .A(KEYINPUT20), .B(KEYINPUT81), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U465 ( .A(n399), .B(G15GAT), .Z(n402) );
  XNOR2_X1 U466 ( .A(G176GAT), .B(n400), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n424), .B(n403), .ZN(n412) );
  XOR2_X1 U469 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n405) );
  NAND2_X1 U470 ( .A1(G227GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U472 ( .A(n406), .B(KEYINPUT84), .Z(n410) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n438) );
  XOR2_X1 U476 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n414) );
  XNOR2_X1 U477 ( .A(KEYINPUT75), .B(KEYINPUT98), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n420) );
  XOR2_X1 U479 ( .A(G204GAT), .B(G92GAT), .Z(n415) );
  XNOR2_X1 U480 ( .A(n416), .B(n415), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U482 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U483 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n426) );
  INV_X1 U486 ( .A(n533), .ZN(n484) );
  XOR2_X1 U487 ( .A(KEYINPUT99), .B(n427), .Z(n428) );
  NOR2_X1 U488 ( .A1(n429), .A2(n428), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n434) );
  XNOR2_X1 U490 ( .A(KEYINPUT27), .B(n533), .ZN(n437) );
  INV_X1 U491 ( .A(n438), .ZN(n542) );
  OR2_X1 U492 ( .A1(n489), .A2(n542), .ZN(n432) );
  XOR2_X1 U493 ( .A(n432), .B(KEYINPUT26), .Z(n578) );
  AND2_X1 U494 ( .A1(n437), .A2(n578), .ZN(n433) );
  NOR2_X1 U495 ( .A1(n434), .A2(n433), .ZN(n435) );
  NOR2_X1 U496 ( .A1(n531), .A2(n435), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n436), .B(KEYINPUT101), .ZN(n443) );
  NAND2_X1 U498 ( .A1(n531), .A2(n437), .ZN(n541) );
  XNOR2_X1 U499 ( .A(KEYINPUT87), .B(n438), .ZN(n439) );
  NOR2_X1 U500 ( .A1(n541), .A2(n439), .ZN(n441) );
  INV_X1 U501 ( .A(n544), .ZN(n440) );
  NAND2_X1 U502 ( .A1(n441), .A2(n440), .ZN(n442) );
  NAND2_X1 U503 ( .A1(n443), .A2(n442), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n444), .B(KEYINPUT102), .ZN(n501) );
  XOR2_X1 U505 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U506 ( .A1(G231GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n464) );
  XOR2_X1 U508 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n450) );
  XNOR2_X1 U509 ( .A(KEYINPUT76), .B(KEYINPUT14), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n454) );
  XOR2_X1 U511 ( .A(KEYINPUT75), .B(G183GAT), .Z(n452) );
  XNOR2_X1 U512 ( .A(G127GAT), .B(G211GAT), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n462) );
  XOR2_X1 U515 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n456) );
  XNOR2_X1 U516 ( .A(G78GAT), .B(G71GAT), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n456), .B(n455), .ZN(n458) );
  XOR2_X1 U518 ( .A(n458), .B(n457), .Z(n460) );
  XNOR2_X1 U519 ( .A(G64GAT), .B(G8GAT), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(n592) );
  NAND2_X1 U523 ( .A1(n501), .A2(n592), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT37), .B(n466), .Z(n530) );
  NAND2_X1 U525 ( .A1(n504), .A2(n530), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n516), .A2(n542), .ZN(n469) );
  INV_X1 U527 ( .A(n555), .ZN(n567) );
  NAND2_X1 U528 ( .A1(n567), .A2(n592), .ZN(n472) );
  INV_X1 U529 ( .A(n580), .ZN(n545) );
  XOR2_X1 U530 ( .A(n586), .B(KEYINPUT41), .Z(n518) );
  AND2_X1 U531 ( .A1(n545), .A2(n518), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT46), .ZN(n471) );
  OR2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n474) );
  OR2_X1 U534 ( .A1(n596), .A2(n592), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U537 ( .A1(n586), .A2(n477), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT112), .B(n478), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n479), .A2(n580), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n481), .A2(n480), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT113), .B(KEYINPUT48), .Z(n482) );
  XOR2_X1 U542 ( .A(n483), .B(n482), .Z(n540) );
  NOR2_X1 U543 ( .A1(n540), .A2(n484), .ZN(n487) );
  INV_X1 U544 ( .A(KEYINPUT118), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n531), .A2(n488), .ZN(n579) );
  NAND2_X1 U546 ( .A1(n579), .A2(n489), .ZN(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n492) );
  NAND2_X1 U549 ( .A1(n492), .A2(n542), .ZN(n575) );
  NOR2_X1 U550 ( .A1(n567), .A2(n575), .ZN(n495) );
  NAND2_X1 U551 ( .A1(n531), .A2(n516), .ZN(n499) );
  XOR2_X1 U552 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n497) );
  INV_X1 U553 ( .A(G29GAT), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U555 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n555), .A2(n592), .ZN(n500) );
  XNOR2_X1 U557 ( .A(KEYINPUT16), .B(n500), .ZN(n502) );
  NAND2_X1 U558 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U559 ( .A(n503), .B(KEYINPUT103), .ZN(n519) );
  NAND2_X1 U560 ( .A1(n504), .A2(n519), .ZN(n505) );
  XOR2_X1 U561 ( .A(KEYINPUT104), .B(n505), .Z(n512) );
  NAND2_X1 U562 ( .A1(n512), .A2(n531), .ZN(n506) );
  XNOR2_X1 U563 ( .A(n506), .B(KEYINPUT34), .ZN(n507) );
  XNOR2_X1 U564 ( .A(G1GAT), .B(n507), .ZN(G1324GAT) );
  NAND2_X1 U565 ( .A1(n533), .A2(n512), .ZN(n508) );
  XNOR2_X1 U566 ( .A(G8GAT), .B(n508), .ZN(G1325GAT) );
  NAND2_X1 U567 ( .A1(n512), .A2(n542), .ZN(n511) );
  XNOR2_X1 U568 ( .A(G15GAT), .B(KEYINPUT105), .ZN(n509) );
  XNOR2_X1 U569 ( .A(n509), .B(KEYINPUT35), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n511), .B(n510), .ZN(G1326GAT) );
  XNOR2_X1 U571 ( .A(G22GAT), .B(KEYINPUT106), .ZN(n514) );
  NAND2_X1 U572 ( .A1(n544), .A2(n512), .ZN(n513) );
  XNOR2_X1 U573 ( .A(n514), .B(n513), .ZN(G1327GAT) );
  NAND2_X1 U574 ( .A1(n516), .A2(n533), .ZN(n515) );
  XNOR2_X1 U575 ( .A(n515), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U576 ( .A1(n516), .A2(n544), .ZN(n517) );
  XNOR2_X1 U577 ( .A(n517), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n521) );
  INV_X1 U579 ( .A(n518), .ZN(n571) );
  NOR2_X1 U580 ( .A1(n545), .A2(n571), .ZN(n529) );
  AND2_X1 U581 ( .A1(n519), .A2(n529), .ZN(n525) );
  NAND2_X1 U582 ( .A1(n525), .A2(n531), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  NAND2_X1 U585 ( .A1(n525), .A2(n533), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n542), .A2(n525), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n527) );
  NAND2_X1 U590 ( .A1(n525), .A2(n544), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(G78GAT), .B(n528), .Z(G1335GAT) );
  AND2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n531), .A2(n537), .ZN(n532) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n532), .ZN(G1336GAT) );
  NAND2_X1 U596 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(KEYINPUT110), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n535), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n542), .A2(n537), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U601 ( .A1(n537), .A2(n544), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n559) );
  NAND2_X1 U606 ( .A1(n559), .A2(n542), .ZN(n543) );
  NOR2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n556) );
  NAND2_X1 U608 ( .A1(n545), .A2(n556), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U611 ( .A1(n556), .A2(n518), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  INV_X1 U613 ( .A(n592), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n556), .A2(n550), .ZN(n554) );
  XOR2_X1 U615 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n552) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  NAND2_X1 U622 ( .A1(n559), .A2(n578), .ZN(n566) );
  NOR2_X1 U623 ( .A1(n580), .A2(n566), .ZN(n560) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n560), .Z(G1344GAT) );
  NOR2_X1 U625 ( .A1(n571), .A2(n566), .ZN(n562) );
  XNOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NOR2_X1 U629 ( .A1(n592), .A2(n566), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1346GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(G162GAT), .B(n568), .Z(G1347GAT) );
  NOR2_X1 U634 ( .A1(n575), .A2(n580), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT120), .B(n569), .Z(n570) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(n570), .ZN(G1348GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n575), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(n574), .ZN(G1349GAT) );
  NOR2_X1 U641 ( .A1(n592), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1350GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n595) );
  NOR2_X1 U645 ( .A1(n580), .A2(n595), .ZN(n585) );
  XOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n582) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(KEYINPUT59), .B(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  INV_X1 U651 ( .A(n586), .ZN(n587) );
  NOR2_X1 U652 ( .A1(n595), .A2(n587), .ZN(n591) );
  XOR2_X1 U653 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n589) );
  XNOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  NOR2_X1 U657 ( .A1(n592), .A2(n595), .ZN(n593) );
  XOR2_X1 U658 ( .A(KEYINPUT126), .B(n593), .Z(n594) );
  XNOR2_X1 U659 ( .A(G211GAT), .B(n594), .ZN(G1354GAT) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U661 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(n599), .ZN(G1355GAT) );
endmodule

