

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794;

  OR2_X1 U371 ( .A1(n388), .A2(n404), .ZN(n391) );
  NOR2_X1 U372 ( .A1(n353), .A2(n591), .ZN(n593) );
  BUF_X1 U373 ( .A(G143), .Z(n611) );
  XNOR2_X2 U374 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X2 U375 ( .A1(n360), .A2(n358), .ZN(n357) );
  INV_X2 U376 ( .A(G143), .ZN(n486) );
  XOR2_X1 U377 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n556) );
  INV_X1 U378 ( .A(G146), .ZN(n488) );
  XOR2_X1 U379 ( .A(KEYINPUT70), .B(KEYINPUT78), .Z(n350) );
  XOR2_X1 U380 ( .A(KEYINPUT89), .B(KEYINPUT63), .Z(n351) );
  XNOR2_X1 U381 ( .A(n686), .B(KEYINPUT66), .ZN(n352) );
  AND2_X1 U382 ( .A1(n766), .A2(n449), .ZN(n442) );
  INV_X1 U383 ( .A(n672), .ZN(n353) );
  NAND2_X1 U384 ( .A1(n367), .A2(n354), .ZN(n366) );
  NAND2_X1 U385 ( .A1(n359), .A2(n354), .ZN(n358) );
  XNOR2_X1 U386 ( .A(n363), .B(n352), .ZN(G60) );
  XNOR2_X1 U387 ( .A(n371), .B(n351), .ZN(G57) );
  AND2_X1 U388 ( .A1(n413), .A2(n412), .ZN(n743) );
  AND2_X1 U389 ( .A1(n432), .A2(n369), .ZN(n368) );
  AND2_X1 U390 ( .A1(n758), .A2(n361), .ZN(n360) );
  NOR2_X1 U391 ( .A1(n462), .A2(n461), .ZN(n416) );
  NAND2_X1 U392 ( .A1(n403), .A2(n401), .ZN(n705) );
  XNOR2_X1 U393 ( .A(n450), .B(n656), .ZN(n674) );
  NOR2_X1 U394 ( .A1(n724), .A2(n729), .ZN(n649) );
  XNOR2_X1 U395 ( .A(n478), .B(n392), .ZN(n723) );
  XNOR2_X1 U396 ( .A(n646), .B(n645), .ZN(n727) );
  NAND2_X1 U397 ( .A1(n418), .A2(n422), .ZN(n417) );
  INV_X1 U398 ( .A(n430), .ZN(n646) );
  XNOR2_X1 U399 ( .A(n428), .B(n499), .ZN(n425) );
  NAND2_X1 U400 ( .A1(n689), .A2(n370), .ZN(n367) );
  NOR2_X1 U401 ( .A1(n689), .A2(n370), .ZN(n369) );
  NAND2_X1 U402 ( .A1(n684), .A2(n362), .ZN(n359) );
  NOR2_X1 U403 ( .A1(n684), .A2(n362), .ZN(n361) );
  XNOR2_X1 U404 ( .A(n542), .B(n541), .ZN(n688) );
  XNOR2_X1 U405 ( .A(n498), .B(n497), .ZN(n499) );
  INV_X1 U406 ( .A(n765), .ZN(n354) );
  XNOR2_X2 U407 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n485) );
  XNOR2_X2 U408 ( .A(KEYINPUT16), .B(G122), .ZN(n483) );
  INV_X1 U409 ( .A(G237), .ZN(n495) );
  XOR2_X1 U410 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n554) );
  XOR2_X2 U411 ( .A(KEYINPUT9), .B(G122), .Z(n565) );
  XNOR2_X1 U412 ( .A(G116), .B(G107), .ZN(n564) );
  INV_X2 U413 ( .A(KEYINPUT76), .ZN(n411) );
  NAND2_X1 U414 ( .A1(n793), .A2(n794), .ZN(n660) );
  XNOR2_X2 U415 ( .A(n654), .B(KEYINPUT42), .ZN(n793) );
  NAND2_X1 U416 ( .A1(n402), .A2(n390), .ZN(n401) );
  NAND2_X1 U417 ( .A1(n727), .A2(n726), .ZN(n724) );
  NAND2_X1 U418 ( .A1(n408), .A2(n405), .ZN(n678) );
  XNOR2_X1 U419 ( .A(n456), .B(n455), .ZN(n454) );
  AND2_X2 U420 ( .A1(n766), .A2(n394), .ZN(n438) );
  NAND2_X1 U421 ( .A1(n357), .A2(n355), .ZN(n363) );
  NAND2_X1 U422 ( .A1(n356), .A2(n684), .ZN(n355) );
  INV_X1 U423 ( .A(n758), .ZN(n356) );
  INV_X1 U424 ( .A(G475), .ZN(n362) );
  NAND2_X1 U425 ( .A1(n365), .A2(n364), .ZN(n371) );
  NAND2_X1 U426 ( .A1(n356), .A2(n689), .ZN(n364) );
  NOR2_X1 U427 ( .A1(n368), .A2(n366), .ZN(n365) );
  INV_X1 U428 ( .A(G472), .ZN(n370) );
  BUF_X1 U429 ( .A(n540), .Z(n372) );
  NAND2_X1 U430 ( .A1(n408), .A2(n376), .ZN(n373) );
  NAND2_X1 U431 ( .A1(n373), .A2(n374), .ZN(n403) );
  OR2_X1 U432 ( .A1(n375), .A2(KEYINPUT84), .ZN(n374) );
  INV_X1 U433 ( .A(n391), .ZN(n375) );
  AND2_X1 U434 ( .A1(n405), .A2(n391), .ZN(n376) );
  INV_X1 U435 ( .A(n651), .ZN(n377) );
  BUF_X1 U436 ( .A(n625), .Z(n378) );
  XNOR2_X1 U437 ( .A(n443), .B(n602), .ZN(n625) );
  NAND2_X1 U438 ( .A1(n448), .A2(n389), .ZN(n673) );
  BUF_X1 U439 ( .A(n634), .Z(n379) );
  XNOR2_X1 U440 ( .A(n660), .B(n434), .ZN(n448) );
  NOR2_X1 U441 ( .A1(n426), .A2(n680), .ZN(n380) );
  NOR2_X1 U442 ( .A1(n426), .A2(n680), .ZN(n432) );
  NAND2_X1 U443 ( .A1(n440), .A2(n439), .ZN(n426) );
  NOR2_X2 U444 ( .A1(n744), .A2(n676), .ZN(n428) );
  XNOR2_X1 U445 ( .A(n622), .B(KEYINPUT35), .ZN(n381) );
  BUF_X1 U446 ( .A(n752), .Z(n382) );
  XNOR2_X1 U447 ( .A(n622), .B(KEYINPUT35), .ZN(n790) );
  NOR2_X2 U448 ( .A1(n752), .A2(G902), .ZN(n427) );
  INV_X1 U449 ( .A(n691), .ZN(n452) );
  AND2_X1 U450 ( .A1(n726), .A2(KEYINPUT19), .ZN(n424) );
  XNOR2_X1 U451 ( .A(KEYINPUT4), .B(G131), .ZN(n511) );
  XNOR2_X1 U452 ( .A(G113), .B(KEYINPUT69), .ZN(n481) );
  INV_X1 U453 ( .A(KEYINPUT64), .ZN(n477) );
  NAND2_X1 U454 ( .A1(n676), .A2(n475), .ZN(n474) );
  NAND2_X1 U455 ( .A1(KEYINPUT2), .A2(n477), .ZN(n475) );
  XNOR2_X1 U456 ( .A(G478), .B(n574), .ZN(n607) );
  XNOR2_X1 U457 ( .A(n567), .B(n566), .ZN(n570) );
  XOR2_X1 U458 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n566) );
  XNOR2_X1 U459 ( .A(n649), .B(n648), .ZN(n709) );
  INV_X1 U460 ( .A(KEYINPUT41), .ZN(n648) );
  AND2_X1 U461 ( .A1(n437), .A2(n436), .ZN(n662) );
  NOR2_X1 U462 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U463 ( .A(n535), .B(KEYINPUT25), .ZN(n445) );
  INV_X1 U464 ( .A(KEYINPUT105), .ZN(n455) );
  NOR2_X1 U465 ( .A1(n699), .A2(n725), .ZN(n663) );
  INV_X1 U466 ( .A(KEYINPUT46), .ZN(n434) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n502) );
  XNOR2_X1 U468 ( .A(n488), .B(G125), .ZN(n524) );
  AND2_X1 U469 ( .A1(n508), .A2(n421), .ZN(n420) );
  NAND2_X1 U470 ( .A1(n501), .A2(n422), .ZN(n421) );
  INV_X1 U471 ( .A(KEYINPUT19), .ZN(n422) );
  XNOR2_X1 U472 ( .A(n458), .B(G140), .ZN(n525) );
  INV_X1 U473 ( .A(G137), .ZN(n458) );
  XOR2_X1 U474 ( .A(G122), .B(G113), .Z(n549) );
  XNOR2_X1 U475 ( .A(G104), .B(G140), .ZN(n555) );
  XNOR2_X1 U476 ( .A(n524), .B(n444), .ZN(n551) );
  INV_X1 U477 ( .A(KEYINPUT10), .ZN(n444) );
  XNOR2_X1 U478 ( .A(n525), .B(n457), .ZN(n513) );
  INV_X1 U479 ( .A(KEYINPUT79), .ZN(n457) );
  NAND2_X1 U480 ( .A1(n400), .A2(n605), .ZN(n399) );
  XOR2_X1 U481 ( .A(KEYINPUT5), .B(G137), .Z(n538) );
  XOR2_X1 U482 ( .A(n525), .B(n551), .Z(n781) );
  NAND2_X1 U483 ( .A1(n476), .A2(n474), .ZN(n473) );
  NAND2_X1 U484 ( .A1(n517), .A2(n477), .ZN(n476) );
  AND2_X1 U485 ( .A1(n708), .A2(KEYINPUT83), .ZN(n461) );
  AND2_X1 U486 ( .A1(n398), .A2(n396), .ZN(n655) );
  XNOR2_X1 U487 ( .A(n604), .B(n397), .ZN(n396) );
  NOR2_X1 U488 ( .A1(n653), .A2(n399), .ZN(n398) );
  INV_X1 U489 ( .A(KEYINPUT30), .ZN(n397) );
  XNOR2_X1 U490 ( .A(n547), .B(KEYINPUT99), .ZN(n691) );
  INV_X2 U491 ( .A(G953), .ZN(n783) );
  XNOR2_X1 U492 ( .A(n570), .B(n569), .ZN(n572) );
  AND2_X1 U493 ( .A1(n685), .A2(G953), .ZN(n765) );
  XNOR2_X1 U494 ( .A(n659), .B(n658), .ZN(n794) );
  NAND2_X1 U495 ( .A1(n468), .A2(n385), .ZN(n467) );
  INV_X1 U496 ( .A(KEYINPUT31), .ZN(n435) );
  BUF_X1 U497 ( .A(n691), .Z(n447) );
  INV_X1 U498 ( .A(G953), .ZN(n412) );
  XNOR2_X1 U499 ( .A(n414), .B(KEYINPUT121), .ZN(n413) );
  OR2_X1 U500 ( .A1(n763), .A2(G902), .ZN(n383) );
  XNOR2_X1 U501 ( .A(G101), .B(KEYINPUT90), .ZN(n384) );
  INV_X1 U502 ( .A(n712), .ZN(n400) );
  AND2_X1 U503 ( .A1(n353), .A2(n712), .ZN(n385) );
  XNOR2_X1 U504 ( .A(KEYINPUT120), .B(n742), .ZN(n386) );
  OR2_X1 U505 ( .A1(n643), .A2(n642), .ZN(n387) );
  AND2_X1 U506 ( .A1(n704), .A2(n675), .ZN(n388) );
  AND2_X1 U507 ( .A1(n665), .A2(n664), .ZN(n389) );
  AND2_X1 U508 ( .A1(n388), .A2(n404), .ZN(n390) );
  XOR2_X1 U509 ( .A(n616), .B(n615), .Z(n392) );
  NAND2_X1 U510 ( .A1(n466), .A2(KEYINPUT64), .ZN(n393) );
  AND2_X1 U511 ( .A1(n676), .A2(n477), .ZN(n394) );
  AND2_X1 U512 ( .A1(KEYINPUT83), .A2(n466), .ZN(n395) );
  INV_X1 U513 ( .A(n678), .ZN(n402) );
  INV_X1 U514 ( .A(KEYINPUT84), .ZN(n404) );
  NAND2_X1 U515 ( .A1(n407), .A2(n406), .ZN(n405) );
  INV_X1 U516 ( .A(n673), .ZN(n406) );
  NOR2_X1 U517 ( .A1(n702), .A2(KEYINPUT48), .ZN(n407) );
  AND2_X2 U518 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X1 U519 ( .A1(n702), .A2(KEYINPUT48), .ZN(n409) );
  NAND2_X1 U520 ( .A1(n673), .A2(KEYINPUT48), .ZN(n410) );
  XNOR2_X2 U521 ( .A(n411), .B(G104), .ZN(n471) );
  NAND2_X1 U522 ( .A1(n416), .A2(n415), .ZN(n414) );
  NAND2_X1 U523 ( .A1(n463), .A2(n465), .ZN(n415) );
  NAND2_X1 U524 ( .A1(n430), .A2(n726), .ZN(n667) );
  NAND2_X2 U525 ( .A1(n419), .A2(n417), .ZN(n509) );
  INV_X1 U526 ( .A(n425), .ZN(n418) );
  AND2_X2 U527 ( .A1(n423), .A2(n420), .ZN(n419) );
  NAND2_X1 U528 ( .A1(n425), .A2(n424), .ZN(n423) );
  NAND2_X1 U529 ( .A1(n440), .A2(n439), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X2 U531 ( .A(n657), .B(n577), .ZN(n698) );
  XNOR2_X2 U532 ( .A(n576), .B(n575), .ZN(n657) );
  XNOR2_X2 U533 ( .A(n427), .B(n516), .ZN(n606) );
  INV_X1 U534 ( .A(n653), .ZN(n436) );
  XNOR2_X1 U535 ( .A(n542), .B(n515), .ZN(n752) );
  XNOR2_X1 U536 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U537 ( .A(n667), .B(KEYINPUT19), .ZN(n429) );
  XNOR2_X1 U538 ( .A(n428), .B(n499), .ZN(n430) );
  NOR2_X2 U539 ( .A1(n472), .A2(n680), .ZN(n431) );
  NOR2_X1 U540 ( .A1(n426), .A2(n680), .ZN(n758) );
  NAND2_X1 U541 ( .A1(n433), .A2(n387), .ZN(n644) );
  XNOR2_X1 U542 ( .A(n639), .B(n638), .ZN(n433) );
  OR2_X2 U543 ( .A1(n442), .A2(n393), .ZN(n439) );
  OR2_X1 U544 ( .A1(n451), .A2(n698), .ZN(n582) );
  OR2_X1 U545 ( .A1(n451), .A2(n695), .ZN(n584) );
  XNOR2_X2 U546 ( .A(n580), .B(n435), .ZN(n451) );
  XNOR2_X2 U547 ( .A(n780), .B(G146), .ZN(n542) );
  XNOR2_X2 U548 ( .A(n571), .B(n511), .ZN(n780) );
  XNOR2_X2 U549 ( .A(n510), .B(G134), .ZN(n571) );
  XNOR2_X2 U550 ( .A(n486), .B(G128), .ZN(n510) );
  NAND2_X1 U551 ( .A1(n662), .A2(n429), .ZN(n699) );
  XNOR2_X1 U552 ( .A(n652), .B(KEYINPUT28), .ZN(n437) );
  NAND2_X1 U553 ( .A1(n438), .A2(n449), .ZN(n441) );
  AND2_X2 U554 ( .A1(n441), .A2(n473), .ZN(n440) );
  NAND2_X1 U555 ( .A1(n601), .A2(n600), .ZN(n443) );
  XNOR2_X2 U556 ( .A(n383), .B(n445), .ZN(n712) );
  XNOR2_X1 U557 ( .A(n446), .B(n529), .ZN(n532) );
  XNOR2_X1 U558 ( .A(n528), .B(n350), .ZN(n446) );
  NAND2_X1 U559 ( .A1(n453), .A2(n623), .ZN(n456) );
  XNOR2_X1 U560 ( .A(n705), .B(KEYINPUT77), .ZN(n449) );
  NAND2_X1 U561 ( .A1(n655), .A2(n727), .ZN(n450) );
  NAND2_X1 U562 ( .A1(n452), .A2(n451), .ZN(n453) );
  NAND2_X1 U563 ( .A1(n624), .A2(n454), .ZN(n626) );
  XNOR2_X2 U564 ( .A(n606), .B(KEYINPUT1), .ZN(n635) );
  XNOR2_X2 U565 ( .A(n459), .B(G119), .ZN(n482) );
  XNOR2_X2 U566 ( .A(G116), .B(KEYINPUT3), .ZN(n459) );
  NAND2_X1 U567 ( .A1(n460), .A2(n386), .ZN(n462) );
  NAND2_X1 U568 ( .A1(n464), .A2(n395), .ZN(n460) );
  INV_X1 U569 ( .A(n707), .ZN(n464) );
  NAND2_X1 U570 ( .A1(n464), .A2(n466), .ZN(n465) );
  NOR2_X1 U571 ( .A1(n708), .A2(KEYINPUT83), .ZN(n463) );
  INV_X1 U572 ( .A(KEYINPUT2), .ZN(n466) );
  NAND2_X1 U573 ( .A1(n791), .A2(n792), .ZN(n641) );
  XNOR2_X2 U574 ( .A(n467), .B(KEYINPUT32), .ZN(n792) );
  INV_X1 U575 ( .A(n379), .ZN(n468) );
  XNOR2_X2 U576 ( .A(n772), .B(KEYINPUT71), .ZN(n514) );
  XNOR2_X2 U577 ( .A(n384), .B(n469), .ZN(n772) );
  XNOR2_X2 U578 ( .A(n471), .B(n470), .ZN(n469) );
  XNOR2_X2 U579 ( .A(G110), .B(G107), .ZN(n470) );
  NAND2_X1 U580 ( .A1(n723), .A2(n617), .ZN(n619) );
  NAND2_X1 U581 ( .A1(n479), .A2(n635), .ZN(n478) );
  NOR2_X1 U582 ( .A1(n614), .A2(n613), .ZN(n479) );
  NOR2_X2 U583 ( .A1(n672), .A2(n671), .ZN(n702) );
  BUF_X1 U584 ( .A(n705), .Z(n782) );
  XNOR2_X1 U585 ( .A(n514), .B(n480), .ZN(n515) );
  NOR2_X2 U586 ( .A1(n579), .A2(n651), .ZN(n720) );
  BUF_X1 U587 ( .A(n744), .Z(n747) );
  XOR2_X1 U588 ( .A(n513), .B(n512), .Z(n480) );
  BUF_X1 U589 ( .A(n709), .Z(n739) );
  INV_X1 U590 ( .A(KEYINPUT86), .ZN(n638) );
  XNOR2_X1 U591 ( .A(KEYINPUT115), .B(KEYINPUT36), .ZN(n669) );
  XNOR2_X1 U592 ( .A(n670), .B(n669), .ZN(n671) );
  INV_X1 U593 ( .A(KEYINPUT106), .ZN(n602) );
  XNOR2_X2 U594 ( .A(n482), .B(n481), .ZN(n540) );
  XNOR2_X2 U595 ( .A(n540), .B(n483), .ZN(n774) );
  XNOR2_X2 U596 ( .A(KEYINPUT18), .B(KEYINPUT91), .ZN(n484) );
  XNOR2_X1 U597 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U598 ( .A(n510), .B(n487), .ZN(n492) );
  NAND2_X1 U599 ( .A1(n783), .A2(G224), .ZN(n489) );
  XNOR2_X1 U600 ( .A(n489), .B(KEYINPUT80), .ZN(n490) );
  XNOR2_X1 U601 ( .A(n524), .B(n490), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n774), .B(n493), .ZN(n494) );
  XNOR2_X1 U604 ( .A(n494), .B(n514), .ZN(n744) );
  XNOR2_X1 U605 ( .A(G902), .B(KEYINPUT15), .ZN(n517) );
  INV_X1 U606 ( .A(n517), .ZN(n676) );
  INV_X1 U607 ( .A(G902), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n543), .A2(n495), .ZN(n500) );
  NAND2_X1 U609 ( .A1(n500), .A2(G210), .ZN(n496) );
  XNOR2_X1 U610 ( .A(n496), .B(KEYINPUT93), .ZN(n498) );
  XNOR2_X1 U611 ( .A(KEYINPUT81), .B(KEYINPUT92), .ZN(n497) );
  NAND2_X1 U612 ( .A1(n500), .A2(G214), .ZN(n726) );
  INV_X1 U613 ( .A(n726), .ZN(n501) );
  XOR2_X1 U614 ( .A(KEYINPUT14), .B(KEYINPUT94), .Z(n503) );
  XOR2_X1 U615 ( .A(n503), .B(n502), .Z(n504) );
  NAND2_X1 U616 ( .A1(G952), .A2(n504), .ZN(n737) );
  NOR2_X1 U617 ( .A1(n737), .A2(G953), .ZN(n587) );
  INV_X1 U618 ( .A(n587), .ZN(n507) );
  AND2_X1 U619 ( .A1(n504), .A2(G953), .ZN(n505) );
  NAND2_X1 U620 ( .A1(G902), .A2(n505), .ZN(n585) );
  OR2_X1 U621 ( .A1(n585), .A2(G898), .ZN(n506) );
  NAND2_X1 U622 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X2 U623 ( .A(n509), .B(KEYINPUT0), .ZN(n598) );
  INV_X1 U624 ( .A(n598), .ZN(n617) );
  NAND2_X1 U625 ( .A1(G227), .A2(n783), .ZN(n512) );
  XOR2_X1 U626 ( .A(KEYINPUT68), .B(G469), .Z(n516) );
  NAND2_X1 U627 ( .A1(n517), .A2(G234), .ZN(n519) );
  XNOR2_X1 U628 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n518) );
  XNOR2_X1 U629 ( .A(n519), .B(n518), .ZN(n534) );
  AND2_X1 U630 ( .A1(n534), .A2(G221), .ZN(n523) );
  XOR2_X1 U631 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n521) );
  INV_X1 U632 ( .A(KEYINPUT21), .ZN(n520) );
  XNOR2_X1 U633 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U634 ( .A(n523), .B(n522), .ZN(n713) );
  XOR2_X1 U635 ( .A(KEYINPUT95), .B(G110), .Z(n527) );
  XNOR2_X1 U636 ( .A(G128), .B(G119), .ZN(n526) );
  XNOR2_X1 U637 ( .A(n527), .B(n526), .ZN(n529) );
  XOR2_X1 U638 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n528) );
  NAND2_X1 U639 ( .A1(G234), .A2(n783), .ZN(n530) );
  XOR2_X1 U640 ( .A(KEYINPUT8), .B(n530), .Z(n568) );
  NAND2_X1 U641 ( .A1(G221), .A2(n568), .ZN(n531) );
  XNOR2_X1 U642 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U643 ( .A(n781), .B(n533), .ZN(n763) );
  NAND2_X1 U644 ( .A1(G217), .A2(n534), .ZN(n535) );
  OR2_X1 U645 ( .A1(n713), .A2(n712), .ZN(n614) );
  INV_X1 U646 ( .A(n614), .ZN(n710) );
  NAND2_X1 U647 ( .A1(n606), .A2(n710), .ZN(n545) );
  NOR2_X2 U648 ( .A1(G953), .A2(G237), .ZN(n552) );
  NAND2_X1 U649 ( .A1(G210), .A2(n552), .ZN(n536) );
  XNOR2_X1 U650 ( .A(n536), .B(G101), .ZN(n537) );
  XNOR2_X1 U651 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U652 ( .A(n372), .B(n539), .ZN(n541) );
  NAND2_X1 U653 ( .A1(n688), .A2(n543), .ZN(n544) );
  XNOR2_X2 U654 ( .A(n544), .B(G472), .ZN(n603) );
  NOR2_X1 U655 ( .A1(n545), .A2(n377), .ZN(n546) );
  NAND2_X1 U656 ( .A1(n617), .A2(n546), .ZN(n547) );
  XNOR2_X1 U657 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n562) );
  XNOR2_X1 U658 ( .A(n611), .B(G131), .ZN(n548) );
  XNOR2_X1 U659 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U660 ( .A(n551), .B(n550), .ZN(n560) );
  NAND2_X1 U661 ( .A1(G214), .A2(n552), .ZN(n553) );
  XNOR2_X1 U662 ( .A(n554), .B(n553), .ZN(n558) );
  XNOR2_X1 U663 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U664 ( .A(n558), .B(n557), .Z(n559) );
  XNOR2_X1 U665 ( .A(n560), .B(n559), .ZN(n683) );
  NOR2_X1 U666 ( .A1(G902), .A2(n683), .ZN(n561) );
  XNOR2_X1 U667 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U668 ( .A(n563), .B(G475), .ZN(n608) );
  XNOR2_X1 U669 ( .A(n565), .B(n564), .ZN(n567) );
  NAND2_X1 U670 ( .A1(G217), .A2(n568), .ZN(n569) );
  XNOR2_X1 U671 ( .A(n572), .B(n571), .ZN(n759) );
  NOR2_X1 U672 ( .A1(G902), .A2(n759), .ZN(n573) );
  INV_X1 U673 ( .A(n573), .ZN(n574) );
  INV_X1 U674 ( .A(n607), .ZN(n583) );
  NAND2_X1 U675 ( .A1(n608), .A2(n583), .ZN(n576) );
  INV_X1 U676 ( .A(KEYINPUT104), .ZN(n575) );
  INV_X1 U677 ( .A(KEYINPUT110), .ZN(n577) );
  INV_X1 U678 ( .A(n698), .ZN(n581) );
  NAND2_X1 U679 ( .A1(n447), .A2(n581), .ZN(n578) );
  XNOR2_X1 U680 ( .A(n578), .B(G104), .ZN(G6) );
  NAND2_X1 U681 ( .A1(n635), .A2(n710), .ZN(n579) );
  INV_X1 U682 ( .A(n603), .ZN(n651) );
  NAND2_X1 U683 ( .A1(n617), .A2(n720), .ZN(n580) );
  XNOR2_X1 U684 ( .A(n582), .B(G113), .ZN(G15) );
  OR2_X1 U685 ( .A1(n608), .A2(n583), .ZN(n695) );
  INV_X1 U686 ( .A(n695), .ZN(n690) );
  XNOR2_X1 U687 ( .A(n584), .B(G116), .ZN(G18) );
  INV_X1 U688 ( .A(n635), .ZN(n672) );
  XNOR2_X1 U689 ( .A(n603), .B(KEYINPUT6), .ZN(n613) );
  NOR2_X1 U690 ( .A1(G900), .A2(n585), .ZN(n586) );
  NOR2_X1 U691 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U692 ( .A1(n713), .A2(n588), .ZN(n605) );
  NAND2_X1 U693 ( .A1(n712), .A2(n605), .ZN(n650) );
  NOR2_X1 U694 ( .A1(n613), .A2(n650), .ZN(n589) );
  XNOR2_X1 U695 ( .A(n589), .B(KEYINPUT111), .ZN(n590) );
  NOR2_X2 U696 ( .A1(n698), .A2(n590), .ZN(n666) );
  NAND2_X1 U697 ( .A1(n666), .A2(n726), .ZN(n591) );
  XOR2_X1 U698 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n592) );
  XNOR2_X1 U699 ( .A(n593), .B(n592), .ZN(n594) );
  NAND2_X1 U700 ( .A1(n594), .A2(n646), .ZN(n675) );
  XNOR2_X1 U701 ( .A(G140), .B(KEYINPUT118), .ZN(n595) );
  XNOR2_X1 U702 ( .A(n675), .B(n595), .ZN(G42) );
  NOR2_X1 U703 ( .A1(n608), .A2(n607), .ZN(n647) );
  INV_X1 U704 ( .A(n713), .ZN(n596) );
  NAND2_X1 U705 ( .A1(n647), .A2(n596), .ZN(n597) );
  NOR2_X2 U706 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U707 ( .A(n599), .B(KEYINPUT22), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n629), .A2(n613), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(KEYINPUT85), .ZN(n601) );
  NOR2_X1 U710 ( .A1(n353), .A2(n712), .ZN(n600) );
  XOR2_X1 U711 ( .A(n378), .B(G101), .Z(G3) );
  NAND2_X1 U712 ( .A1(n603), .A2(n726), .ZN(n604) );
  INV_X1 U713 ( .A(n606), .ZN(n653) );
  NAND2_X1 U714 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U715 ( .A(n609), .B(KEYINPUT109), .ZN(n620) );
  NAND2_X1 U716 ( .A1(n655), .A2(n620), .ZN(n610) );
  NOR2_X1 U717 ( .A1(n646), .A2(n610), .ZN(n661) );
  INV_X1 U718 ( .A(n611), .ZN(n612) );
  XNOR2_X1 U719 ( .A(n661), .B(n612), .ZN(G45) );
  XNOR2_X1 U720 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n616) );
  INV_X1 U721 ( .A(KEYINPUT108), .ZN(n615) );
  XOR2_X1 U722 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n618) );
  XNOR2_X1 U723 ( .A(n619), .B(n618), .ZN(n621) );
  NAND2_X1 U724 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U725 ( .A1(n790), .A2(KEYINPUT44), .ZN(n624) );
  OR2_X1 U726 ( .A1(n657), .A2(n690), .ZN(n623) );
  INV_X1 U727 ( .A(n623), .ZN(n725) );
  NOR2_X2 U728 ( .A1(n626), .A2(n625), .ZN(n628) );
  INV_X1 U729 ( .A(KEYINPUT87), .ZN(n627) );
  XNOR2_X1 U730 ( .A(n628), .B(n627), .ZN(n637) );
  BUF_X1 U731 ( .A(n629), .Z(n631) );
  NOR2_X1 U732 ( .A1(n377), .A2(n353), .ZN(n630) );
  NAND2_X1 U733 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U734 ( .A1(n632), .A2(n400), .ZN(n633) );
  XNOR2_X1 U735 ( .A(n633), .B(KEYINPUT107), .ZN(n791) );
  NAND2_X1 U736 ( .A1(n641), .A2(KEYINPUT44), .ZN(n636) );
  NAND2_X1 U737 ( .A1(n637), .A2(n636), .ZN(n639) );
  NOR2_X1 U738 ( .A1(n381), .A2(KEYINPUT44), .ZN(n640) );
  XNOR2_X1 U739 ( .A(n640), .B(KEYINPUT67), .ZN(n643) );
  XNOR2_X1 U740 ( .A(n641), .B(KEYINPUT88), .ZN(n642) );
  XNOR2_X2 U741 ( .A(n644), .B(KEYINPUT45), .ZN(n766) );
  XOR2_X1 U742 ( .A(KEYINPUT38), .B(KEYINPUT75), .Z(n645) );
  INV_X1 U743 ( .A(n647), .ZN(n729) );
  NAND2_X1 U744 ( .A1(n709), .A2(n662), .ZN(n654) );
  XOR2_X1 U745 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n656) );
  NAND2_X1 U746 ( .A1(n674), .A2(n657), .ZN(n659) );
  XOR2_X1 U747 ( .A(KEYINPUT113), .B(KEYINPUT40), .Z(n658) );
  XOR2_X1 U748 ( .A(n661), .B(KEYINPUT82), .Z(n665) );
  XNOR2_X1 U749 ( .A(n663), .B(KEYINPUT47), .ZN(n664) );
  XOR2_X1 U750 ( .A(n666), .B(KEYINPUT114), .Z(n668) );
  NOR2_X1 U751 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n674), .A2(n690), .ZN(n704) );
  NAND2_X1 U753 ( .A1(n388), .A2(KEYINPUT2), .ZN(n677) );
  NOR2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n679) );
  AND2_X1 U755 ( .A1(n766), .A2(n679), .ZN(n708) );
  BUF_X1 U756 ( .A(n708), .Z(n680) );
  XNOR2_X1 U757 ( .A(KEYINPUT65), .B(KEYINPUT124), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n681), .B(KEYINPUT59), .ZN(n682) );
  INV_X1 U759 ( .A(G952), .ZN(n685) );
  XNOR2_X1 U760 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n686) );
  XOR2_X1 U761 ( .A(KEYINPUT116), .B(KEYINPUT62), .Z(n687) );
  NAND2_X1 U762 ( .A1(n447), .A2(n690), .ZN(n693) );
  XOR2_X1 U763 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n692) );
  XNOR2_X1 U764 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U765 ( .A(G107), .B(n694), .ZN(G9) );
  NOR2_X1 U766 ( .A1(n699), .A2(n695), .ZN(n697) );
  XNOR2_X1 U767 ( .A(G128), .B(KEYINPUT29), .ZN(n696) );
  XNOR2_X1 U768 ( .A(n697), .B(n696), .ZN(G30) );
  NOR2_X1 U769 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U770 ( .A(G146), .B(KEYINPUT117), .ZN(n700) );
  XNOR2_X1 U771 ( .A(n701), .B(n700), .ZN(G48) );
  XNOR2_X1 U772 ( .A(n702), .B(G125), .ZN(n703) );
  XNOR2_X1 U773 ( .A(n703), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U774 ( .A(G134), .B(n704), .ZN(G36) );
  INV_X1 U775 ( .A(n782), .ZN(n706) );
  AND2_X1 U776 ( .A1(n766), .A2(n706), .ZN(n707) );
  NOR2_X1 U777 ( .A1(n353), .A2(n710), .ZN(n711) );
  XOR2_X1 U778 ( .A(KEYINPUT50), .B(n711), .Z(n717) );
  NAND2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U780 ( .A(n714), .B(KEYINPUT49), .ZN(n715) );
  XNOR2_X1 U781 ( .A(KEYINPUT119), .B(n715), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U783 ( .A1(n377), .A2(n718), .ZN(n719) );
  NOR2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U785 ( .A(KEYINPUT51), .B(n721), .ZN(n722) );
  NAND2_X1 U786 ( .A1(n739), .A2(n722), .ZN(n734) );
  BUF_X1 U787 ( .A(n723), .Z(n738) );
  NOR2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n731) );
  NOR2_X1 U789 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U790 ( .A1(n729), .A2(n728), .ZN(n730) );
  OR2_X1 U791 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U792 ( .A1(n738), .A2(n732), .ZN(n733) );
  NAND2_X1 U793 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U794 ( .A(KEYINPUT52), .B(n735), .Z(n736) );
  NOR2_X1 U795 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U796 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U797 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U798 ( .A(KEYINPUT53), .B(n743), .ZN(G75) );
  NAND2_X1 U799 ( .A1(n431), .A2(G210), .ZN(n749) );
  XOR2_X1 U800 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n745) );
  XNOR2_X1 U801 ( .A(n745), .B(KEYINPUT55), .ZN(n746) );
  XNOR2_X1 U802 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X2 U803 ( .A1(n750), .A2(n765), .ZN(n751) );
  XNOR2_X1 U804 ( .A(n751), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U805 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n754) );
  XNOR2_X1 U806 ( .A(n382), .B(KEYINPUT123), .ZN(n753) );
  XNOR2_X1 U807 ( .A(n754), .B(n753), .ZN(n756) );
  NAND2_X1 U808 ( .A1(n431), .A2(G469), .ZN(n755) );
  XOR2_X1 U809 ( .A(n756), .B(n755), .Z(n757) );
  NOR2_X1 U810 ( .A1(n765), .A2(n757), .ZN(G54) );
  NAND2_X1 U811 ( .A1(n380), .A2(G478), .ZN(n760) );
  XNOR2_X1 U812 ( .A(n760), .B(n759), .ZN(n761) );
  NOR2_X1 U813 ( .A1(n765), .A2(n761), .ZN(G63) );
  NAND2_X1 U814 ( .A1(n380), .A2(G217), .ZN(n762) );
  XNOR2_X1 U815 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U816 ( .A1(n765), .A2(n764), .ZN(G66) );
  BUF_X1 U817 ( .A(n766), .Z(n767) );
  NAND2_X1 U818 ( .A1(n767), .A2(n783), .ZN(n771) );
  NAND2_X1 U819 ( .A1(G953), .A2(G224), .ZN(n768) );
  XNOR2_X1 U820 ( .A(KEYINPUT61), .B(n768), .ZN(n769) );
  NAND2_X1 U821 ( .A1(n769), .A2(G898), .ZN(n770) );
  NAND2_X1 U822 ( .A1(n771), .A2(n770), .ZN(n778) );
  XNOR2_X1 U823 ( .A(n772), .B(KEYINPUT127), .ZN(n773) );
  XOR2_X1 U824 ( .A(n774), .B(n773), .Z(n776) );
  NOR2_X1 U825 ( .A1(G898), .A2(n783), .ZN(n775) );
  NOR2_X1 U826 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U827 ( .A(n778), .B(n777), .ZN(n779) );
  XNOR2_X1 U828 ( .A(KEYINPUT126), .B(n779), .ZN(G69) );
  XNOR2_X1 U829 ( .A(n780), .B(n781), .ZN(n785) );
  XNOR2_X1 U830 ( .A(n785), .B(n782), .ZN(n784) );
  NAND2_X1 U831 ( .A1(n784), .A2(n783), .ZN(n789) );
  XNOR2_X1 U832 ( .A(G227), .B(n785), .ZN(n786) );
  NAND2_X1 U833 ( .A1(n786), .A2(G900), .ZN(n787) );
  NAND2_X1 U834 ( .A1(n787), .A2(G953), .ZN(n788) );
  NAND2_X1 U835 ( .A1(n789), .A2(n788), .ZN(G72) );
  XOR2_X1 U836 ( .A(G122), .B(n381), .Z(G24) );
  XNOR2_X1 U837 ( .A(G110), .B(n791), .ZN(G12) );
  XNOR2_X1 U838 ( .A(G119), .B(n792), .ZN(G21) );
  XNOR2_X1 U839 ( .A(n793), .B(G137), .ZN(G39) );
  XNOR2_X1 U840 ( .A(G131), .B(n794), .ZN(G33) );
endmodule

