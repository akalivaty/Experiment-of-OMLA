

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n703, n704, n705, n706, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n813) );
  INV_X2 U556 ( .A(n724), .ZN(n722) );
  NOR2_X1 U557 ( .A1(n708), .A2(n812), .ZN(n710) );
  OR2_X1 U558 ( .A1(n706), .A2(n705), .ZN(n708) );
  AND2_X2 U559 ( .A1(n546), .A2(n545), .ZN(G164) );
  NAND2_X1 U560 ( .A1(n525), .A2(n992), .ZN(n781) );
  XNOR2_X1 U561 ( .A(n764), .B(n523), .ZN(n784) );
  NAND2_X1 U562 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U563 ( .A1(n795), .A2(n526), .ZN(n831) );
  NAND2_X1 U564 ( .A1(n536), .A2(n535), .ZN(n537) );
  INV_X1 U565 ( .A(G2105), .ZN(n536) );
  NOR2_X1 U566 ( .A1(n830), .A2(n524), .ZN(n522) );
  XOR2_X1 U567 ( .A(KEYINPUT32), .B(KEYINPUT108), .Z(n523) );
  AND2_X1 U568 ( .A1(n1010), .A2(n844), .ZN(n524) );
  OR2_X1 U569 ( .A1(n780), .A2(n792), .ZN(n525) );
  AND2_X1 U570 ( .A1(n794), .A2(n793), .ZN(n526) );
  NOR2_X1 U571 ( .A1(n714), .A2(n995), .ZN(n721) );
  OR2_X1 U572 ( .A1(n737), .A2(n736), .ZN(n738) );
  INV_X1 U573 ( .A(KEYINPUT29), .ZN(n740) );
  XNOR2_X1 U574 ( .A(n741), .B(n740), .ZN(n745) );
  NOR2_X1 U575 ( .A1(n706), .A2(n703), .ZN(n704) );
  INV_X1 U576 ( .A(G2104), .ZN(n535) );
  INV_X1 U577 ( .A(KEYINPUT0), .ZN(n547) );
  AND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n912) );
  INV_X1 U579 ( .A(n549), .ZN(n667) );
  XNOR2_X1 U580 ( .A(n547), .B(G543), .ZN(n659) );
  INV_X1 U581 ( .A(KEYINPUT23), .ZN(n528) );
  XNOR2_X2 U582 ( .A(G2104), .B(KEYINPUT67), .ZN(n532) );
  NOR2_X4 U583 ( .A1(G2105), .A2(n532), .ZN(n907) );
  AND2_X1 U584 ( .A1(G101), .A2(n907), .ZN(n527) );
  XNOR2_X1 U585 ( .A(n528), .B(n527), .ZN(n531) );
  NAND2_X1 U586 ( .A1(G113), .A2(n912), .ZN(n529) );
  XOR2_X1 U587 ( .A(KEYINPUT68), .B(n529), .Z(n530) );
  NOR2_X1 U588 ( .A1(n531), .A2(n530), .ZN(n534) );
  AND2_X2 U589 ( .A1(n532), .A2(G2105), .ZN(n910) );
  NAND2_X1 U590 ( .A1(n910), .A2(G125), .ZN(n533) );
  AND2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n540) );
  XNOR2_X2 U592 ( .A(n537), .B(KEYINPUT17), .ZN(n906) );
  NAND2_X1 U593 ( .A1(G137), .A2(n906), .ZN(n538) );
  XOR2_X1 U594 ( .A(KEYINPUT69), .B(n538), .Z(n539) );
  AND2_X2 U595 ( .A1(n540), .A2(n539), .ZN(G160) );
  NAND2_X1 U596 ( .A1(G138), .A2(n906), .ZN(n546) );
  AND2_X1 U597 ( .A1(G126), .A2(n910), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G114), .A2(n912), .ZN(n542) );
  NAND2_X1 U599 ( .A1(G102), .A2(n907), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G108), .ZN(G238) );
  INV_X1 U604 ( .A(G120), .ZN(G236) );
  INV_X1 U605 ( .A(G57), .ZN(G237) );
  INV_X1 U606 ( .A(G132), .ZN(G219) );
  INV_X1 U607 ( .A(G82), .ZN(G220) );
  NOR2_X1 U608 ( .A1(G651), .A2(n659), .ZN(n548) );
  XNOR2_X1 U609 ( .A(KEYINPUT66), .B(n548), .ZN(n598) );
  INV_X1 U610 ( .A(n598), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n667), .A2(G52), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n550), .B(KEYINPUT73), .ZN(n560) );
  NOR2_X1 U613 ( .A1(G651), .A2(G543), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT65), .B(n551), .Z(n662) );
  NAND2_X1 U615 ( .A1(G90), .A2(n662), .ZN(n553) );
  INV_X1 U616 ( .A(G651), .ZN(n555) );
  NOR2_X1 U617 ( .A1(n659), .A2(n555), .ZN(n663) );
  NAND2_X1 U618 ( .A1(G77), .A2(n663), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT9), .ZN(n558) );
  NOR2_X1 U621 ( .A1(G543), .A2(n555), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT1), .B(n556), .Z(n666) );
  NAND2_X1 U623 ( .A1(G64), .A2(n666), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(G171) );
  INV_X1 U626 ( .A(G171), .ZN(G301) );
  NAND2_X1 U627 ( .A1(G91), .A2(n662), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G78), .A2(n663), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U630 ( .A1(G65), .A2(n666), .ZN(n564) );
  NAND2_X1 U631 ( .A1(G53), .A2(n667), .ZN(n563) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT74), .B(n567), .Z(G299) );
  NAND2_X1 U635 ( .A1(n666), .A2(G63), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT81), .B(n568), .Z(n570) );
  NAND2_X1 U637 ( .A1(G51), .A2(n667), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT82), .B(KEYINPUT6), .Z(n571) );
  XOR2_X1 U640 ( .A(n572), .B(n571), .Z(n580) );
  NAND2_X1 U641 ( .A1(n663), .A2(G76), .ZN(n573) );
  XOR2_X1 U642 ( .A(KEYINPUT80), .B(n573), .Z(n577) );
  NAND2_X1 U643 ( .A1(G89), .A2(n662), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT79), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n575), .B(KEYINPUT4), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U647 ( .A(KEYINPUT5), .B(n578), .ZN(n579) );
  NOR2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n581), .B(KEYINPUT83), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n582), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G567), .ZN(n696) );
  NOR2_X1 U655 ( .A1(G223), .A2(n696), .ZN(n584) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n584), .Z(n585) );
  XNOR2_X1 U657 ( .A(KEYINPUT75), .B(n585), .ZN(G234) );
  NAND2_X1 U658 ( .A1(n662), .A2(G81), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G68), .A2(n663), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT13), .B(KEYINPUT76), .Z(n589) );
  XNOR2_X1 U663 ( .A(n590), .B(n589), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n666), .A2(G56), .ZN(n591) );
  XOR2_X1 U665 ( .A(KEYINPUT14), .B(n591), .Z(n592) );
  NOR2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G43), .A2(n667), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n995) );
  INV_X1 U669 ( .A(G860), .ZN(n637) );
  OR2_X1 U670 ( .A1(n995), .A2(n637), .ZN(G153) );
  NAND2_X1 U671 ( .A1(G66), .A2(n666), .ZN(n597) );
  NAND2_X1 U672 ( .A1(G92), .A2(n662), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G54), .A2(n598), .ZN(n599) );
  XNOR2_X1 U675 ( .A(KEYINPUT77), .B(n599), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G79), .A2(n663), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT15), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT78), .B(n605), .ZN(n921) );
  INV_X1 U681 ( .A(n921), .ZN(n1000) );
  NOR2_X1 U682 ( .A1(n1000), .A2(G868), .ZN(n607) );
  INV_X1 U683 ( .A(G868), .ZN(n681) );
  NOR2_X1 U684 ( .A1(n681), .A2(G301), .ZN(n606) );
  NOR2_X1 U685 ( .A1(n607), .A2(n606), .ZN(G284) );
  NOR2_X1 U686 ( .A1(G286), .A2(n681), .ZN(n608) );
  XNOR2_X1 U687 ( .A(n608), .B(KEYINPUT84), .ZN(n610) );
  NOR2_X1 U688 ( .A1(G299), .A2(G868), .ZN(n609) );
  NOR2_X1 U689 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n637), .A2(G559), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n611), .A2(n921), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT85), .ZN(n613) );
  XOR2_X1 U693 ( .A(KEYINPUT16), .B(n613), .Z(G148) );
  NOR2_X1 U694 ( .A1(G868), .A2(n995), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n921), .A2(G868), .ZN(n614) );
  NOR2_X1 U696 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U697 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G135), .A2(n906), .ZN(n618) );
  NAND2_X1 U699 ( .A1(G111), .A2(n912), .ZN(n617) );
  NAND2_X1 U700 ( .A1(n618), .A2(n617), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G99), .A2(n907), .ZN(n619) );
  XNOR2_X1 U702 ( .A(n619), .B(KEYINPUT86), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G123), .A2(n910), .ZN(n620) );
  XNOR2_X1 U704 ( .A(n620), .B(KEYINPUT18), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n949) );
  XNOR2_X1 U707 ( .A(n949), .B(G2096), .ZN(n626) );
  INV_X1 U708 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U710 ( .A1(G67), .A2(n666), .ZN(n627) );
  XNOR2_X1 U711 ( .A(n627), .B(KEYINPUT88), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n667), .A2(G55), .ZN(n628) );
  XOR2_X1 U713 ( .A(KEYINPUT89), .B(n628), .Z(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G93), .A2(n662), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G80), .A2(n663), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U718 ( .A(KEYINPUT87), .B(n633), .Z(n634) );
  OR2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n680) );
  XNOR2_X1 U720 ( .A(n680), .B(KEYINPUT90), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n921), .A2(G559), .ZN(n636) );
  XOR2_X1 U722 ( .A(n995), .B(n636), .Z(n678) );
  NAND2_X1 U723 ( .A1(n678), .A2(n637), .ZN(n638) );
  XNOR2_X1 U724 ( .A(n639), .B(n638), .ZN(G145) );
  NAND2_X1 U725 ( .A1(G47), .A2(n667), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n666), .A2(G60), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U728 ( .A(n642), .B(KEYINPUT71), .ZN(n647) );
  NAND2_X1 U729 ( .A1(G85), .A2(n662), .ZN(n644) );
  NAND2_X1 U730 ( .A1(G72), .A2(n663), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U732 ( .A(KEYINPUT70), .B(n645), .Z(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U734 ( .A(n648), .B(KEYINPUT72), .ZN(G290) );
  NAND2_X1 U735 ( .A1(G61), .A2(n666), .ZN(n650) );
  NAND2_X1 U736 ( .A1(G86), .A2(n662), .ZN(n649) );
  NAND2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U738 ( .A1(n663), .A2(G73), .ZN(n651) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(n651), .Z(n652) );
  NOR2_X1 U740 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U741 ( .A1(G48), .A2(n667), .ZN(n654) );
  NAND2_X1 U742 ( .A1(n655), .A2(n654), .ZN(G305) );
  NAND2_X1 U743 ( .A1(G651), .A2(G74), .ZN(n657) );
  NAND2_X1 U744 ( .A1(G49), .A2(n667), .ZN(n656) );
  NAND2_X1 U745 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U746 ( .A1(n666), .A2(n658), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n659), .A2(G87), .ZN(n660) );
  NAND2_X1 U748 ( .A1(n661), .A2(n660), .ZN(G288) );
  NAND2_X1 U749 ( .A1(G88), .A2(n662), .ZN(n665) );
  NAND2_X1 U750 ( .A1(G75), .A2(n663), .ZN(n664) );
  NAND2_X1 U751 ( .A1(n665), .A2(n664), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G62), .A2(n666), .ZN(n669) );
  NAND2_X1 U753 ( .A1(G50), .A2(n667), .ZN(n668) );
  NAND2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U755 ( .A1(n671), .A2(n670), .ZN(G166) );
  XOR2_X1 U756 ( .A(G290), .B(n680), .Z(n677) );
  XOR2_X1 U757 ( .A(KEYINPUT91), .B(KEYINPUT19), .Z(n672) );
  XNOR2_X1 U758 ( .A(G288), .B(n672), .ZN(n673) );
  XNOR2_X1 U759 ( .A(G305), .B(n673), .ZN(n675) );
  XNOR2_X1 U760 ( .A(G166), .B(G299), .ZN(n674) );
  XNOR2_X1 U761 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n677), .B(n676), .ZN(n923) );
  XNOR2_X1 U763 ( .A(n678), .B(n923), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n679), .A2(G868), .ZN(n683) );
  NAND2_X1 U765 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n683), .A2(n682), .ZN(G295) );
  NAND2_X1 U767 ( .A1(G2078), .A2(G2084), .ZN(n684) );
  XOR2_X1 U768 ( .A(KEYINPUT20), .B(n684), .Z(n685) );
  NAND2_X1 U769 ( .A1(G2090), .A2(n685), .ZN(n686) );
  XNOR2_X1 U770 ( .A(KEYINPUT21), .B(n686), .ZN(n687) );
  NAND2_X1 U771 ( .A1(n687), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U772 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n688) );
  XNOR2_X1 U774 ( .A(KEYINPUT22), .B(n688), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n689), .A2(G96), .ZN(n690) );
  NOR2_X1 U776 ( .A1(G218), .A2(n690), .ZN(n691) );
  XNOR2_X1 U777 ( .A(KEYINPUT92), .B(n691), .ZN(n855) );
  INV_X1 U778 ( .A(n855), .ZN(n692) );
  NAND2_X1 U779 ( .A1(n692), .A2(G2106), .ZN(n693) );
  XNOR2_X1 U780 ( .A(n693), .B(KEYINPUT93), .ZN(n698) );
  NOR2_X1 U781 ( .A1(G236), .A2(G238), .ZN(n694) );
  NAND2_X1 U782 ( .A1(G69), .A2(n694), .ZN(n695) );
  NOR2_X1 U783 ( .A1(G237), .A2(n695), .ZN(n856) );
  NOR2_X1 U784 ( .A1(n696), .A2(n856), .ZN(n697) );
  NOR2_X1 U785 ( .A1(n698), .A2(n697), .ZN(G319) );
  NAND2_X1 U786 ( .A1(G483), .A2(G661), .ZN(n700) );
  INV_X1 U787 ( .A(G319), .ZN(n699) );
  NOR2_X1 U788 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U789 ( .A(n701), .B(KEYINPUT94), .ZN(n854) );
  NAND2_X1 U790 ( .A1(G36), .A2(n854), .ZN(G176) );
  INV_X1 U791 ( .A(G166), .ZN(G303) );
  INV_X1 U792 ( .A(n813), .ZN(n706) );
  INV_X1 U793 ( .A(G40), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(G160), .ZN(n724) );
  NAND2_X1 U795 ( .A1(G8), .A2(n724), .ZN(n792) );
  INV_X1 U796 ( .A(G1996), .ZN(n705) );
  NAND2_X1 U797 ( .A1(G160), .A2(G40), .ZN(n812) );
  XOR2_X1 U798 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n709) );
  XNOR2_X1 U799 ( .A(n710), .B(n709), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n724), .A2(G1341), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U802 ( .A(KEYINPUT104), .B(n713), .ZN(n714) );
  NAND2_X1 U803 ( .A1(n721), .A2(n921), .ZN(n719) );
  INV_X1 U804 ( .A(G1348), .ZN(n1017) );
  NOR2_X1 U805 ( .A1(n722), .A2(n1017), .ZN(n715) );
  XNOR2_X1 U806 ( .A(n715), .B(KEYINPUT105), .ZN(n717) );
  NAND2_X1 U807 ( .A1(n722), .A2(G2067), .ZN(n716) );
  NAND2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U810 ( .A(n720), .B(KEYINPUT106), .ZN(n732) );
  OR2_X1 U811 ( .A1(n721), .A2(n921), .ZN(n730) );
  NAND2_X1 U812 ( .A1(n722), .A2(G2072), .ZN(n723) );
  XNOR2_X1 U813 ( .A(KEYINPUT27), .B(n723), .ZN(n727) );
  AND2_X1 U814 ( .A1(G1956), .A2(n724), .ZN(n725) );
  XNOR2_X1 U815 ( .A(KEYINPUT102), .B(n725), .ZN(n726) );
  NOR2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n734) );
  INV_X1 U817 ( .A(G299), .ZN(n735) );
  NOR2_X1 U818 ( .A1(n734), .A2(n735), .ZN(n729) );
  XNOR2_X1 U819 ( .A(KEYINPUT103), .B(KEYINPUT28), .ZN(n728) );
  XNOR2_X1 U820 ( .A(n729), .B(n728), .ZN(n733) );
  AND2_X1 U821 ( .A1(n730), .A2(n733), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n739) );
  INV_X1 U823 ( .A(n733), .ZN(n737) );
  NAND2_X1 U824 ( .A1(n734), .A2(n735), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n741) );
  XOR2_X1 U826 ( .A(KEYINPUT25), .B(G2078), .Z(n975) );
  INV_X1 U827 ( .A(n722), .ZN(n756) );
  NOR2_X1 U828 ( .A1(n975), .A2(n756), .ZN(n743) );
  NOR2_X1 U829 ( .A1(n722), .A2(G1961), .ZN(n742) );
  NOR2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n746) );
  NOR2_X1 U831 ( .A1(G301), .A2(n746), .ZN(n744) );
  NOR2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n754) );
  AND2_X1 U833 ( .A1(G301), .A2(n746), .ZN(n751) );
  NOR2_X1 U834 ( .A1(G1966), .A2(n792), .ZN(n768) );
  NOR2_X1 U835 ( .A1(G2084), .A2(n756), .ZN(n765) );
  NOR2_X1 U836 ( .A1(n768), .A2(n765), .ZN(n747) );
  NAND2_X1 U837 ( .A1(G8), .A2(n747), .ZN(n748) );
  XNOR2_X1 U838 ( .A(KEYINPUT30), .B(n748), .ZN(n749) );
  NOR2_X1 U839 ( .A1(G168), .A2(n749), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U841 ( .A(n752), .B(KEYINPUT31), .ZN(n753) );
  NOR2_X2 U842 ( .A1(n754), .A2(n753), .ZN(n766) );
  XNOR2_X1 U843 ( .A(KEYINPUT107), .B(n766), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n755), .A2(G286), .ZN(n763) );
  INV_X1 U845 ( .A(G8), .ZN(n761) );
  NOR2_X1 U846 ( .A1(G1971), .A2(n792), .ZN(n758) );
  NOR2_X1 U847 ( .A1(G2090), .A2(n756), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n759), .A2(G303), .ZN(n760) );
  OR2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n765), .A2(G8), .ZN(n770) );
  XOR2_X1 U852 ( .A(KEYINPUT107), .B(n766), .Z(n767) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n770), .A2(n769), .ZN(n785) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n999) );
  AND2_X1 U856 ( .A1(n785), .A2(n999), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n784), .A2(n771), .ZN(n775) );
  INV_X1 U858 ( .A(n999), .ZN(n773) );
  NOR2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n779) );
  NOR2_X1 U860 ( .A1(G1971), .A2(G303), .ZN(n772) );
  NOR2_X1 U861 ( .A1(n779), .A2(n772), .ZN(n1004) );
  OR2_X1 U862 ( .A1(n773), .A2(n1004), .ZN(n774) );
  AND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U864 ( .A(n776), .B(KEYINPUT109), .Z(n777) );
  NOR2_X1 U865 ( .A1(n792), .A2(n777), .ZN(n778) );
  NOR2_X1 U866 ( .A1(KEYINPUT33), .A2(n778), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n779), .A2(KEYINPUT33), .ZN(n780) );
  XOR2_X1 U868 ( .A(G1981), .B(G305), .Z(n992) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  INV_X1 U870 ( .A(n783), .ZN(n795) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n788) );
  NOR2_X1 U872 ( .A1(G2090), .A2(G303), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G8), .A2(n786), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n789), .A2(n792), .ZN(n794) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n790) );
  XOR2_X1 U877 ( .A(n790), .B(KEYINPUT24), .Z(n791) );
  OR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G119), .A2(n910), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G107), .A2(n912), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U882 ( .A(KEYINPUT99), .B(n798), .ZN(n802) );
  NAND2_X1 U883 ( .A1(G131), .A2(n906), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G95), .A2(n907), .ZN(n799) );
  AND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U886 ( .A1(n802), .A2(n801), .ZN(n886) );
  NAND2_X1 U887 ( .A1(G1991), .A2(n886), .ZN(n811) );
  NAND2_X1 U888 ( .A1(G141), .A2(n906), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G117), .A2(n912), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U891 ( .A1(n907), .A2(G105), .ZN(n805) );
  XOR2_X1 U892 ( .A(KEYINPUT38), .B(n805), .Z(n806) );
  NOR2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n910), .A2(G129), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n809), .A2(n808), .ZN(n891) );
  NAND2_X1 U896 ( .A1(G1996), .A2(n891), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n811), .A2(n810), .ZN(n952) );
  NOR2_X1 U898 ( .A1(n813), .A2(n812), .ZN(n844) );
  NAND2_X1 U899 ( .A1(n952), .A2(n844), .ZN(n814) );
  XOR2_X1 U900 ( .A(KEYINPUT100), .B(n814), .Z(n836) );
  INV_X1 U901 ( .A(n836), .ZN(n827) );
  XNOR2_X1 U902 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n818) );
  NAND2_X1 U903 ( .A1(G140), .A2(n906), .ZN(n816) );
  NAND2_X1 U904 ( .A1(G104), .A2(n907), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U906 ( .A(n818), .B(n817), .ZN(n824) );
  XNOR2_X1 U907 ( .A(KEYINPUT97), .B(KEYINPUT35), .ZN(n822) );
  NAND2_X1 U908 ( .A1(G128), .A2(n910), .ZN(n820) );
  NAND2_X1 U909 ( .A1(G116), .A2(n912), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U911 ( .A(n822), .B(n821), .ZN(n823) );
  NOR2_X1 U912 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U913 ( .A(n825), .B(KEYINPUT36), .ZN(n826) );
  XNOR2_X1 U914 ( .A(n826), .B(KEYINPUT98), .ZN(n889) );
  XNOR2_X1 U915 ( .A(G2067), .B(KEYINPUT37), .ZN(n841) );
  NOR2_X1 U916 ( .A1(n889), .A2(n841), .ZN(n956) );
  NAND2_X1 U917 ( .A1(n844), .A2(n956), .ZN(n839) );
  NAND2_X1 U918 ( .A1(n827), .A2(n839), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT101), .B(n828), .Z(n830) );
  XOR2_X1 U920 ( .A(G1986), .B(G290), .Z(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT95), .B(n829), .ZN(n1010) );
  NAND2_X1 U922 ( .A1(n831), .A2(n522), .ZN(n847) );
  NOR2_X1 U923 ( .A1(G1996), .A2(n891), .ZN(n946) );
  NOR2_X1 U924 ( .A1(G1991), .A2(n886), .ZN(n950) );
  NOR2_X1 U925 ( .A1(G1986), .A2(G290), .ZN(n832) );
  XNOR2_X1 U926 ( .A(KEYINPUT110), .B(n832), .ZN(n833) );
  NOR2_X1 U927 ( .A1(n950), .A2(n833), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT111), .B(n834), .Z(n835) );
  NOR2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U930 ( .A1(n946), .A2(n837), .ZN(n838) );
  XNOR2_X1 U931 ( .A(KEYINPUT39), .B(n838), .ZN(n840) );
  NAND2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n843) );
  NAND2_X1 U933 ( .A1(n841), .A2(n889), .ZN(n842) );
  XNOR2_X1 U934 ( .A(n842), .B(KEYINPUT112), .ZN(n963) );
  NAND2_X1 U935 ( .A1(n843), .A2(n963), .ZN(n845) );
  NAND2_X1 U936 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U937 ( .A1(n847), .A2(n846), .ZN(n850) );
  XOR2_X1 U938 ( .A(KEYINPUT114), .B(KEYINPUT40), .Z(n848) );
  XNOR2_X1 U939 ( .A(KEYINPUT113), .B(n848), .ZN(n849) );
  XNOR2_X1 U940 ( .A(n850), .B(n849), .ZN(G329) );
  INV_X1 U941 ( .A(G223), .ZN(n851) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n851), .ZN(G217) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n852) );
  NAND2_X1 U944 ( .A1(G661), .A2(n852), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n853) );
  NAND2_X1 U946 ( .A1(n854), .A2(n853), .ZN(G188) );
  INV_X1 U948 ( .A(G96), .ZN(G221) );
  NAND2_X1 U949 ( .A1(n856), .A2(n855), .ZN(G261) );
  INV_X1 U950 ( .A(G261), .ZN(G325) );
  XOR2_X1 U951 ( .A(G2100), .B(KEYINPUT118), .Z(n858) );
  XNOR2_X1 U952 ( .A(KEYINPUT117), .B(KEYINPUT43), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2072), .Z(n860) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2090), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U957 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U958 ( .A(G2678), .B(G2096), .ZN(n863) );
  XNOR2_X1 U959 ( .A(n864), .B(n863), .ZN(n866) );
  XOR2_X1 U960 ( .A(G2078), .B(G2084), .Z(n865) );
  XNOR2_X1 U961 ( .A(n866), .B(n865), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1976), .B(G1961), .Z(n868) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1971), .ZN(n867) );
  XNOR2_X1 U964 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U965 ( .A(n869), .B(G2474), .Z(n871) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U968 ( .A(KEYINPUT41), .B(G1981), .Z(n873) );
  XNOR2_X1 U969 ( .A(G1956), .B(G1966), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U971 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U972 ( .A1(n910), .A2(G124), .ZN(n876) );
  XNOR2_X1 U973 ( .A(n876), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G112), .A2(n912), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U976 ( .A1(G136), .A2(n906), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G100), .A2(n907), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U979 ( .A1(n882), .A2(n881), .ZN(G162) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n884) );
  XNOR2_X1 U981 ( .A(G164), .B(KEYINPUT124), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U983 ( .A(G160), .B(n949), .Z(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n905) );
  XOR2_X1 U986 ( .A(n889), .B(G162), .Z(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n903) );
  NAND2_X1 U988 ( .A1(n912), .A2(G118), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT119), .B(n892), .Z(n894) );
  NAND2_X1 U990 ( .A1(n910), .A2(G130), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U992 ( .A(KEYINPUT120), .B(n895), .ZN(n901) );
  NAND2_X1 U993 ( .A1(n907), .A2(G106), .ZN(n896) );
  XOR2_X1 U994 ( .A(KEYINPUT121), .B(n896), .Z(n898) );
  NAND2_X1 U995 ( .A1(n906), .A2(G142), .ZN(n897) );
  NAND2_X1 U996 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(n899), .B(KEYINPUT45), .Z(n900) );
  NOR2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U999 ( .A(n903), .B(n902), .Z(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n919) );
  NAND2_X1 U1001 ( .A1(G139), .A2(n906), .ZN(n909) );
  NAND2_X1 U1002 ( .A1(G103), .A2(n907), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(n917) );
  NAND2_X1 U1004 ( .A1(n910), .A2(G127), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(n911), .B(KEYINPUT122), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(G115), .A2(n912), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1008 ( .A(KEYINPUT47), .B(n915), .Z(n916) );
  NOR2_X1 U1009 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1010 ( .A(KEYINPUT123), .B(n918), .Z(n959) );
  XNOR2_X1 U1011 ( .A(n919), .B(n959), .ZN(n920) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n920), .ZN(G395) );
  XNOR2_X1 U1013 ( .A(G171), .B(n921), .ZN(n922) );
  XNOR2_X1 U1014 ( .A(n922), .B(n995), .ZN(n925) );
  XNOR2_X1 U1015 ( .A(G286), .B(n923), .ZN(n924) );
  XNOR2_X1 U1016 ( .A(n925), .B(n924), .ZN(n926) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n926), .ZN(n927) );
  XOR2_X1 U1018 ( .A(KEYINPUT125), .B(n927), .Z(G397) );
  XNOR2_X1 U1019 ( .A(G2435), .B(G2446), .ZN(n937) );
  XOR2_X1 U1020 ( .A(G2454), .B(G2430), .Z(n929) );
  XNOR2_X1 U1021 ( .A(G2451), .B(G2443), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(n929), .B(n928), .ZN(n933) );
  XOR2_X1 U1023 ( .A(G2427), .B(KEYINPUT115), .Z(n931) );
  XNOR2_X1 U1024 ( .A(G1341), .B(G1348), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(n931), .B(n930), .ZN(n932) );
  XOR2_X1 U1026 ( .A(n933), .B(n932), .Z(n935) );
  XNOR2_X1 U1027 ( .A(KEYINPUT116), .B(G2438), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(n935), .B(n934), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(n937), .B(n936), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(n938), .A2(G14), .ZN(n944) );
  NAND2_X1 U1031 ( .A1(G319), .A2(n944), .ZN(n941) );
  NOR2_X1 U1032 ( .A1(G227), .A2(G229), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(KEYINPUT49), .B(n939), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n943) );
  NOR2_X1 U1035 ( .A1(G395), .A2(G397), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(G225) );
  INV_X1 U1037 ( .A(G225), .ZN(G308) );
  INV_X1 U1038 ( .A(G69), .ZN(G235) );
  INV_X1 U1039 ( .A(n944), .ZN(G401) );
  XOR2_X1 U1040 ( .A(G2090), .B(G162), .Z(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1042 ( .A(KEYINPUT126), .B(n947), .Z(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT51), .B(n948), .ZN(n958) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1045 ( .A(G160), .B(G2084), .Z(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n966) );
  XOR2_X1 U1050 ( .A(G2072), .B(n959), .Z(n961) );
  XOR2_X1 U1051 ( .A(G164), .B(G2078), .Z(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(KEYINPUT50), .B(n962), .ZN(n964) );
  NAND2_X1 U1054 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1055 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(KEYINPUT52), .B(n967), .ZN(n968) );
  INV_X1 U1057 ( .A(KEYINPUT55), .ZN(n988) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n988), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(n969), .A2(G29), .ZN(n1043) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(G34), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(n970), .B(KEYINPUT127), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(G2084), .B(n971), .ZN(n986) );
  XNOR2_X1 U1063 ( .A(G2090), .B(G35), .ZN(n984) );
  XOR2_X1 U1064 ( .A(G1991), .B(G25), .Z(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(G28), .ZN(n981) );
  XNOR2_X1 U1066 ( .A(G1996), .B(G32), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(G33), .B(G2072), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(G2067), .B(G26), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(G27), .B(n975), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(KEYINPUT53), .B(n982), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(n988), .B(n987), .ZN(n990) );
  INV_X1 U1078 ( .A(G29), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(G11), .A2(n991), .ZN(n1041) );
  XNOR2_X1 U1081 ( .A(G16), .B(KEYINPUT56), .ZN(n1014) );
  XNOR2_X1 U1082 ( .A(G168), .B(G1966), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT57), .ZN(n1012) );
  XNOR2_X1 U1085 ( .A(G301), .B(G1961), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n995), .B(G1341), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n1008) );
  NAND2_X1 U1088 ( .A1(G1971), .A2(G303), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(G299), .B(G1956), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1000), .B(G1348), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1039) );
  INV_X1 U1099 ( .A(G16), .ZN(n1037) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G5), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1027) );
  XNOR2_X1 U1103 ( .A(KEYINPUT59), .B(G4), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(n1018), .B(n1017), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(G20), .B(G1956), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1024) );
  XNOR2_X1 U1107 ( .A(G1341), .B(G19), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(G1981), .B(G6), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(KEYINPUT60), .B(n1025), .Z(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1034) );
  XNOR2_X1 U1113 ( .A(G1971), .B(G22), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(G23), .B(G1976), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(G1986), .B(G24), .Z(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1118 ( .A(KEYINPUT58), .B(n1032), .ZN(n1033) );
  NOR2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(KEYINPUT61), .B(n1035), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1123 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1124 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

