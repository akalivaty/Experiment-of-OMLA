//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  OR3_X1    g0010(.A1(new_n210), .A2(KEYINPUT64), .A3(G13), .ZN(new_n211));
  OAI21_X1  g0011(.A(KEYINPUT64), .B1(new_n210), .B2(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AND2_X1   g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n203), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n202), .A2(new_n203), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n234), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n235));
  NOR4_X1   g0035(.A1(new_n216), .A2(new_n217), .A3(new_n227), .A4(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT67), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT69), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n256), .B1(new_n210), .B2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n259));
  AND3_X1   g0059(.A1(new_n258), .A2(new_n231), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G1), .B2(new_n232), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G20), .A2(G77), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n257), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT15), .B(G87), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n264), .B1(new_n265), .B2(new_n267), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n259), .A2(new_n231), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n258), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n271), .A2(new_n273), .B1(new_n262), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n263), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n257), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1698), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G232), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n281), .B2(new_n282), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G238), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n281), .A2(new_n282), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n284), .B(new_n287), .C1(new_n207), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  OAI211_X1 g0090(.A(G1), .B(G13), .C1(new_n257), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(G41), .B2(G45), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G274), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n291), .A2(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n298), .B1(new_n300), .B2(G244), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n279), .B1(new_n304), .B2(KEYINPUT70), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT71), .B(G200), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n306), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n305), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n279), .ZN(new_n311));
  AOI21_X1  g0111(.A(G169), .B1(new_n293), .B2(new_n301), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT72), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT72), .ZN(new_n314));
  INV_X1    g0114(.A(new_n302), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n314), .B(new_n279), .C1(new_n315), .C2(G169), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n313), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n322));
  INV_X1    g0122(.A(new_n275), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n203), .A2(G20), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT76), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XOR2_X1   g0125(.A(new_n325), .B(KEYINPUT12), .Z(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n203), .B2(new_n261), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n324), .B1(new_n267), .B2(new_n201), .C1(new_n269), .C2(new_n262), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n273), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n285), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n288), .B(new_n336), .C1(G232), .C2(new_n285), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n292), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n297), .B1(new_n299), .B2(new_n219), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n334), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n291), .B1(new_n337), .B2(new_n338), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n344), .A2(KEYINPUT13), .A3(new_n341), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G169), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT14), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(G179), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n346), .A2(KEYINPUT14), .A3(new_n347), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n333), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(G190), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n332), .C1(new_n354), .C2(new_n346), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n321), .A2(new_n322), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n265), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n276), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n261), .B2(new_n265), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n281), .A2(new_n232), .A3(new_n282), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT7), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n281), .A2(new_n363), .A3(new_n232), .A4(new_n282), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(G68), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(G58), .B(G68), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(G20), .B1(G159), .B2(new_n266), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT16), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n370), .A3(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n360), .B1(new_n372), .B2(new_n273), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n291), .A2(G232), .A3(new_n295), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n374), .A2(new_n297), .ZN(new_n375));
  INV_X1    g0175(.A(G223), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n285), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n335), .A2(G1698), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n377), .B(new_n378), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n292), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n354), .B1(new_n375), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n291), .B1(new_n381), .B2(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n374), .A2(new_n297), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n386), .A2(new_n387), .A3(new_n303), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT77), .B1(new_n373), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n365), .A2(new_n370), .A3(new_n367), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n370), .B1(new_n365), .B2(new_n367), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n273), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n360), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(new_n389), .A3(KEYINPUT77), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT17), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT17), .B1(new_n373), .B2(new_n389), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n393), .A2(new_n394), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n347), .B1(new_n386), .B2(new_n387), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n375), .A2(new_n384), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(G179), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  AOI211_X1 g0206(.A(KEYINPUT18), .B(new_n404), .C1(new_n393), .C2(new_n394), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n397), .A2(new_n399), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n283), .A2(G222), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n410), .A2(KEYINPUT68), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(KEYINPUT68), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n288), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G77), .B1(new_n286), .B2(G223), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n291), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n297), .B1(new_n299), .B2(new_n335), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n308), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  INV_X1    g0219(.A(new_n417), .ZN(new_n420));
  INV_X1    g0220(.A(new_n415), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n411), .B2(new_n412), .ZN(new_n422));
  OAI211_X1 g0222(.A(G190), .B(new_n420), .C1(new_n422), .C2(new_n291), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT10), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n266), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n265), .B2(new_n269), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n273), .B1(new_n201), .B2(new_n277), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n201), .B2(new_n261), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT9), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n431), .ZN(new_n433));
  AND4_X1   g0233(.A1(new_n418), .A2(new_n432), .A3(new_n423), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n418), .A2(new_n432), .A3(new_n423), .A4(new_n433), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n425), .A3(new_n424), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n347), .B1(new_n416), .B2(new_n417), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n317), .B(new_n420), .C1(new_n422), .C2(new_n291), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n430), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n356), .A2(new_n409), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(G244), .B(new_n285), .C1(new_n379), .C2(new_n380), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT4), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n445), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n292), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  AND2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(G257), .A3(new_n291), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT5), .B(G41), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(new_n291), .A3(G274), .A4(new_n452), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n347), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(new_n458), .A3(KEYINPUT79), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT79), .B1(new_n456), .B2(new_n458), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n450), .B(new_n317), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n362), .A2(G107), .A3(new_n364), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n266), .A2(G77), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n207), .A2(KEYINPUT6), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT78), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n206), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT78), .A2(G97), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT6), .B1(new_n208), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(G20), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n467), .A2(new_n468), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n273), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n275), .A2(G20), .B1(new_n294), .B2(G33), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n260), .A2(G97), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n277), .A2(new_n206), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n462), .A2(new_n466), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n232), .B2(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n232), .A2(G33), .A3(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n232), .B(G87), .C1(new_n379), .C2(new_n380), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n288), .A2(new_n494), .A3(new_n232), .A4(G87), .ZN(new_n495));
  AOI211_X1 g0295(.A(KEYINPUT24), .B(new_n491), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n495), .ZN(new_n498));
  INV_X1    g0298(.A(new_n491), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n273), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n479), .A2(new_n258), .A3(new_n272), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n277), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT25), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n276), .B2(G107), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n502), .A2(G107), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G257), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n507));
  OAI211_X1 g0307(.A(G250), .B(new_n285), .C1(new_n379), .C2(new_n380), .ZN(new_n508));
  INV_X1    g0308(.A(G294), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n508), .C1(new_n257), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n292), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n455), .A2(G264), .A3(new_n291), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n458), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n511), .A2(G190), .A3(new_n458), .A4(new_n512), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n501), .A2(new_n506), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n482), .B1(new_n273), .B2(new_n477), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n450), .A2(G190), .A3(new_n460), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT79), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n459), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(new_n463), .B1(new_n449), .B2(new_n292), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n517), .B(new_n518), .C1(new_n521), .C2(new_n354), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n485), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n498), .A2(new_n499), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT24), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n498), .A2(new_n497), .A3(new_n499), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n260), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n506), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n513), .A2(new_n347), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n511), .A2(new_n317), .A3(new_n458), .A4(new_n512), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n523), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G238), .B(new_n285), .C1(new_n379), .C2(new_n380), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT80), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n288), .A2(KEYINPUT80), .A3(G238), .A4(new_n285), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n286), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n291), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n291), .B(G250), .C1(G1), .C2(new_n451), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n452), .A2(G274), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n347), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n270), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(new_n276), .ZN(new_n547));
  AND2_X1   g0347(.A1(KEYINPUT78), .A2(G97), .ZN(new_n548));
  NOR2_X1   g0348(.A1(KEYINPUT78), .A2(G97), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n268), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n288), .A2(new_n232), .A3(G68), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G87), .A2(G107), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n471), .A2(new_n472), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n232), .B1(new_n338), .B2(new_n551), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n552), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n547), .B1(new_n558), .B2(new_n273), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n502), .A2(new_n546), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n544), .ZN(new_n562));
  OAI211_X1 g0362(.A(G244), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n563));
  INV_X1    g0363(.A(G116), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n257), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n537), .B2(new_n538), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n317), .B(new_n562), .C1(new_n566), .C2(new_n291), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n545), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G190), .B(new_n562), .C1(new_n566), .C2(new_n291), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n308), .B1(new_n541), .B2(new_n544), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n558), .A2(new_n273), .ZN(new_n572));
  INV_X1    g0372(.A(new_n547), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n502), .A2(G87), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n570), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n571), .A2(new_n575), .A3(KEYINPUT81), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n568), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n455), .A2(G270), .A3(new_n291), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n581), .A2(new_n458), .ZN(new_n582));
  OAI211_X1 g0382(.A(G264), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n583));
  OAI211_X1 g0383(.A(G257), .B(new_n285), .C1(new_n379), .C2(new_n380), .ZN(new_n584));
  INV_X1    g0384(.A(G303), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n288), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n292), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n347), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT20), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(G33), .B1(new_n471), .B2(new_n472), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n447), .A2(new_n232), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n593), .A2(new_n594), .B1(new_n232), .B2(G116), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n589), .B(new_n592), .C1(new_n595), .C2(new_n260), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n257), .B1(new_n548), .B2(new_n549), .ZN(new_n597));
  INV_X1    g0397(.A(new_n594), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(G20), .B2(new_n564), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(new_n590), .A3(new_n591), .A4(new_n273), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n275), .A2(G20), .A3(new_n564), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n479), .A2(new_n272), .A3(G116), .A4(new_n258), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT82), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT82), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n260), .A2(new_n605), .A3(G116), .A4(new_n479), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n588), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT84), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n604), .A2(new_n606), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(new_n596), .A3(new_n600), .A4(new_n601), .ZN(new_n613));
  AOI211_X1 g0413(.A(new_n347), .B(new_n610), .C1(new_n582), .C2(new_n587), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n582), .A2(new_n587), .A3(G179), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n582), .A2(new_n587), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G190), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n582), .A2(new_n587), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G200), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n619), .A2(new_n620), .A3(new_n612), .A4(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n611), .A2(new_n617), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n534), .A2(new_n580), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n442), .A2(new_n626), .ZN(G372));
  NAND2_X1  g0427(.A1(new_n576), .A2(new_n577), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(new_n579), .A3(new_n569), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n562), .B1(new_n566), .B2(new_n291), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n630), .A2(new_n347), .B1(new_n559), .B2(new_n560), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n567), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n462), .A2(new_n466), .A3(new_n484), .ZN(new_n633));
  XOR2_X1   g0433(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n629), .A2(new_n632), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT85), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n559), .A2(new_n637), .A3(new_n574), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n559), .B2(new_n574), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n571), .B(new_n569), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n633), .A2(new_n640), .A3(new_n632), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT86), .ZN(new_n645));
  INV_X1    g0445(.A(new_n610), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n621), .A2(G169), .A3(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n612), .A2(new_n620), .B1(new_n647), .B2(new_n615), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n613), .B2(new_n588), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n611), .A2(KEYINPUT86), .A3(new_n617), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n533), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n485), .A2(new_n516), .A3(new_n522), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n559), .A2(new_n574), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT85), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n559), .A2(new_n637), .A3(new_n574), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n571), .A2(new_n569), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n657), .A2(new_n658), .B1(new_n631), .B2(new_n567), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n644), .B(new_n632), .C1(new_n652), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n442), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n435), .A2(new_n437), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n393), .A2(new_n394), .A3(new_n389), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT77), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n395), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n398), .B1(new_n668), .B2(KEYINPUT17), .ZN(new_n669));
  AND4_X1   g0469(.A1(new_n313), .A2(new_n355), .A3(new_n316), .A4(new_n318), .ZN(new_n670));
  INV_X1    g0470(.A(new_n352), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n664), .B1(new_n672), .B2(new_n408), .ZN(new_n673));
  INV_X1    g0473(.A(new_n440), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n663), .A2(new_n675), .ZN(G369));
  OAI211_X1 g0476(.A(new_n530), .B(new_n531), .C1(new_n527), .C2(new_n528), .ZN(new_n677));
  OR3_X1    g0477(.A1(new_n323), .A2(KEYINPUT27), .A3(G20), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT27), .B1(new_n323), .B2(G20), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n529), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n516), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n677), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n677), .A2(new_n682), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n624), .B(KEYINPUT89), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n613), .A2(new_n682), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT90), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n650), .A2(new_n651), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n613), .A3(new_n682), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n693), .B1(new_n692), .B2(new_n695), .ZN(new_n698));
  OAI211_X1 g0498(.A(G330), .B(new_n689), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n682), .B1(new_n611), .B2(new_n617), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n688), .B1(new_n686), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n213), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n548), .A2(new_n549), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n564), .A3(new_n554), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n704), .A2(new_n294), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n230), .B2(new_n704), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  NAND3_X1  g0509(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n633), .A2(new_n632), .A3(new_n640), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n710), .A2(new_n634), .B1(new_n711), .B2(KEYINPUT26), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n677), .A2(new_n617), .A3(new_n611), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n653), .A2(new_n713), .A3(new_n659), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n632), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT29), .B(new_n683), .C1(new_n712), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT94), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n635), .B1(new_n580), .B2(new_n633), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n641), .A2(new_n642), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n632), .B(new_n714), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT29), .A4(new_n683), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n724), .B(KEYINPUT29), .C1(new_n661), .C2(new_n683), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n632), .B1(new_n652), .B2(new_n660), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n636), .A2(new_n643), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n683), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT93), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n723), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n534), .A2(new_n580), .A3(new_n625), .A4(new_n683), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n618), .A2(KEYINPUT91), .A3(G179), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT91), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n615), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n541), .A2(new_n544), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n459), .B1(new_n449), .B2(new_n292), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n511), .A2(new_n512), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n734), .A2(new_n735), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n737), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n521), .B1(new_n458), .B2(new_n744), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n742), .A2(new_n618), .A3(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n741), .A2(new_n746), .A3(new_n737), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n682), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n732), .B1(new_n733), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n753), .A2(new_n732), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G330), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n731), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n709), .B1(new_n760), .B2(G1), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT95), .ZN(G364));
  NAND2_X1  g0562(.A1(new_n692), .A2(new_n695), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT90), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n757), .B1(new_n764), .B2(new_n696), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n274), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n294), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n704), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(new_n696), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(G330), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n231), .B1(G20), .B2(new_n347), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n703), .A2(new_n288), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n229), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G45), .B2(new_n249), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n703), .A2(new_n414), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G355), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G116), .B2(new_n213), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n777), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n769), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NAND2_X1  g0586(.A1(G20), .A2(G179), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n303), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n354), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G326), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n786), .A2(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n789), .A2(new_n354), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n232), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n288), .B1(new_n800), .B2(G329), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n303), .A2(G179), .A3(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n232), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n307), .A2(new_n232), .A3(G179), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G190), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n801), .B1(new_n509), .B2(new_n803), .C1(new_n805), .C2(new_n585), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n792), .A2(G200), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G322), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n804), .A2(new_n303), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT98), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT98), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n799), .B(new_n808), .C1(new_n809), .C2(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G50), .A2(new_n793), .B1(new_n790), .B2(G77), .ZN(new_n815));
  INV_X1    g0615(.A(new_n807), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n202), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT97), .ZN(new_n818));
  INV_X1    g0618(.A(new_n797), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n819), .A2(new_n203), .B1(new_n206), .B2(new_n803), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT99), .ZN(new_n821));
  INV_X1    g0621(.A(new_n813), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G107), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(KEYINPUT99), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n800), .A2(G159), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n288), .B1(new_n825), .B2(KEYINPUT32), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n805), .A2(new_n220), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(KEYINPUT32), .C2(new_n825), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n821), .A2(new_n823), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n814), .B1(new_n818), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n785), .B1(new_n830), .B2(new_n776), .ZN(new_n831));
  INV_X1    g0631(.A(new_n775), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n771), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n772), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G396));
  NAND2_X1  g0635(.A1(new_n279), .A2(new_n682), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n319), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n310), .A2(new_n319), .A3(new_n836), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n728), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n683), .B(new_n839), .C1(new_n726), .C2(new_n727), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n769), .B1(new_n759), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n759), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n776), .A2(new_n773), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT100), .Z(new_n847));
  OAI21_X1  g0647(.A(new_n769), .B1(new_n847), .B2(G77), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n564), .A2(new_n791), .B1(new_n819), .B2(new_n809), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G294), .B2(new_n807), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n822), .A2(G87), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n793), .A2(G303), .ZN(new_n852));
  INV_X1    g0652(.A(new_n800), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n414), .B1(new_n803), .B2(new_n206), .C1(new_n786), .C2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n805), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(G107), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n822), .A2(G68), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n288), .B1(new_n803), .B2(new_n202), .C1(new_n859), .C2(new_n853), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G50), .B2(new_n855), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G143), .A2(new_n807), .B1(new_n790), .B2(G159), .ZN(new_n862));
  INV_X1    g0662(.A(G137), .ZN(new_n863));
  INV_X1    g0663(.A(G150), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n863), .B2(new_n794), .C1(new_n864), .C2(new_n819), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT34), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n858), .B(new_n861), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n857), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n848), .B1(new_n869), .B2(new_n776), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n839), .B2(new_n774), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n845), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  OR2_X1    g0673(.A1(new_n473), .A2(new_n475), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n233), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  AOI211_X1 g0678(.A(new_n262), .B(new_n229), .C1(G58), .C2(G68), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n879), .A2(KEYINPUT101), .B1(new_n201), .B2(G68), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n294), .B(G13), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n723), .B(new_n442), .C1(new_n725), .C2(new_n730), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n675), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  INV_X1    g0686(.A(new_n680), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT37), .B1(new_n401), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n401), .A2(new_n405), .ZN(new_n889));
  AND4_X1   g0689(.A1(new_n667), .A2(new_n888), .A3(new_n395), .A4(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n667), .A2(new_n395), .A3(new_n889), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n260), .B1(new_n369), .B2(new_n371), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n887), .B1(new_n892), .B2(new_n360), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT102), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n401), .A2(KEYINPUT102), .A3(new_n887), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n890), .B1(new_n898), .B2(KEYINPUT37), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n669), .B2(new_n408), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n891), .A2(new_n888), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n901), .ZN(new_n904));
  INV_X1    g0704(.A(new_n893), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n409), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT103), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n889), .A2(new_n908), .A3(new_n665), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n909), .A2(new_n893), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n908), .B1(new_n889), .B2(new_n665), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n907), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n904), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n886), .B1(new_n902), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n671), .A2(new_n683), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT102), .B1(new_n401), .B2(new_n887), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n894), .B(new_n680), .C1(new_n393), .C2(new_n394), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n409), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n667), .A2(new_n889), .A3(new_n395), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT37), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n903), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n918), .A2(KEYINPUT39), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n915), .A2(new_n917), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n333), .A2(new_n682), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n352), .A2(new_n355), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n350), .A2(new_n351), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(new_n929), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n319), .A2(new_n682), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n842), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n918), .A2(new_n926), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n680), .B1(new_n406), .B2(new_n407), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n928), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n885), .B(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n890), .A2(KEYINPUT38), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n893), .B1(new_n669), .B2(new_n408), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n909), .A2(new_n893), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT37), .B1(new_n944), .B2(new_n911), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n942), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n946), .A2(new_n926), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n839), .B(new_n932), .C1(new_n754), .C2(new_n755), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT40), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n948), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT40), .B1(new_n918), .B2(new_n926), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n753), .A2(new_n732), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n733), .A2(new_n753), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n954), .B1(new_n955), .B2(new_n732), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n442), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n757), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n957), .B2(new_n953), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n941), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n294), .B2(new_n766), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n941), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n883), .B1(new_n961), .B2(new_n962), .ZN(G367));
  INV_X1    g0763(.A(new_n778), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n245), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n777), .B1(new_n213), .B2(new_n270), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n769), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n855), .A2(G116), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT46), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n786), .A2(new_n794), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G294), .B2(new_n797), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n813), .A2(new_n705), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n288), .B1(new_n800), .B2(G317), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n207), .B2(new_n803), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n968), .B2(new_n969), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G283), .A2(new_n790), .B1(new_n807), .B2(G303), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n971), .A2(new_n972), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(G159), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n201), .A2(new_n791), .B1(new_n819), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G150), .B2(new_n807), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n822), .A2(G77), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n805), .A2(new_n202), .ZN(new_n982));
  INV_X1    g0782(.A(new_n803), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(G68), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(new_n288), .C1(new_n863), .C2(new_n853), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n982), .B(new_n985), .C1(G143), .C2(new_n793), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n977), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n967), .B1(new_n989), .B2(new_n776), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n655), .A2(new_n656), .A3(new_n682), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n659), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n632), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n990), .B1(new_n832), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT45), .ZN(new_n995));
  INV_X1    g0795(.A(new_n701), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n485), .B(new_n522), .C1(new_n517), .C2(new_n683), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n633), .A2(new_n682), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n995), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n996), .A2(new_n1000), .A3(KEYINPUT44), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n701), .B2(new_n999), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT107), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n699), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n765), .A2(new_n1008), .A3(KEYINPUT107), .A4(new_n689), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n689), .A2(new_n700), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n700), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n687), .A2(new_n688), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n765), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n760), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n704), .B(KEYINPUT41), .Z(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n768), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT106), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1016), .A2(new_n999), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(KEYINPUT42), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n485), .B1(new_n997), .B2(new_n677), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT105), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n683), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT42), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1016), .A2(new_n1031), .A3(new_n999), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1025), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT104), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT43), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(KEYINPUT43), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n993), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n699), .A2(new_n1000), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1023), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(KEYINPUT106), .B(new_n1042), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n994), .B1(new_n1022), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT108), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G387));
  INV_X1    g0851(.A(new_n769), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n781), .A2(new_n706), .B1(new_n207), .B2(new_n703), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n706), .C1(G68), .C2(G77), .ZN(new_n1054));
  AOI21_X1  g0854(.A(KEYINPUT50), .B1(new_n357), .B2(new_n201), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n357), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(KEYINPUT109), .A3(new_n778), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n451), .B2(new_n241), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT109), .B1(new_n1057), .B2(new_n778), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1053), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1052), .B1(new_n1061), .B2(new_n777), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n689), .B2(new_n832), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n203), .A2(new_n791), .B1(new_n819), .B2(new_n265), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G50), .B2(new_n807), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n983), .A2(new_n546), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT110), .B(G150), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n414), .B1(new_n800), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n805), .A2(new_n262), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G159), .C2(new_n793), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1065), .B(new_n1071), .C1(new_n206), .C2(new_n813), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G303), .A2(new_n790), .B1(new_n807), .B2(G317), .ZN(new_n1073));
  INV_X1    g0873(.A(G322), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1073), .B1(new_n786), .B2(new_n819), .C1(new_n1074), .C2(new_n794), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT48), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n855), .A2(G294), .B1(G283), .B2(new_n983), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT111), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT49), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n414), .B1(new_n795), .B2(new_n853), .C1(new_n813), .C2(new_n564), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT112), .Z(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1072), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1063), .B1(new_n1088), .B2(new_n776), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1017), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n765), .B(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1089), .B1(new_n768), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n760), .A2(new_n1091), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n704), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n760), .A2(new_n1091), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(G393));
  XNOR2_X1  g0896(.A(new_n699), .B(new_n1008), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n768), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n964), .A2(new_n254), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n777), .B1(new_n213), .B2(new_n705), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n769), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n414), .B1(new_n800), .B2(G143), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n851), .B(new_n1102), .C1(new_n203), .C2(new_n805), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT114), .Z(new_n1104));
  OAI22_X1  g0904(.A1(new_n201), .A2(new_n819), .B1(new_n791), .B2(new_n265), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT115), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1105), .A2(new_n1106), .B1(new_n262), .B2(new_n803), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1106), .B2(new_n1105), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G150), .A2(new_n793), .B1(new_n807), .B2(G159), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT51), .Z(new_n1110));
  NAND3_X1  g0910(.A1(new_n1104), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n790), .A2(G294), .B1(G116), .B2(new_n983), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n585), .B2(new_n819), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT117), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G311), .A2(new_n807), .B1(new_n793), .B2(G317), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n414), .B1(new_n853), .B2(new_n1074), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n855), .B2(G283), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n823), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1111), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1101), .B1(new_n1121), .B2(new_n776), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n999), .A2(new_n832), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT113), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1098), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT118), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n760), .A2(new_n1091), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n704), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1097), .B1(new_n760), .B2(new_n1091), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1097), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1093), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1133), .A2(KEYINPUT118), .A3(new_n704), .A4(new_n1128), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1126), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G390));
  NAND4_X1  g0936(.A1(new_n956), .A2(G330), .A3(new_n839), .A4(new_n932), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n842), .A2(new_n935), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n932), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1140), .A2(new_n916), .B1(new_n915), .B2(new_n927), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n946), .A2(new_n926), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n916), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n720), .A2(new_n683), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n935), .B1(new_n1144), .B2(new_n840), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n932), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1138), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n927), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT39), .B1(new_n946), .B2(new_n926), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n1148), .A2(new_n1149), .B1(new_n936), .B2(new_n917), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n712), .A2(new_n715), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(new_n682), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n934), .B1(new_n1152), .B2(new_n839), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n916), .B(new_n1142), .C1(new_n1153), .C2(new_n933), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n1154), .A3(new_n1137), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(new_n767), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n769), .B1(new_n847), .B2(new_n357), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n774), .B1(new_n915), .B2(new_n927), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n207), .A2(new_n819), .B1(new_n791), .B2(new_n705), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G116), .B2(new_n807), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n793), .A2(G283), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n414), .B1(new_n853), .B2(new_n509), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1163), .B(new_n827), .C1(G77), .C2(new_n983), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n858), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n822), .A2(G50), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n855), .A2(new_n1067), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT53), .Z(new_n1168));
  NAND2_X1  g0968(.A1(new_n807), .A2(G132), .ZN(new_n1169));
  INV_X1    g0969(.A(G125), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n288), .B1(new_n803), .B2(new_n978), .C1(new_n1170), .C2(new_n853), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G128), .B2(new_n793), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .A4(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G137), .A2(new_n797), .B1(new_n790), .B2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT119), .Z(new_n1177));
  OAI21_X1  g0977(.A(new_n1165), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1158), .B(new_n1159), .C1(new_n776), .C2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1157), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n758), .A2(new_n442), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n884), .A2(new_n675), .A3(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(G330), .B(new_n839), .C1(new_n754), .C2(new_n755), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n933), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1137), .A2(new_n1184), .A3(new_n1153), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1183), .B(new_n932), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1139), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1156), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1147), .A2(new_n1182), .A3(new_n1155), .A4(new_n1188), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n704), .A3(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1180), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(G378));
  NAND3_X1  g0994(.A1(new_n441), .A2(new_n430), .A3(new_n887), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n430), .A2(new_n887), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n435), .A2(new_n437), .A3(new_n440), .A4(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n953), .B2(G330), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n757), .B(new_n1201), .C1(new_n949), .C2(new_n952), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n940), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1142), .A2(new_n956), .A3(new_n839), .A4(new_n932), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1206), .A2(KEYINPUT40), .B1(new_n950), .B2(new_n951), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1201), .B1(new_n1207), .B2(new_n757), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n940), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n953), .A2(G330), .A3(new_n1202), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1205), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1201), .A2(new_n773), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n769), .B1(new_n847), .B2(G50), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G50), .B1(new_n282), .B2(new_n290), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n207), .A2(new_n816), .B1(new_n791), .B2(new_n270), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G97), .B2(new_n797), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n822), .A2(G58), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G41), .B(new_n288), .C1(G283), .C2(new_n800), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n984), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1070), .B(new_n1220), .C1(G116), .C2(new_n793), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1217), .A2(new_n1218), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1215), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G33), .B(G41), .C1(new_n800), .C2(G124), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1170), .A2(new_n794), .B1(new_n791), .B2(new_n863), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n855), .A2(new_n1175), .B1(G150), .B2(new_n983), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n859), .B2(new_n819), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(G128), .C2(new_n807), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT59), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1225), .B1(new_n978), .B2(new_n813), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1229), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1224), .B1(new_n1223), .B2(new_n1222), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1214), .B1(new_n1234), .B2(new_n776), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1212), .A2(new_n768), .B1(new_n1213), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1188), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1182), .B1(new_n1156), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1212), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT57), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT120), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(KEYINPUT121), .A3(new_n1240), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1211), .A2(new_n1205), .B1(new_n1191), .B2(new_n1182), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT120), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(KEYINPUT57), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1241), .A2(new_n1242), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1238), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n704), .B1(new_n1247), .B2(KEYINPUT121), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1236), .B1(new_n1246), .B2(new_n1248), .ZN(G375));
  NOR2_X1   g1049(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n1021), .A3(new_n1189), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT122), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n981), .A2(new_n414), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT123), .Z(new_n1255));
  AOI22_X1  g1055(.A1(new_n983), .A2(new_n546), .B1(G303), .B2(new_n800), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1256), .B1(new_n206), .B2(new_n805), .C1(new_n791), .C2(new_n207), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G116), .A2(new_n797), .B1(new_n793), .B2(G294), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n809), .B2(new_n816), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1255), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n859), .A2(new_n794), .B1(new_n791), .B2(new_n864), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n983), .A2(G50), .B1(G128), .B2(new_n800), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n978), .B2(new_n805), .C1(new_n816), .C2(new_n863), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1261), .B(new_n1263), .C1(new_n797), .C2(new_n1175), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1218), .A2(new_n288), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n776), .B1(new_n1260), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n847), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1052), .B1(new_n1270), .B2(new_n203), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1269), .B(new_n1271), .C1(new_n774), .C2(new_n932), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1188), .B2(new_n768), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1253), .A2(new_n1274), .ZN(G381));
  AOI21_X1  g1075(.A(new_n1244), .B1(new_n1243), .B2(KEYINPUT57), .ZN(new_n1276));
  AND4_X1   g1076(.A1(new_n1244), .A2(new_n1212), .A3(KEYINPUT57), .A4(new_n1238), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n704), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT121), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1282), .A3(new_n1242), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n1193), .A3(new_n1236), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OR2_X1    g1085(.A1(G393), .A2(G396), .ZN(new_n1286));
  NOR4_X1   g1086(.A1(G381), .A2(G390), .A3(G384), .A4(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1050), .A3(new_n1287), .ZN(G407));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(G343), .C2(new_n1284), .ZN(G409));
  XNOR2_X1  g1089(.A(G393), .B(new_n834), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1126), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1291), .A2(new_n1048), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1048), .B2(new_n1135), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1292), .B1(new_n1135), .B2(new_n1048), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1290), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1290), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1135), .A2(new_n1048), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1298), .B(new_n1299), .C1(new_n1050), .C2(G390), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G375), .A2(G378), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1193), .B(new_n1236), .C1(new_n1020), .C2(new_n1239), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n681), .A2(G213), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1250), .B1(KEYINPUT60), .B2(new_n1189), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n884), .A2(new_n675), .A3(new_n1181), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1237), .A2(KEYINPUT60), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n704), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1274), .B1(new_n1308), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n872), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G384), .B(new_n1274), .C1(new_n1308), .C2(new_n1311), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1303), .A2(new_n1307), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1306), .B1(G375), .B2(G378), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1319), .A3(new_n1315), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n681), .A2(G213), .A3(G2897), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1313), .A2(new_n1314), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1193), .B1(new_n1283), .B2(new_n1236), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1325), .B1(new_n1326), .B2(new_n1306), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT126), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1302), .B1(new_n1321), .B2(new_n1329), .ZN(new_n1330));
  AND4_X1   g1130(.A1(KEYINPUT63), .A2(new_n1303), .A3(new_n1307), .A4(new_n1315), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT63), .B1(new_n1318), .B2(new_n1315), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1301), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT126), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1297), .A2(new_n1300), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1325), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1335), .B(new_n1328), .C1(new_n1318), .C2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1333), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1330), .A2(new_n1339), .ZN(G405));
  INV_X1    g1140(.A(new_n1315), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1341), .B1(new_n1285), .B2(new_n1326), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1303), .A2(new_n1284), .A3(new_n1315), .ZN(new_n1343));
  AOI22_X1  g1143(.A1(new_n1342), .A2(new_n1343), .B1(new_n1302), .B2(KEYINPUT127), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1301), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1342), .A2(new_n1345), .A3(new_n1301), .A4(new_n1343), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(G402));
endmodule


