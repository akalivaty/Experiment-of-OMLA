//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n450, new_n451, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n570, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n622, new_n624, new_n625, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137, new_n1138;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  INV_X1    g024(.A(G567), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT69), .Z(G217));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n456), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT70), .Z(new_n462));
  OAI21_X1  g037(.A(new_n462), .B1(new_n450), .B2(new_n457), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT71), .Z(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT72), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT74), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT73), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT73), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n465), .A2(G2104), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n480), .A2(G137), .B1(G101), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n471), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n479), .A2(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n480), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OR2_X1    g066(.A1(new_n465), .A2(G114), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n473), .A2(new_n472), .B1(new_n475), .B2(KEYINPUT3), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT3), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT75), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n497), .A2(new_n498), .A3(G126), .A4(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n477), .A2(G126), .A3(G2105), .A4(new_n478), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT75), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n494), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT76), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI211_X1 g079(.A(KEYINPUT76), .B(new_n494), .C1(new_n499), .C2(new_n501), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n477), .A2(G138), .A3(new_n465), .A4(new_n478), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT4), .A2(G2105), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n510));
  OAI211_X1 g085(.A(G138), .B(new_n508), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT77), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n466), .A2(new_n513), .A3(G138), .A4(new_n508), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NOR3_X1   g092(.A1(new_n504), .A2(new_n505), .A3(new_n517), .ZN(G164));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT79), .B1(new_n519), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT79), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT5), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(new_n523), .B1(new_n519), .B2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G62), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT80), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n524), .A2(KEYINPUT80), .A3(G62), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT6), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(G651), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(KEYINPUT78), .A3(KEYINPUT6), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n534), .A2(new_n536), .B1(new_n533), .B2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n524), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(G88), .A2(new_n539), .B1(new_n541), .B2(G50), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n531), .A2(new_n542), .ZN(G303));
  INV_X1    g118(.A(G303), .ZN(G166));
  AOI22_X1  g119(.A1(G89), .A2(new_n539), .B1(new_n541), .B2(G51), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT81), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT7), .Z(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(G168));
  AOI22_X1  g128(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n535), .ZN(new_n555));
  INV_X1    g130(.A(G90), .ZN(new_n556));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n538), .A2(new_n556), .B1(new_n540), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(G171));
  AOI22_X1  g134(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(G651), .A3(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(G81), .A2(new_n539), .B1(new_n541), .B2(G43), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT83), .Z(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  XOR2_X1   g144(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n570));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G188));
  NAND2_X1  g148(.A1(new_n541), .A2(G53), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT85), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n574), .B(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n524), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT86), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n583), .A2(KEYINPUT87), .A3(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n539), .A2(G91), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n581), .A2(new_n584), .A3(new_n585), .A4(new_n588), .ZN(G299));
  XNOR2_X1  g164(.A(G171), .B(KEYINPUT88), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G301));
  INV_X1    g166(.A(G168), .ZN(G286));
  NAND2_X1  g167(.A1(new_n539), .A2(G87), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n541), .A2(G49), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G288));
  AOI22_X1  g171(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n535), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  INV_X1    g174(.A(G48), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n538), .A2(new_n599), .B1(new_n540), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(G85), .A2(new_n539), .B1(new_n541), .B2(G47), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n535), .B2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n539), .A2(G92), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT10), .Z(new_n609));
  NAND2_X1  g184(.A1(new_n541), .A2(G54), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n524), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(new_n535), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(G868), .B2(new_n614), .ZN(G284));
  OAI21_X1  g190(.A(new_n607), .B1(G868), .B2(new_n614), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  XOR2_X1   g192(.A(G299), .B(KEYINPUT89), .Z(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  XOR2_X1   g194(.A(G280), .B(KEYINPUT90), .Z(G297));
  NOR2_X1   g195(.A1(new_n613), .A2(G559), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G860), .B2(new_n614), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT91), .Z(G148));
  INV_X1    g198(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT92), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n466), .A2(new_n481), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n485), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n480), .A2(G135), .ZN(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n635), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n632), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2435), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n645), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n657), .B2(new_n660), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n669), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  AOI22_X1  g250(.A1(new_n673), .A2(KEYINPUT20), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n669), .A3(new_n672), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n678), .C1(KEYINPUT20), .C2(new_n673), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  NAND2_X1  g260(.A1(new_n485), .A2(G119), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n480), .A2(G131), .ZN(new_n687));
  NOR2_X1   g262(.A1(G95), .A2(G2105), .ZN(new_n688));
  OAI21_X1  g263(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n686), .B(new_n687), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(G25), .B(new_n690), .S(G29), .Z(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT35), .B(G1991), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT95), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT94), .B(KEYINPUT96), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G24), .B(G290), .S(G16), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1986), .ZN(new_n700));
  INV_X1    g275(.A(new_n697), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n695), .B2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G23), .B(G288), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT33), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1976), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G1971), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(G1971), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(G6), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n602), .B2(new_n706), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n705), .A2(new_n709), .A3(new_n710), .A4(new_n714), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n698), .B(new_n702), .C1(new_n715), .C2(KEYINPUT34), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n716), .B1(KEYINPUT34), .B2(new_n715), .C1(G1986), .C2(new_n699), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT36), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n706), .A2(G21), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G168), .B2(new_n706), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT100), .B(G1966), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT99), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G299), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT23), .B1(new_n724), .B2(new_n706), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n706), .A2(G20), .ZN(new_n726));
  MUX2_X1   g301(.A(KEYINPUT23), .B(new_n725), .S(new_n726), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1956), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n480), .A2(G141), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n485), .A2(G129), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT26), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G105), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n729), .A2(new_n730), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G32), .B(new_n734), .S(G29), .Z(new_n735));
  XOR2_X1   g310(.A(KEYINPUT27), .B(G1996), .Z(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G34), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT98), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(G34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n483), .B2(new_n737), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n735), .A2(new_n736), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G5), .A2(G16), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G171), .B2(G16), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(G1961), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT102), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n706), .A2(G4), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n614), .B2(new_n706), .ZN(new_n753));
  INV_X1    g328(.A(G1348), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n706), .A2(G19), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n565), .B2(new_n706), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G1341), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n737), .A2(G26), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n485), .A2(G128), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n480), .A2(G140), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n759), .B1(new_n765), .B2(new_n737), .ZN(new_n766));
  MUX2_X1   g341(.A(new_n759), .B(new_n766), .S(KEYINPUT28), .Z(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n755), .A2(new_n758), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n751), .B1(new_n771), .B2(KEYINPUT97), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n735), .A2(new_n736), .B1(new_n745), .B2(new_n746), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n481), .A2(G103), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT25), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n480), .A2(G139), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n466), .A2(G127), .ZN(new_n777));
  AND2_X1   g352(.A1(G115), .A2(G2104), .ZN(new_n778));
  OAI21_X1  g353(.A(G2105), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(G2072), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G11), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(G2072), .ZN(new_n784));
  INV_X1    g359(.A(G28), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n785), .A2(KEYINPUT101), .A3(KEYINPUT30), .ZN(new_n786));
  OAI21_X1  g361(.A(KEYINPUT101), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(new_n737), .ZN(new_n788));
  AOI211_X1 g363(.A(new_n786), .B(new_n788), .C1(KEYINPUT30), .C2(new_n785), .ZN(new_n789));
  INV_X1    g364(.A(new_n637), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G29), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n791), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n773), .B(new_n792), .C1(G1961), .C2(new_n749), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n737), .A2(G35), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G162), .B2(new_n737), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT29), .B(G2090), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G164), .A2(new_n737), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G27), .B2(new_n737), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n793), .A2(new_n797), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n770), .A2(new_n804), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n728), .A2(new_n772), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n718), .A2(new_n723), .A3(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  INV_X1    g383(.A(G93), .ZN(new_n809));
  INV_X1    g384(.A(G55), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n538), .A2(new_n809), .B1(new_n540), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT103), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n813), .A2(new_n814), .B1(new_n535), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n614), .A2(G559), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n565), .B1(KEYINPUT104), .B2(new_n816), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(KEYINPUT104), .B2(new_n816), .ZN(new_n823));
  INV_X1    g398(.A(new_n816), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n825), .A3(new_n565), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n821), .B(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n818), .B1(new_n828), .B2(G860), .ZN(G145));
  XNOR2_X1  g404(.A(new_n483), .B(KEYINPUT105), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n490), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n690), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n765), .B(new_n734), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n499), .A2(new_n501), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(new_n516), .A3(new_n493), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n630), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n832), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n637), .B(new_n780), .Z(new_n839));
  AND2_X1   g414(.A1(new_n480), .A2(G142), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT106), .ZN(new_n841));
  OR2_X1    g416(.A1(G106), .A2(G2105), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n480), .A2(KEYINPUT106), .A3(G142), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n485), .A2(G130), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n841), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n839), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n838), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g426(.A1(G299), .A2(new_n614), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n588), .A2(new_n585), .A3(new_n584), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n853), .A2(new_n581), .A3(new_n613), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT107), .B1(new_n852), .B2(new_n854), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n724), .B2(new_n613), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(KEYINPUT41), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n827), .B(new_n621), .ZN(new_n863));
  MUX2_X1   g438(.A(new_n855), .B(new_n862), .S(new_n863), .Z(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n866), .ZN(new_n868));
  XNOR2_X1  g443(.A(G303), .B(G290), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G288), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n602), .B(KEYINPUT109), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT108), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n870), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n867), .A2(new_n868), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n867), .B2(new_n868), .ZN(new_n876));
  OAI21_X1  g451(.A(G868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(G868), .B2(new_n824), .ZN(G295));
  OAI21_X1  g453(.A(new_n877), .B1(G868), .B2(new_n824), .ZN(G331));
  NAND2_X1  g454(.A1(G301), .A2(G168), .ZN(new_n880));
  NAND2_X1  g455(.A1(G286), .A2(G171), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n827), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n826), .A3(new_n823), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n855), .B1(new_n886), .B2(new_n856), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n885), .B(KEYINPUT41), .C1(new_n857), .C2(new_n859), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n874), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n855), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n860), .A2(new_n861), .A3(new_n885), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n874), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT112), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n887), .A2(KEYINPUT112), .A3(new_n874), .A4(new_n888), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n849), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT43), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT113), .ZN(new_n898));
  INV_X1    g473(.A(new_n892), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n890), .A2(new_n891), .A3(new_n874), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n899), .A2(new_n849), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT113), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n896), .A2(new_n904), .A3(KEYINPUT43), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n898), .A2(KEYINPUT44), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT111), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n901), .B2(new_n902), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n894), .A2(new_n902), .A3(new_n849), .A4(new_n895), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n899), .A2(new_n849), .A3(new_n900), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n906), .A2(new_n914), .ZN(G397));
  NAND3_X1  g490(.A1(new_n471), .A2(G40), .A3(new_n482), .ZN(new_n916));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n835), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT116), .B1(new_n918), .B2(KEYINPUT50), .ZN(new_n919));
  AOI21_X1  g494(.A(G1384), .B1(new_n502), .B2(new_n516), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT116), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT50), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n916), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n925));
  AOI21_X1  g500(.A(G1348), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT121), .ZN(new_n927));
  INV_X1    g502(.A(new_n916), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n920), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(G2067), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(new_n932));
  AND4_X1   g507(.A1(new_n921), .A2(new_n835), .A3(new_n922), .A4(new_n917), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n500), .A2(KEYINPUT75), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n500), .A2(KEYINPUT75), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n493), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT76), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n502), .A2(new_n503), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n516), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n922), .B1(new_n940), .B2(new_n917), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n754), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n930), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT121), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT60), .B1(new_n931), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(KEYINPUT123), .A3(new_n613), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n927), .B1(new_n926), .B2(new_n930), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(KEYINPUT121), .A3(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n613), .A2(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n613), .A2(KEYINPUT123), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n949), .A2(KEYINPUT60), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n946), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(G164), .B2(G1384), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n918), .A2(new_n955), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n928), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(G1996), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n918), .A2(new_n916), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT58), .B(G1341), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n565), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT59), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT56), .B(G2072), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n956), .A2(new_n928), .A3(new_n958), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT120), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n918), .A2(KEYINPUT50), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n940), .A2(new_n917), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n928), .B(new_n969), .C1(new_n970), .C2(KEYINPUT50), .ZN(new_n971));
  INV_X1    g546(.A(G1956), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n916), .B1(new_n970), .B2(new_n955), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n958), .A4(new_n966), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n578), .A2(KEYINPUT57), .ZN(new_n978));
  AOI22_X1  g553(.A1(G299), .A2(KEYINPUT57), .B1(new_n853), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n979), .A2(new_n968), .A3(new_n973), .A4(new_n976), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT61), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT122), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n977), .B2(new_n980), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n981), .A2(new_n985), .A3(KEYINPUT61), .A4(new_n982), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n954), .A2(new_n965), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n982), .A2(new_n614), .A3(new_n948), .A4(new_n947), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n990), .A2(new_n981), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n940), .A2(KEYINPUT45), .A3(new_n917), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n920), .A2(KEYINPUT45), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n928), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n721), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n924), .A2(new_n925), .A3(new_n746), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT124), .B(G8), .C1(new_n1000), .C2(G286), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n998), .B2(new_n999), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G168), .A2(new_n1004), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT124), .B(KEYINPUT51), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G303), .A2(G8), .ZN(new_n1011));
  XOR2_X1   g586(.A(new_n1011), .B(KEYINPUT55), .Z(new_n1012));
  AOI21_X1  g587(.A(G1971), .B1(new_n974), .B2(new_n958), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n934), .A2(G2090), .A3(new_n941), .ZN(new_n1014));
  OAI211_X1 g589(.A(G8), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1981), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n602), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(G1981), .B1(new_n598), .B2(new_n601), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT117), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1017), .A2(new_n1021), .A3(KEYINPUT49), .A4(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n961), .A2(new_n1004), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n929), .B(G8), .C1(new_n1029), .C2(G288), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT52), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1027), .B(new_n1032), .C1(new_n1029), .C2(G288), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n959), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n504), .A2(new_n505), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n1038), .B2(new_n516), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n916), .B1(new_n1039), .B2(new_n922), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n969), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1004), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1015), .B(new_n1035), .C1(new_n1043), .C2(new_n1012), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n956), .A2(new_n800), .A3(new_n928), .A4(new_n958), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G2078), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n993), .A2(new_n928), .A3(new_n995), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n934), .B2(new_n941), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1047), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G40), .ZN(new_n1054));
  NOR4_X1   g629(.A1(new_n469), .A2(new_n1048), .A3(new_n1054), .A4(G2078), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n958), .A2(new_n995), .A3(new_n482), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT45), .B1(new_n940), .B2(new_n917), .ZN(new_n1057));
  NOR4_X1   g632(.A1(new_n1057), .A2(G2078), .A3(new_n916), .A4(new_n957), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1046), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1052), .B(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1053), .A2(G301), .B1(G171), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1044), .B1(new_n1061), .B2(KEYINPUT54), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1053), .A2(G301), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1060), .A2(new_n590), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1010), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n992), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT126), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT63), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1005), .A2(G168), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1044), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n924), .A2(new_n925), .A3(new_n1041), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1057), .A2(new_n916), .A3(new_n957), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(G1971), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1012), .B1(new_n1077), .B2(G8), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1074), .B1(new_n1078), .B2(new_n1034), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1004), .B1(new_n1037), .B2(new_n1075), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1035), .B(KEYINPUT119), .C1(new_n1080), .C2(new_n1012), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1079), .A2(KEYINPUT63), .A3(new_n1081), .A4(new_n1015), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1073), .B1(new_n1082), .B2(new_n1072), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1015), .A2(new_n1034), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1028), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G288), .A2(G1976), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT118), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1017), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1027), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1083), .A2(new_n1085), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1069), .A2(new_n1070), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1067), .B1(new_n989), .B2(new_n991), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1083), .A2(new_n1085), .A3(new_n1090), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT126), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1010), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1044), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(new_n1064), .C1(new_n1097), .C2(new_n1096), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1092), .A2(new_n1095), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n994), .A2(new_n928), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT114), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n734), .ZN(new_n1103));
  INV_X1    g678(.A(G1996), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT115), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1101), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1104), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1108), .A2(new_n734), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n764), .B(G2067), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1102), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1106), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n690), .B(new_n694), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1102), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G290), .B(G1986), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1107), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1100), .A2(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1101), .A2(G1986), .A3(G290), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT48), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n690), .A2(new_n693), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1112), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n765), .A2(new_n768), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1114), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT46), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1108), .B(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1129), .A2(new_n1103), .A3(new_n1111), .A4(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT47), .Z(new_n1132));
  NOR3_X1   g707(.A1(new_n1121), .A2(new_n1125), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1118), .A2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g709(.A(G319), .ZN(new_n1136));
  NOR2_X1   g710(.A1(new_n1136), .A2(G229), .ZN(new_n1137));
  AOI211_X1 g711(.A(G401), .B(G227), .C1(new_n848), .C2(new_n849), .ZN(new_n1138));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n1137), .A3(new_n1138), .ZN(G225));
  INV_X1    g713(.A(G225), .ZN(G308));
endmodule


