//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n564, new_n566, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n457), .B1(new_n448), .B2(new_n454), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT3), .B1(new_n460), .B2(KEYINPUT70), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n461), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT72), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n468), .B1(new_n460), .B2(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n465), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n471), .B2(G101), .ZN(new_n472));
  INV_X1    g047(.A(G101), .ZN(new_n473));
  AOI211_X1 g048(.A(KEYINPUT72), .B(new_n473), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n466), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n463), .A2(new_n460), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n481), .B(G125), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n488));
  OAI21_X1  g063(.A(G125), .B1(new_n483), .B2(new_n484), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT68), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n485), .A3(new_n476), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n475), .B1(new_n488), .B2(new_n493), .ZN(G160));
  NAND3_X1  g069(.A1(new_n461), .A2(new_n464), .A3(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G124), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n465), .A2(G112), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n495), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n500));
  XOR2_X1   g075(.A(new_n500), .B(KEYINPUT73), .Z(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n501), .B2(G136), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT74), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G162));
  NOR2_X1   g079(.A1(new_n483), .A2(new_n484), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n505), .A2(new_n506), .A3(G2105), .ZN(new_n507));
  XOR2_X1   g082(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n508));
  NAND4_X1  g083(.A1(new_n461), .A2(new_n464), .A3(G138), .A4(new_n465), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(new_n508), .B1(KEYINPUT4), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G126), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n465), .A2(G114), .ZN(new_n512));
  OAI21_X1  g087(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n495), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n510), .A2(new_n514), .ZN(G164));
  XOR2_X1   g090(.A(KEYINPUT6), .B(G651), .Z(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR3_X1   g096(.A1(new_n516), .A2(new_n521), .A3(KEYINPUT76), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n518), .A2(new_n520), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(G75), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G62), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(G50), .A2(G543), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n531), .A2(G651), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n528), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n527), .A2(G89), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n516), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n525), .A2(KEYINPUT77), .ZN(new_n539));
  NOR3_X1   g114(.A1(new_n538), .A2(new_n517), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n524), .A2(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n536), .A2(new_n541), .A3(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  NAND2_X1  g123(.A1(new_n527), .A2(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n540), .A2(G52), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G651), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(new_n527), .A2(G81), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT78), .B(G43), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n540), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n552), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT79), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G188));
  NAND3_X1  g144(.A1(new_n540), .A2(KEYINPUT80), .A3(G53), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n527), .A2(KEYINPUT81), .A3(G91), .ZN(new_n572));
  AOI21_X1  g147(.A(KEYINPUT81), .B1(new_n527), .B2(G91), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n521), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n573), .B1(G651), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n527), .A2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n540), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n527), .A2(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n521), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(G48), .A2(G543), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n586), .A2(G651), .B1(new_n525), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n527), .A2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n540), .A2(G47), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n590), .B(new_n591), .C1(new_n552), .C2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n527), .A2(G92), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT10), .Z(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n521), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n540), .A2(G54), .B1(G651), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n594), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  XNOR2_X1  g182(.A(KEYINPUT82), .B(G559), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(G860), .B2(new_n609), .ZN(G148));
  NAND2_X1  g185(.A1(new_n601), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g189(.A(new_n505), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n471), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2100), .Z(new_n619));
  INV_X1    g194(.A(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n465), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI22_X1  g197(.A1(new_n495), .A2(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n501), .B2(G135), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT83), .B(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n626), .ZN(G156));
  XOR2_X1   g202(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n628));
  XOR2_X1   g203(.A(KEYINPUT15), .B(G2435), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n630), .B2(new_n631), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT16), .B(G1341), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(G14), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n633), .B2(new_n639), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT85), .Z(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XOR2_X1   g218(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n643), .B2(new_n646), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(KEYINPUT87), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(KEYINPUT87), .B2(new_n650), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT89), .Z(new_n653));
  AND3_X1   g228(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n643), .A2(new_n646), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(new_n648), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT86), .Z(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n653), .B(new_n658), .C1(KEYINPUT18), .C2(new_n657), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT91), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(KEYINPUT91), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT20), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n667), .A2(new_n668), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(new_n671), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n671), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n669), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n676), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT92), .ZN(new_n684));
  INV_X1    g259(.A(G1991), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n683), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(G1991), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n664), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(G1991), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n684), .A2(new_n685), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n694), .A3(G1996), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n692), .B1(new_n690), .B2(new_n695), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n663), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n690), .A2(new_n695), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(new_n691), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n701), .A2(new_n662), .A3(new_n696), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(G229));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G35), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT29), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G2090), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT101), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n501), .A2(G141), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT97), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT26), .ZN(new_n715));
  INV_X1    g290(.A(G129), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n495), .A2(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n715), .B(new_n717), .C1(G105), .C2(new_n471), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT98), .ZN(new_n720));
  MUX2_X1   g295(.A(G32), .B(new_n720), .S(G29), .Z(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT99), .Z(new_n724));
  NOR2_X1   g299(.A1(new_n710), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G27), .A2(G29), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G164), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2078), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n601), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G4), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G1348), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT94), .B(G16), .ZN(new_n733));
  MUX2_X1   g308(.A(G19), .B(new_n561), .S(new_n733), .Z(new_n734));
  INV_X1    g309(.A(G1341), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n732), .B(new_n736), .C1(new_n731), .C2(new_n730), .ZN(new_n737));
  INV_X1    g312(.A(G20), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT23), .Z(new_n740));
  INV_X1    g315(.A(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n605), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n501), .A2(G139), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT25), .Z(new_n746));
  AOI22_X1  g321(.A1(new_n615), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n746), .C1(new_n465), .C2(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G33), .B(new_n748), .S(G29), .Z(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G2072), .Z(new_n750));
  NAND2_X1  g325(.A1(G171), .A2(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G5), .B2(G16), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT24), .ZN(new_n755));
  INV_X1    g330(.A(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n755), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G160), .B2(new_n704), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n750), .B(new_n754), .C1(G2084), .C2(new_n759), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n737), .A2(new_n743), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n704), .A2(G26), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n501), .A2(G140), .ZN(new_n763));
  INV_X1    g338(.A(G128), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n465), .A2(G116), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n766));
  OAI22_X1  g341(.A1(new_n495), .A2(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(new_n704), .ZN(new_n769));
  MUX2_X1   g344(.A(new_n762), .B(new_n769), .S(KEYINPUT28), .Z(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT96), .B(G2067), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n770), .A2(new_n771), .B1(new_n759), .B2(G2084), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n708), .B2(G2090), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n741), .A2(G21), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G168), .B2(new_n741), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G1966), .Z(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G28), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n704), .B1(new_n778), .B2(G28), .ZN(new_n780));
  AND2_X1   g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  NOR2_X1   g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n624), .B2(G29), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n777), .B(new_n784), .C1(new_n753), .C2(new_n752), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT100), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n722), .B2(new_n721), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n725), .A2(new_n761), .A3(new_n774), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(G288), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT33), .B(G1976), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G22), .B(G303), .S(new_n733), .Z(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G6), .B(G305), .S(G16), .Z(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n793), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT34), .Z(new_n801));
  AND2_X1   g376(.A1(new_n704), .A2(G25), .ZN(new_n802));
  OR2_X1    g377(.A1(G95), .A2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n803), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n804));
  INV_X1    g379(.A(G119), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n495), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n501), .B2(G131), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT93), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT93), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n802), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT35), .B(G1991), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G24), .B(G290), .S(new_n733), .Z(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT95), .B(G1986), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n811), .A2(new_n813), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n801), .A2(new_n814), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT36), .Z(new_n820));
  NOR2_X1   g395(.A1(new_n788), .A2(new_n820), .ZN(G311));
  INV_X1    g396(.A(G311), .ZN(G150));
  NAND2_X1  g397(.A1(new_n527), .A2(G93), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n540), .A2(G55), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n823), .B(new_n824), .C1(new_n552), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n601), .A2(G559), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT39), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT102), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT38), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n562), .B(new_n826), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G860), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n832), .B2(new_n833), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n828), .B1(new_n834), .B2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n503), .B(G160), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n624), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n501), .A2(G142), .ZN(new_n840));
  INV_X1    g415(.A(G130), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n465), .A2(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  OAI221_X1 g418(.A(new_n840), .B1(new_n841), .B2(new_n495), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n810), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT103), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n617), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n845), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n617), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n851), .A3(KEYINPUT104), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n719), .A2(new_n748), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n720), .B2(new_n748), .ZN(new_n855));
  INV_X1    g430(.A(G164), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n768), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT104), .B1(new_n847), .B2(new_n851), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n853), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n858), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n849), .A2(new_n850), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n846), .A2(new_n617), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n861), .B1(new_n865), .B2(new_n852), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n839), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n858), .B1(new_n853), .B2(new_n859), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n863), .A2(new_n864), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n839), .B1(new_n869), .B2(new_n861), .ZN(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g448(.A1(new_n596), .A2(new_n600), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n605), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n874), .B(G299), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT41), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n611), .B(new_n833), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT105), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n878), .ZN(new_n883));
  MUX2_X1   g458(.A(new_n882), .B(KEYINPUT105), .S(new_n883), .Z(new_n884));
  XOR2_X1   g459(.A(G290), .B(KEYINPUT106), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G305), .ZN(new_n886));
  XNOR2_X1  g461(.A(G288), .B(G303), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n884), .B(new_n891), .ZN(new_n892));
  MUX2_X1   g467(.A(new_n826), .B(new_n892), .S(G868), .Z(G295));
  MUX2_X1   g468(.A(new_n826), .B(new_n892), .S(G868), .Z(G331));
  XOR2_X1   g469(.A(G286), .B(G301), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n833), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n880), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n890), .B(new_n897), .C1(new_n878), .C2(new_n896), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  INV_X1    g474(.A(new_n896), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n879), .B2(new_n877), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n896), .A2(new_n878), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n901), .A2(new_n902), .B1(new_n888), .B2(new_n889), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT107), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n898), .A2(new_n899), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n908), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n907), .A2(new_n909), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n904), .A2(new_n913), .A3(KEYINPUT43), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n906), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n904), .A2(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n907), .A2(new_n909), .A3(new_n911), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n910), .ZN(new_n918));
  MUX2_X1   g493(.A(new_n915), .B(new_n918), .S(KEYINPUT44), .Z(G397));
  NOR2_X1   g494(.A1(new_n720), .A2(G1996), .ZN(new_n920));
  INV_X1    g495(.A(G2067), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n768), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n763), .A2(G2067), .A3(new_n767), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n719), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n664), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n810), .A2(new_n812), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n808), .A2(new_n809), .A3(new_n813), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n920), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(G290), .B(G1986), .Z(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(KEYINPUT109), .B(G1384), .Z(new_n933));
  NAND2_X1  g508(.A1(new_n856), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(G40), .B(new_n466), .C1(new_n472), .C2(new_n474), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n489), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n940));
  AOI211_X1 g515(.A(KEYINPUT69), .B(new_n465), .C1(new_n940), .C2(new_n485), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n492), .B1(new_n491), .B2(G2105), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT110), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n939), .B(new_n945), .C1(new_n941), .C2(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n937), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n932), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT54), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n510), .B2(new_n514), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n953), .A2(new_n954), .A3(new_n935), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n953), .B2(new_n935), .ZN(new_n956));
  OAI211_X1 g531(.A(KEYINPUT45), .B(new_n933), .C1(new_n510), .C2(new_n514), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G2078), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n947), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT53), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n944), .B2(new_n946), .ZN(new_n965));
  INV_X1    g540(.A(new_n953), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n961), .A2(new_n962), .B1(new_n969), .B2(new_n753), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n953), .B(new_n935), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n946), .B2(new_n944), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(KEYINPUT53), .A3(new_n960), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(G301), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT125), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n938), .B1(G2105), .B2(new_n491), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n978), .A2(KEYINPUT123), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(KEYINPUT123), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n936), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT124), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n958), .A2(new_n962), .A3(G2078), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G301), .B1(new_n986), .B2(new_n970), .ZN(new_n987));
  OR4_X1    g562(.A1(new_n951), .A2(new_n976), .A3(new_n977), .A4(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1981), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n583), .A2(new_n989), .A3(new_n588), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(G305), .B2(G1981), .ZN(new_n995));
  AOI211_X1 g570(.A(KEYINPUT116), .B(new_n989), .C1(new_n583), .C2(new_n588), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n992), .A2(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT49), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n947), .A2(new_n966), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(KEYINPUT114), .A3(G8), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n953), .B1(new_n944), .B2(new_n946), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT117), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n959), .A2(new_n947), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n795), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G2090), .B2(new_n969), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT113), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(KEYINPUT113), .B2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1011), .A2(G8), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1000), .A2(new_n1004), .B1(G1976), .B2(new_n790), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n1021), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1007), .A2(new_n1020), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n970), .A2(new_n973), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G171), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n986), .A2(G301), .A3(new_n970), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT54), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n488), .A2(new_n493), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n945), .B1(new_n1035), .B2(new_n939), .ZN(new_n1036));
  AOI211_X1 g611(.A(KEYINPUT110), .B(new_n938), .C1(new_n488), .C2(new_n493), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1034), .B(new_n963), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n968), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n965), .A2(new_n1034), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1039), .A2(new_n1040), .A3(G2090), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1009), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1018), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g620(.A1(new_n969), .A2(G2084), .B1(new_n972), .B2(G1966), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G286), .A2(G8), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(KEYINPUT51), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(G8), .A3(G286), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(G8), .C1(new_n1046), .C2(G286), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n988), .A2(new_n1029), .A3(new_n1045), .A4(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G299), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n571), .A2(new_n572), .A3(new_n577), .A4(new_n1055), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n968), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n965), .B2(new_n1034), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n963), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT118), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1956), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT56), .B(G2072), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n959), .A2(new_n947), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1059), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1059), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1066), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1072), .A3(KEYINPUT61), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1068), .A2(new_n1072), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT61), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(new_n735), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1008), .A2(G1996), .B1(new_n1002), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n562), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1083), .A2(KEYINPUT59), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(KEYINPUT59), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1078), .A2(new_n1079), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1077), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT122), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1077), .A2(new_n1089), .A3(new_n1086), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n969), .A2(new_n731), .B1(new_n921), .B2(new_n1002), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(KEYINPUT60), .B2(new_n601), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1088), .A2(new_n1090), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1068), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1091), .A2(new_n874), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1072), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1054), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1006), .B(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1101), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n790), .A2(new_n1022), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1101), .A2(new_n1103), .B1(new_n992), .B2(new_n993), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1005), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1047), .A2(G286), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1011), .A2(G8), .A3(new_n1019), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n1018), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT63), .B1(new_n1108), .B2(new_n1028), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1031), .B1(new_n1053), .B2(KEYINPUT62), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT63), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1110), .A2(new_n1111), .B1(new_n1112), .B2(new_n1106), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1044), .A2(new_n1043), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1029), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1105), .B(new_n1109), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n950), .B1(new_n1099), .B2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n948), .A2(G1986), .A3(G290), .ZN(new_n1118));
  XOR2_X1   g693(.A(new_n1118), .B(KEYINPUT48), .Z(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n930), .B2(new_n948), .ZN(new_n1120));
  NOR2_X1   g695(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n925), .B(new_n924), .C1(G1996), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n949), .ZN(new_n1123));
  AND2_X1   g698(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n948), .A2(G1996), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT47), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n920), .A2(new_n926), .A3(new_n928), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n949), .B1(new_n1128), .B2(new_n923), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1120), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1117), .A2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g706(.A1(G227), .A2(new_n458), .A3(new_n641), .ZN(new_n1133));
  NAND3_X1  g707(.A1(new_n699), .A2(new_n702), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n1135));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g710(.A1(new_n699), .A2(new_n702), .A3(KEYINPUT127), .A4(new_n1133), .ZN(new_n1137));
  NAND4_X1  g711(.A1(new_n1136), .A2(new_n915), .A3(new_n872), .A4(new_n1137), .ZN(G225));
  INV_X1    g712(.A(G225), .ZN(G308));
endmodule


