//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n205), .A2(KEYINPUT28), .B1(new_n206), .B2(new_n204), .ZN(new_n207));
  INV_X1    g006(.A(G169gat), .ZN(new_n208));
  INV_X1    g007(.A(G176gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT67), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n208), .A2(new_n209), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n206), .A2(KEYINPUT27), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT27), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G183gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(new_n204), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n207), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT23), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n216), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT25), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n206), .A2(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n204), .A2(G183gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT69), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n242));
  XNOR2_X1  g041(.A(G183gat), .B(G190gat), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n242), .B(new_n239), .C1(new_n243), .C2(new_n235), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n234), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n233), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n238), .A2(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT23), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n215), .B1(new_n248), .B2(new_n218), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT66), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n218), .A2(new_n251), .A3(new_n248), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n247), .B(new_n249), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n227), .B1(new_n246), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT73), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT73), .ZN(new_n259));
  INV_X1    g058(.A(new_n257), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n233), .A2(new_n245), .B1(new_n253), .B2(new_n254), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n259), .B(new_n260), .C1(new_n261), .C2(new_n227), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT29), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n261), .B2(new_n227), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n257), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G211gat), .ZN(new_n268));
  INV_X1    g067(.A(G218gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G211gat), .A2(G218gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT72), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n270), .A2(new_n274), .A3(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(G197gat), .A2(G204gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(G197gat), .A2(G204gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT22), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n271), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(new_n280), .A3(new_n275), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n267), .A2(KEYINPUT74), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n258), .A2(new_n262), .B1(new_n257), .B2(new_n265), .ZN(new_n287));
  INV_X1    g086(.A(new_n284), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n256), .A2(new_n257), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n257), .B2(new_n265), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n288), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n285), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n294));
  XOR2_X1   g093(.A(G8gat), .B(G36gat), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT75), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  AND3_X1   g097(.A1(new_n293), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n294), .B1(new_n293), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT2), .ZN(new_n303));
  AND2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G141gat), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT78), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n316), .A3(new_n310), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n315), .A2(new_n317), .A3(new_n303), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT77), .B1(new_n304), .B2(new_n305), .ZN(new_n319));
  INV_X1    g118(.A(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(new_n302), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n312), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G113gat), .ZN(new_n328));
  INV_X1    g127(.A(G113gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332));
  INV_X1    g131(.A(G134gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G127gat), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G134gat), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n331), .A2(new_n332), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n336), .ZN(new_n338));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(KEYINPUT1), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT82), .B1(new_n326), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n306), .A2(new_n311), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n319), .A2(new_n324), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n315), .A2(new_n317), .A3(new_n303), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n337), .A2(new_n340), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n326), .A2(KEYINPUT3), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n346), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n358), .A3(new_n341), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n353), .A2(new_n354), .A3(new_n355), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n355), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n362), .B(new_n351), .C1(new_n346), .C2(new_n348), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n345), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n364), .A3(new_n312), .ZN(new_n365));
  INV_X1    g164(.A(new_n351), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT81), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  INV_X1    g168(.A(new_n349), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n361), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n326), .A2(new_n341), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n342), .A2(new_n349), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n355), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n360), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(G57gat), .B(G85gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT6), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n360), .B(new_n383), .C1(new_n373), .C2(new_n378), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n379), .A2(KEYINPUT6), .A3(new_n384), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n298), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n285), .A2(new_n289), .A3(new_n292), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n298), .A2(new_n393), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n285), .A2(new_n289), .A3(new_n292), .A4(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n390), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n301), .B2(new_n397), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n390), .A2(new_n394), .A3(new_n396), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n293), .A2(new_n298), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT76), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n293), .A2(new_n294), .A3(new_n298), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n256), .A2(new_n348), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n341), .B1(new_n261), .B2(new_n227), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n409), .B(KEYINPUT64), .Z(new_n410));
  OAI21_X1  g209(.A(KEYINPUT34), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT34), .ZN(new_n412));
  INV_X1    g211(.A(new_n410), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n406), .A2(new_n407), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G15gat), .B(G43gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(new_n410), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT33), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT33), .B1(new_n408), .B2(new_n410), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n411), .B(new_n414), .C1(new_n423), .C2(new_n418), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(KEYINPUT32), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n422), .A2(KEYINPUT32), .A3(new_n419), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n358), .A2(new_n264), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n284), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n282), .A2(new_n264), .A3(new_n283), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n432), .A2(new_n357), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n433), .B2(new_n346), .ZN(new_n434));
  INV_X1    g233(.A(G228gat), .ZN(new_n435));
  INV_X1    g234(.A(G233gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n346), .B1(new_n432), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT85), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n356), .B(new_n443), .C1(new_n346), .C2(new_n432), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n438), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT86), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n358), .A2(new_n447), .A3(new_n264), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n284), .A3(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n445), .A2(KEYINPUT87), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT87), .B1(new_n445), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n439), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(G22gat), .ZN(new_n453));
  INV_X1    g252(.A(G22gat), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n454), .B(new_n439), .C1(new_n450), .C2(new_n451), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(KEYINPUT88), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457));
  INV_X1    g256(.A(G50gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n449), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n445), .A2(KEYINPUT87), .A3(new_n449), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n464), .A2(new_n465), .B1(new_n438), .B2(new_n434), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n454), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n456), .A2(new_n461), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n453), .A2(KEYINPUT89), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n461), .B1(new_n466), .B2(new_n454), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n452), .A2(new_n472), .A3(G22gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n429), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n398), .A2(new_n405), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT35), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n301), .A2(new_n397), .A3(KEYINPUT35), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n469), .A2(new_n474), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n267), .A2(new_n288), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n291), .B2(new_n284), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT92), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT92), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n484), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n285), .A2(new_n289), .A3(new_n486), .A4(new_n292), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n298), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n293), .A2(KEYINPUT37), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n298), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n484), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n388), .A2(new_n392), .A3(new_n389), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n394), .A2(new_n396), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n403), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n355), .B1(new_n353), .B2(new_n359), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT39), .B1(new_n375), .B2(new_n376), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT39), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n504), .A2(new_n383), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n504), .A2(KEYINPUT40), .A3(new_n383), .A4(new_n506), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n509), .ZN(new_n511));
  OAI221_X1 g310(.A(new_n385), .B1(KEYINPUT40), .B2(new_n507), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n482), .B(new_n499), .C1(new_n501), .C2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n482), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n301), .A2(new_n397), .A3(KEYINPUT83), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n404), .B1(new_n399), .B2(new_n403), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n427), .A2(new_n428), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT71), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(KEYINPUT71), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n520), .A2(KEYINPUT71), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n429), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT90), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n514), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n398), .A2(new_n405), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n525), .B1(new_n530), .B2(new_n515), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT90), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n481), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT14), .B(G29gat), .Z(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538));
  NAND2_X1  g337(.A1(G43gat), .A2(G50gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT94), .B(G50gat), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(G43gat), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G43gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n458), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n538), .B1(new_n544), .B2(new_n539), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n537), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT17), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT16), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(G1gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G1gat), .B2(new_n550), .ZN(new_n553));
  INV_X1    g352(.A(G8gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n556), .A3(new_n547), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n549), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n548), .ZN(new_n560));
  INV_X1    g359(.A(new_n555), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT95), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n548), .A2(new_n555), .A3(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n558), .B(new_n559), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT18), .ZN(new_n568));
  OAI22_X1  g367(.A1(new_n562), .A2(new_n564), .B1(new_n560), .B2(new_n561), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n559), .B(KEYINPUT13), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G113gat), .B(G141gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G197gat), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT11), .B(G169gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT12), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n565), .A2(new_n566), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n568), .A2(new_n571), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT97), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n567), .A2(KEYINPUT18), .B1(new_n569), .B2(new_n570), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n577), .A4(new_n579), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n579), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n581), .A2(new_n584), .B1(new_n585), .B2(new_n576), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n533), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT7), .ZN(new_n589));
  INV_X1    g388(.A(G99gat), .ZN(new_n590));
  INV_X1    g389(.A(G106gat), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT8), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT101), .B(G92gat), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n589), .B(new_n592), .C1(G85gat), .C2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G99gat), .B(G106gat), .Z(new_n595));
  AND2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n560), .A2(new_n598), .B1(KEYINPUT41), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n594), .B(new_n595), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n549), .A2(new_n557), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n603), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT100), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n606), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G64gat), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT98), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G71gat), .B(G78gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT99), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n615), .B(new_n616), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n335), .ZN(new_n628));
  INV_X1    g427(.A(new_n623), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n561), .B1(new_n629), .B2(KEYINPUT21), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n320), .ZN(new_n633));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n636), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n612), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n623), .A2(new_n640), .A3(new_n601), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n601), .A2(new_n619), .A3(new_n622), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n598), .A2(new_n618), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n640), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT102), .B1(new_n645), .B2(new_n640), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT105), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n649), .B2(new_n645), .ZN(new_n653));
  XOR2_X1   g452(.A(G120gat), .B(G148gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT104), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n653), .A2(KEYINPUT106), .A3(new_n658), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n648), .A2(new_n663), .A3(new_n649), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n648), .B2(new_n649), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n645), .A2(new_n649), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n658), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n661), .A2(new_n662), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n639), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n587), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n390), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(G1gat), .Z(G1324gat));
  NOR4_X1   g474(.A1(new_n533), .A2(new_n586), .A3(new_n501), .A4(new_n671), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  AND2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n554), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT42), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(KEYINPUT42), .B2(new_n678), .ZN(G1325gat));
  OAI21_X1  g480(.A(G15gat), .B1(new_n673), .B2(new_n526), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n429), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n673), .B2(new_n683), .ZN(G1326gat));
  NAND3_X1  g483(.A1(new_n587), .A2(new_n515), .A3(new_n672), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT107), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n637), .A2(new_n638), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n670), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n611), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n587), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n390), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n534), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT45), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n531), .A2(new_n513), .B1(new_n477), .B2(new_n479), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(new_n611), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n691), .A2(new_n586), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n611), .A2(new_n698), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n700), .B(new_n701), .C1(new_n533), .C2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n482), .B1(new_n398), .B2(new_n405), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n528), .B1(new_n707), .B2(new_n525), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n532), .A2(new_n513), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n480), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n702), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n711), .A2(KEYINPUT108), .A3(new_n700), .A4(new_n701), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n706), .A2(new_n695), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n697), .B1(new_n534), .B2(new_n713), .ZN(G1328gat));
  INV_X1    g513(.A(G36gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n501), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n706), .A2(new_n716), .A3(new_n712), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n718), .B2(new_n717), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n693), .A2(G36gat), .A3(new_n501), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(G1329gat));
  NAND3_X1  g522(.A1(new_n694), .A2(new_n543), .A3(new_n519), .ZN(new_n724));
  OAI21_X1  g523(.A(G43gat), .B1(new_n704), .B2(new_n526), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(KEYINPUT47), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n706), .A2(new_n525), .A3(new_n712), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G43gat), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n724), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n726), .B1(new_n729), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g529(.A1(new_n482), .A2(new_n540), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n587), .A2(new_n692), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n540), .B1(new_n704), .B2(new_n482), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n706), .A2(new_n515), .A3(new_n712), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n540), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n733), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n732), .B1(new_n737), .B2(new_n540), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(KEYINPUT110), .A3(KEYINPUT48), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n735), .B1(new_n741), .B2(new_n743), .ZN(G1331gat));
  OAI21_X1  g543(.A(new_n480), .B1(new_n527), .B2(new_n514), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n661), .A2(new_n662), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n667), .A2(new_n669), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND4_X1   g547(.A1(new_n586), .A2(new_n745), .A3(new_n639), .A4(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n390), .B(KEYINPUT111), .Z(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g551(.A(new_n501), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n754), .B(new_n755), .Z(G1333gat));
  NAND2_X1  g555(.A1(new_n749), .A2(new_n519), .ZN(new_n757));
  AOI21_X1  g556(.A(G71gat), .B1(new_n757), .B2(KEYINPUT112), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(KEYINPUT112), .B2(new_n757), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n749), .A2(G71gat), .A3(new_n525), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n749), .A2(new_n515), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g563(.A1(new_n711), .A2(new_n700), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n581), .A2(new_n584), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n585), .A2(new_n576), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n689), .A2(new_n768), .A3(new_n670), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n390), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n689), .A2(new_n768), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n745), .A2(new_n612), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n670), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n390), .A2(G85gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n771), .B1(new_n778), .B2(new_n779), .ZN(G1336gat));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n716), .A3(new_n769), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n501), .A2(G92gat), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n781), .A2(new_n593), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT113), .B1(new_n781), .B2(new_n593), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(KEYINPUT52), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT52), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n770), .B2(new_n526), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n775), .A2(new_n776), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n790), .A2(new_n590), .A3(new_n519), .A4(new_n748), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1338gat));
  OAI21_X1  g591(.A(G106gat), .B1(new_n770), .B2(new_n482), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n591), .A3(new_n515), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n795), .B(new_n798), .ZN(G1339gat));
  OR2_X1    g598(.A1(new_n562), .A2(new_n564), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n559), .B1(new_n800), .B2(new_n558), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n569), .A2(new_n570), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n575), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n748), .A2(new_n766), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n658), .B1(new_n652), .B2(KEYINPUT54), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT54), .B1(new_n648), .B2(new_n651), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n806), .B(KEYINPUT55), .C1(new_n666), .C2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n648), .A2(new_n649), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT103), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n648), .A2(new_n663), .A3(new_n649), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n809), .B1(new_n813), .B2(new_n805), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n768), .A2(new_n747), .A3(new_n808), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n612), .B1(new_n804), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n808), .A3(new_n747), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n766), .A2(new_n803), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(new_n818), .A3(new_n611), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n690), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n671), .A2(new_n768), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n750), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(new_n475), .A3(new_n501), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n329), .A3(new_n768), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n515), .B1(new_n820), .B2(new_n822), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n716), .A2(new_n390), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n519), .ZN(new_n830));
  OAI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n586), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT115), .ZN(G1340gat));
  AOI21_X1  g632(.A(G120gat), .B1(new_n825), .B2(new_n748), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n670), .A2(new_n327), .A3(new_n429), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n829), .B2(new_n835), .ZN(G1341gat));
  NAND3_X1  g635(.A1(new_n825), .A2(new_n335), .A3(new_n689), .ZN(new_n837));
  OAI21_X1  g636(.A(G127gat), .B1(new_n830), .B2(new_n690), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1342gat));
  NAND3_X1  g638(.A1(new_n825), .A2(new_n333), .A3(new_n612), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT56), .Z(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n830), .B2(new_n611), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1343gat));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n817), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n814), .A2(new_n808), .A3(new_n747), .A4(KEYINPUT116), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n768), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n804), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n819), .B1(new_n848), .B2(new_n611), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n822), .B1(new_n849), .B2(new_n689), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n482), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n819), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n670), .A2(new_n818), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n586), .B1(new_n817), .B2(new_n844), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n846), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n612), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n821), .B1(new_n859), .B2(new_n690), .ZN(new_n860));
  INV_X1    g659(.A(new_n853), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT117), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n823), .A2(new_n515), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n852), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n854), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n828), .A2(new_n526), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n768), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n865), .A2(KEYINPUT118), .A3(new_n768), .A4(new_n867), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(G141gat), .A3(new_n871), .ZN(new_n872));
  AND4_X1   g671(.A1(new_n515), .A2(new_n824), .A3(new_n526), .A4(new_n501), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(new_n307), .A3(new_n768), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(KEYINPUT58), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n868), .A2(G141gat), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT58), .B1(new_n877), .B2(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1344gat));
  NOR2_X1   g678(.A1(new_n308), .A2(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n867), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n670), .ZN(new_n882));
  XNOR2_X1  g681(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n863), .A2(KEYINPUT57), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n866), .A2(new_n670), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n689), .B1(new_n859), .B2(KEYINPUT120), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n849), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n821), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n515), .A2(new_n852), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n884), .B(new_n885), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n883), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI211_X1 g693(.A(KEYINPUT121), .B(new_n883), .C1(new_n891), .C2(G148gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n882), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n873), .A2(new_n308), .A3(new_n748), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1345gat));
  OAI21_X1  g697(.A(G155gat), .B1(new_n881), .B2(new_n690), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n873), .A2(new_n320), .A3(new_n689), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1346gat));
  OAI21_X1  g700(.A(G162gat), .B1(new_n881), .B2(new_n611), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n873), .A2(new_n321), .A3(new_n612), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1347gat));
  NOR3_X1   g703(.A1(new_n501), .A2(new_n750), .A3(new_n429), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n827), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n208), .B1(new_n907), .B2(new_n768), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n695), .B1(new_n820), .B2(new_n822), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(new_n475), .A3(new_n716), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n586), .A2(G169gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT122), .Z(G1348gat));
  AOI21_X1  g712(.A(G176gat), .B1(new_n910), .B2(new_n748), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT123), .Z(new_n915));
  NOR3_X1   g714(.A1(new_n906), .A2(new_n209), .A3(new_n670), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(G1349gat));
  NAND3_X1  g716(.A1(new_n910), .A2(new_n203), .A3(new_n689), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT124), .B1(new_n906), .B2(new_n690), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G183gat), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n906), .A2(KEYINPUT124), .A3(new_n690), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n922), .B(new_n923), .Z(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n906), .B2(new_n611), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT61), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n204), .A3(new_n612), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1351gat));
  NOR3_X1   g727(.A1(new_n525), .A2(new_n482), .A3(new_n501), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n909), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n768), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n525), .A2(new_n501), .A3(new_n750), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n884), .B(new_n936), .C1(new_n889), .C2(new_n890), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n768), .A2(G197gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  NOR3_X1   g739(.A1(new_n930), .A2(G204gat), .A3(new_n670), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT62), .ZN(new_n942));
  OAI21_X1  g741(.A(G204gat), .B1(new_n937), .B2(new_n670), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n934), .A2(new_n268), .A3(new_n689), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n938), .A2(new_n689), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n947));
  OAI211_X1 g746(.A(KEYINPUT63), .B(G211gat), .C1(new_n937), .C2(new_n690), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n947), .B2(new_n949), .ZN(G1354gat));
  OAI21_X1  g749(.A(new_n269), .B1(new_n933), .B2(new_n611), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(KEYINPUT127), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(KEYINPUT127), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n269), .A3(new_n611), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G1355gat));
endmodule


