//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1236, new_n1237, new_n1238;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n461), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g047(.A1(new_n461), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(new_n461), .B2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G101), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n462), .A2(new_n463), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n478), .B1(G2105), .B2(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n480), .B(KEYINPUT69), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n461), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AOI211_X1 g067(.A(new_n486), .B(new_n489), .C1(new_n492), .C2(G136), .ZN(G162));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n462), .B2(new_n463), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  OAI21_X1  g080(.A(G138), .B1(new_n505), .B2(KEYINPUT71), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n503), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G138), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n511), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n510), .A2(new_n512), .A3(new_n461), .A4(new_n502), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n500), .B1(new_n507), .B2(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(G651), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(new_n521), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n519), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n527), .A2(G88), .B1(G50), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n532), .B(G651), .C1(new_n516), .C2(new_n522), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n524), .A2(new_n531), .A3(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  INV_X1    g111(.A(new_n526), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT77), .B(G89), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(new_n525), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT74), .B(G51), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n530), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT76), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n546));
  XNOR2_X1  g121(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n525), .A2(new_n526), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT78), .B(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n526), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G52), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n552), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n551), .A2(new_n556), .ZN(G171));
  AOI22_X1  g132(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n550), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n552), .A2(new_n560), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT79), .Z(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n520), .A2(new_n521), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n527), .B2(G91), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n530), .A2(new_n575), .A3(G53), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(G299));
  OR2_X1    g154(.A1(new_n551), .A2(new_n556), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  OAI21_X1  g156(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n525), .A2(new_n526), .A3(G87), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n526), .A2(G49), .A3(G543), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n525), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n550), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n527), .A2(G86), .B1(G48), .B2(new_n530), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n525), .A2(G60), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n550), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n527), .A2(G85), .ZN(new_n598));
  XOR2_X1   g173(.A(KEYINPUT82), .B(G47), .Z(new_n599));
  NAND2_X1  g174(.A1(new_n530), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n598), .B(new_n600), .C1(new_n594), .C2(new_n595), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT83), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n592), .A2(new_n593), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT81), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n527), .A2(G85), .B1(new_n530), .B2(new_n599), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n596), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n602), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(new_n550), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT84), .B(KEYINPUT10), .Z(new_n613));
  NAND3_X1  g188(.A1(new_n527), .A2(G92), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n530), .A2(G54), .ZN(new_n615));
  INV_X1    g190(.A(new_n613), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n552), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n612), .A2(new_n614), .A3(new_n615), .A4(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n610), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n610), .B1(new_n620), .B2(G868), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  INV_X1    g198(.A(G299), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(G868), .B2(new_n624), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(G868), .B2(new_n624), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n620), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n492), .A2(G135), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n488), .B2(G123), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n473), .A2(new_n474), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(new_n480), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT85), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n640), .A3(new_n646), .ZN(G156));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n651), .B(new_n657), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(G14), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT86), .Z(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT87), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT88), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n688), .B(new_n694), .ZN(G229));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G6), .ZN(new_n697));
  INV_X1    g272(.A(G305), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT91), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT92), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n696), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n696), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G23), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT93), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G288), .B2(new_n696), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT94), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n703), .A2(new_n707), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT34), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n492), .A2(G131), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(G107), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G2105), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n488), .B2(G119), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT90), .Z(new_n725));
  AOI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(G29), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n696), .A2(G24), .ZN(new_n730));
  INV_X1    g305(.A(G290), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n696), .ZN(new_n732));
  INV_X1    g307(.A(G1986), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n728), .A2(new_n729), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n715), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT36), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n716), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n488), .A2(G128), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n461), .A2(G116), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n492), .A2(G140), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2067), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n492), .A2(G141), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n488), .A2(G129), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  OAI21_X1  g328(.A(G105), .B1(new_n473), .B2(new_n474), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n750), .A2(new_n751), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n716), .B2(G32), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  INV_X1    g333(.A(G2072), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n716), .A2(G33), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n492), .A2(G139), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n763));
  NAND2_X1  g338(.A1(G103), .A2(G2104), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G2105), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n510), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n762), .B(new_n767), .C1(new_n461), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n761), .B1(new_n769), .B2(G29), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n757), .A2(new_n758), .B1(new_n759), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n757), .A2(new_n758), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n771), .B(new_n772), .C1(new_n759), .C2(new_n770), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n716), .A2(G35), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G162), .B2(new_n716), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT29), .B(G2090), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n638), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n716), .A2(G27), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G164), .B2(new_n716), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n778), .A2(G29), .B1(G2078), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n696), .A2(G4), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n620), .B2(new_n696), .ZN(new_n783));
  INV_X1    g358(.A(G1348), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n696), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n696), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G19), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n563), .B2(G16), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(G1341), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(G1341), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n780), .A2(G2078), .ZN(new_n794));
  INV_X1    g369(.A(G28), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT30), .ZN(new_n796));
  AOI21_X1  g371(.A(G29), .B1(new_n795), .B2(KEYINPUT30), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n796), .A2(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n793), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n781), .A2(new_n785), .A3(new_n792), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n696), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n624), .B2(new_n696), .ZN(new_n805));
  INV_X1    g380(.A(G1956), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n696), .A2(G21), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G168), .B2(new_n696), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT96), .B(G1966), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT24), .ZN(new_n812));
  INV_X1    g387(.A(G34), .ZN(new_n813));
  AOI21_X1  g388(.A(G29), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G160), .B2(new_n716), .ZN(new_n816));
  INV_X1    g391(.A(G2084), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n807), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n802), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n749), .A2(new_n773), .A3(new_n777), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n737), .A2(new_n821), .ZN(G311));
  OR2_X1    g397(.A1(new_n737), .A2(new_n821), .ZN(G150));
  AND2_X1   g398(.A1(G80), .A2(G543), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n525), .B2(G67), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n550), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n527), .A2(G93), .B1(G55), .B2(new_n530), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT97), .B1(new_n825), .B2(new_n550), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n620), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT98), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT38), .Z(new_n839));
  OR2_X1    g414(.A1(new_n559), .A2(new_n562), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n829), .B2(new_n832), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n563), .A2(new_n831), .A3(new_n828), .A4(new_n830), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n839), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n834), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n836), .B1(new_n846), .B2(new_n847), .ZN(G145));
  XOR2_X1   g423(.A(new_n638), .B(G160), .Z(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(G162), .Z(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n492), .A2(G142), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT99), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  INV_X1    g429(.A(G118), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(G2105), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n488), .A2(G130), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT100), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n853), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(G164), .B1(new_n745), .B2(new_n746), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n745), .A2(G164), .A3(new_n746), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n859), .B1(new_n865), .B2(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n769), .B(new_n755), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n724), .B(new_n643), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(new_n867), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n851), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n868), .A2(new_n871), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n867), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n850), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(G395));
  NAND2_X1  g457(.A1(G166), .A2(new_n698), .ZN(new_n883));
  NAND2_X1  g458(.A1(G303), .A2(G305), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT104), .ZN(new_n886));
  INV_X1    g461(.A(G288), .ZN(new_n887));
  NAND2_X1  g462(.A1(G290), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n602), .A2(new_n608), .A3(G288), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n890), .A3(new_n884), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n886), .A2(new_n888), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n889), .ZN(new_n893));
  AOI21_X1  g468(.A(G288), .B1(new_n602), .B2(new_n608), .ZN(new_n894));
  OAI211_X1 g469(.A(KEYINPUT104), .B(new_n885), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT105), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n843), .B(new_n629), .ZN(new_n902));
  AND2_X1   g477(.A1(G299), .A2(new_n619), .ZN(new_n903));
  NOR2_X1   g478(.A1(G299), .A2(new_n619), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(KEYINPUT102), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n906), .A2(KEYINPUT102), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT41), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n612), .A2(new_n615), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n614), .A2(new_n618), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n576), .B(KEYINPUT9), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n574), .ZN(new_n914));
  NAND2_X1  g489(.A1(G299), .A2(new_n619), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n909), .A2(new_n910), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n905), .A2(KEYINPUT103), .A3(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n920), .A2(new_n902), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n907), .B1(new_n908), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n896), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n901), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n922), .B1(new_n924), .B2(new_n901), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G868), .B2(new_n833), .ZN(G331));
  XNOR2_X1  g503(.A(G331), .B(KEYINPUT106), .ZN(G295));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n914), .A2(new_n915), .ZN(new_n931));
  INV_X1    g506(.A(new_n843), .ZN(new_n932));
  OAI21_X1  g507(.A(G301), .B1(new_n547), .B2(new_n543), .ZN(new_n933));
  INV_X1    g508(.A(new_n547), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n934), .A2(G171), .A3(new_n540), .A4(new_n542), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n931), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n843), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n938), .A2(new_n843), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n933), .A2(new_n935), .B1(new_n841), .B2(new_n842), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT107), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n941), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n946), .A2(new_n920), .A3(KEYINPUT108), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n918), .A2(new_n919), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n938), .A2(new_n843), .A3(KEYINPUT107), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT107), .B1(new_n938), .B2(new_n843), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n950), .A2(new_n951), .B1(new_n843), .B2(new_n938), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n948), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n940), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n900), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n937), .B1(new_n950), .B2(new_n951), .ZN(new_n957));
  INV_X1    g532(.A(new_n917), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n941), .A2(new_n944), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n897), .A2(new_n961), .A3(new_n899), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n876), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n930), .B1(new_n956), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  INV_X1    g540(.A(new_n940), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n946), .B2(new_n920), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n949), .A2(new_n948), .A3(new_n952), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(G37), .B1(new_n969), .B2(new_n900), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n954), .A2(new_n955), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(new_n965), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n964), .A2(KEYINPUT109), .A3(new_n972), .A4(new_n965), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n963), .B1(new_n900), .B2(new_n969), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT44), .B1(new_n978), .B2(new_n930), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n970), .A2(new_n971), .A3(new_n930), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT110), .A4(new_n930), .ZN(new_n983));
  AOI211_X1 g558(.A(KEYINPUT111), .B(new_n979), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n983), .ZN(new_n986));
  INV_X1    g561(.A(new_n979), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n977), .B1(new_n984), .B2(new_n988), .ZN(G397));
  INV_X1    g564(.A(KEYINPUT125), .ZN(new_n990));
  INV_X1    g565(.A(new_n500), .ZN(new_n991));
  AOI21_X1  g566(.A(G2105), .B1(new_n508), .B2(new_n509), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n502), .B1(new_n992), .B2(new_n512), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n504), .A2(new_n503), .A3(new_n506), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(KEYINPUT112), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(G164), .B2(G1384), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n482), .A2(G2105), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n472), .A2(new_n1002), .A3(G40), .A4(new_n477), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G164), .A2(G1384), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n998), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT119), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1961), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n997), .A2(new_n1000), .A3(new_n998), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n995), .A2(new_n996), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1003), .B1(new_n1010), .B2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1007), .A2(new_n1008), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT45), .B1(new_n997), .B2(new_n1000), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n995), .A2(KEYINPUT45), .A3(new_n996), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1004), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2078), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(KEYINPUT53), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(G164), .B2(G1384), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1004), .A2(new_n1016), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1024), .B2(G2078), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1014), .A2(new_n1020), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G171), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1019), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n478), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n461), .B1(new_n482), .B2(KEYINPUT124), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(KEYINPUT124), .B2(new_n482), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1029), .A2(new_n1016), .A3(new_n1023), .A4(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1014), .A2(new_n1032), .A3(G301), .A4(new_n1025), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1014), .A2(new_n1025), .A3(new_n1032), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G171), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(KEYINPUT54), .C1(G171), .C2(new_n1026), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n810), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1009), .A2(new_n1011), .A3(new_n817), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1042), .B2(G286), .ZN(new_n1043));
  AOI21_X1  g618(.A(G168), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT51), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(KEYINPUT51), .B2(new_n1043), .ZN(new_n1046));
  INV_X1    g621(.A(G2090), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1009), .A2(new_n1011), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1024), .A2(new_n706), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n1051));
  NAND3_X1  g626(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1054), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT113), .A3(new_n1052), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1050), .A2(new_n1055), .A3(G8), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1004), .A2(new_n997), .A3(new_n1000), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n887), .A2(G1976), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1062), .A2(G8), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1981), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n589), .A2(new_n590), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G86), .ZN(new_n1068));
  INV_X1    g643(.A(G48), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n552), .A2(new_n1068), .B1(new_n554), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G1981), .B1(new_n1070), .B2(new_n588), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1067), .A2(new_n1071), .A3(KEYINPUT49), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1063), .A3(G8), .A4(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1065), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1063), .A2(G8), .A3(new_n1064), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT52), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1058), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n995), .A2(new_n998), .A3(new_n996), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1005), .A2(KEYINPUT115), .A3(new_n998), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT112), .B1(new_n995), .B2(new_n996), .ZN(new_n1087));
  NOR3_X1   g662(.A1(G164), .A2(new_n999), .A3(G1384), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT50), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n1089), .A3(new_n1047), .A4(new_n1004), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1081), .B1(new_n1090), .B2(new_n1049), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1080), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1036), .A2(new_n1039), .A3(new_n1046), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1007), .A2(new_n784), .A3(new_n1013), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1063), .A2(G2067), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1097), .A2(KEYINPUT120), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT120), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT60), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1012), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1104), .A2(new_n1105), .A3(G1348), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1103), .B1(new_n1106), .B2(new_n1098), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1097), .A2(KEYINPUT120), .A3(new_n1099), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1102), .A2(new_n620), .A3(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT60), .B(new_n619), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1024), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1086), .A2(new_n1004), .A3(new_n1089), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n806), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n624), .A2(KEYINPUT118), .A3(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1119), .A2(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(KEYINPUT118), .ZN(new_n1122));
  NAND3_X1  g697(.A1(G299), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1113), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n1118), .B2(KEYINPUT121), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n997), .A2(new_n1000), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1003), .B1(new_n1128), .B2(KEYINPUT50), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1956), .B1(new_n1129), .B2(new_n1086), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n1116), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1126), .B1(new_n1127), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n1063), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1996), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1004), .A2(new_n1016), .A3(new_n1136), .A4(new_n1023), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n840), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT123), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT122), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT59), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1138), .B2(KEYINPUT123), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1118), .A2(new_n1125), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1124), .B1(new_n1130), .B2(new_n1116), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT61), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1111), .A2(new_n1112), .A3(new_n1133), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n619), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1096), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1042), .A2(G8), .A3(G168), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1079), .A2(new_n1065), .A3(new_n1076), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1050), .A2(G8), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1092), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1161), .A2(new_n1163), .A3(KEYINPUT117), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT117), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1058), .B(new_n1159), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1162), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1160), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1157), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1158), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1095), .B2(new_n1172), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1166), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(G288), .A2(G1976), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1076), .A2(new_n1177), .B1(new_n1066), .B2(new_n698), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1063), .A2(G8), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1058), .A2(new_n1160), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n990), .B1(new_n1156), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1161), .B(new_n1058), .C1(new_n1093), .C2(new_n1091), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT116), .B1(new_n1184), .B2(new_n1157), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1185), .A2(new_n1158), .A3(new_n1173), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1180), .B1(new_n1186), .B2(new_n1166), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1132), .B2(new_n1127), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1142), .B(KEYINPUT59), .C1(new_n1138), .C2(KEYINPUT123), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1145), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1140), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1113), .ZN(new_n1195));
  AND4_X1   g770(.A1(new_n1112), .A2(new_n1193), .A3(new_n1133), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1189), .B1(new_n1196), .B2(new_n1111), .ZN(new_n1197));
  OAI211_X1 g772(.A(KEYINPUT125), .B(new_n1187), .C1(new_n1197), .C2(new_n1096), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1046), .A2(KEYINPUT62), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1199), .A2(new_n1027), .A3(new_n1184), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1200), .B1(KEYINPUT62), .B2(new_n1046), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1183), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1023), .A2(new_n1003), .ZN(new_n1203));
  INV_X1    g778(.A(G2067), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n747), .B(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n755), .B(new_n1136), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n724), .B(new_n727), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(G290), .B(G1986), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1203), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1202), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n747), .B(G2067), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1203), .B1(new_n1212), .B2(new_n755), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1203), .A2(new_n1136), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1214), .B(KEYINPUT46), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1213), .A2(KEYINPUT127), .A3(new_n1215), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1218), .A2(KEYINPUT47), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n1221));
  INV_X1    g796(.A(new_n727), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1221), .B1(new_n725), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1205), .A2(new_n1206), .A3(new_n1223), .ZN(new_n1224));
  NOR3_X1   g799(.A1(new_n725), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1225));
  OAI22_X1  g800(.A1(new_n1224), .A2(new_n1225), .B1(G2067), .B2(new_n747), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1226), .A2(new_n1203), .ZN(new_n1227));
  AND2_X1   g802(.A1(new_n1208), .A2(new_n1203), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n731), .A2(new_n733), .A3(new_n1203), .ZN(new_n1229));
  XOR2_X1   g804(.A(new_n1229), .B(KEYINPUT48), .Z(new_n1230));
  OAI211_X1 g805(.A(new_n1220), .B(new_n1227), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g806(.A(KEYINPUT47), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1211), .A2(new_n1233), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g809(.A1(new_n964), .A2(new_n972), .ZN(new_n1236));
  INV_X1    g810(.A(G319), .ZN(new_n1237));
  NOR4_X1   g811(.A1(G229), .A2(new_n1237), .A3(G401), .A4(G227), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n880), .A2(new_n1236), .A3(new_n1238), .ZN(G225));
  INV_X1    g813(.A(G225), .ZN(G308));
endmodule


