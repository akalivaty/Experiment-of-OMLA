//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G57), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n454), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G137), .A3(new_n464), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n476), .B1(new_n473), .B2(G125), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n472), .B(new_n474), .C1(new_n477), .C2(new_n464), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n480), .A2(new_n482), .A3(new_n464), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n473), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n480), .A2(new_n482), .A3(G138), .A4(new_n464), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n473), .A2(KEYINPUT4), .A3(G138), .A4(new_n464), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n464), .B2(G114), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G102), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(new_n464), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n499), .A2(new_n501), .A3(G2104), .A4(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n480), .A2(new_n482), .A3(G126), .A4(G2105), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n504), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n497), .B1(new_n507), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(G543), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(new_n520), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(G89), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT73), .B(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n515), .A2(G63), .ZN(new_n532));
  NAND3_X1  g107(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n517), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n531), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT74), .B(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n520), .A2(new_n539), .B1(new_n540), .B2(new_n523), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n517), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n520), .A2(new_n545), .B1(new_n546), .B2(new_n523), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n519), .A2(G53), .A3(G543), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT9), .Z(new_n556));
  AOI22_X1  g131(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G91), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n557), .A2(new_n517), .B1(new_n520), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G166), .ZN(G303));
  INV_X1    g138(.A(G87), .ZN(new_n564));
  INV_X1    g139(.A(G49), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n520), .A2(new_n564), .B1(new_n565), .B2(new_n523), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n512), .A2(new_n514), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n572), .A2(KEYINPUT76), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT76), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n520), .A2(new_n579), .B1(new_n580), .B2(new_n523), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n526), .A2(G85), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n585), .B2(new_n523), .C1(new_n517), .C2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n526), .A2(G92), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n591), .A2(new_n517), .B1(new_n523), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n588), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n588), .B1(new_n594), .B2(G868), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G868), .B2(new_n560), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(G868), .B2(new_n560), .ZN(G280));
  XNOR2_X1  g174(.A(KEYINPUT77), .B(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n594), .B1(G860), .B2(new_n600), .ZN(G148));
  NAND2_X1  g176(.A1(new_n594), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g180(.A(G2100), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(KEYINPUT79), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n484), .A2(G135), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n464), .A2(G111), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT80), .Z(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n610), .A2(new_n612), .B1(G123), .B2(new_n487), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G2096), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n473), .A2(new_n469), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n606), .A2(KEYINPUT79), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n618), .B(new_n620), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n615), .B(new_n621), .C1(G2096), .C2(new_n614), .ZN(G156));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2438), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2430), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT81), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n624), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n633), .B(new_n634), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G14), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT82), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT83), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT17), .ZN(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n638), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n640), .ZN(new_n646));
  INV_X1    g221(.A(new_n642), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n647), .A2(new_n643), .A3(new_n638), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n640), .A2(new_n644), .A3(new_n638), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n646), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(new_n606), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n606), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n658), .A2(new_n659), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n657), .A3(new_n660), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n666), .C1(new_n657), .C2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n668), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G6), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n581), .B1(new_n577), .B2(G651), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT32), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1981), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(G22), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G166), .B2(new_n676), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(G1971), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(G1971), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n676), .A2(G23), .ZN(new_n686));
  INV_X1    g261(.A(G288), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n676), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT33), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT87), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n688), .B(new_n690), .Z(new_n691));
  NOR4_X1   g266(.A1(new_n681), .A2(new_n684), .A3(new_n685), .A4(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n693));
  OAI21_X1  g268(.A(KEYINPUT88), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n693), .B2(new_n692), .ZN(new_n695));
  MUX2_X1   g270(.A(G24), .B(G290), .S(G16), .Z(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(G1986), .Z(new_n697));
  AOI22_X1  g272(.A1(new_n484), .A2(G131), .B1(G119), .B2(new_n487), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n695), .A2(new_n697), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G21), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G168), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT91), .B(G1966), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT92), .ZN(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G19), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n548), .B2(G16), .ZN(new_n716));
  NOR2_X1   g291(.A1(G5), .A2(G16), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G171), .B2(G16), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n714), .B1(G1341), .B2(new_n716), .C1(G1961), .C2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G27), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G164), .B2(new_n720), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT95), .B(G2078), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(G35), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n720), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT96), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT29), .B(G2090), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n718), .A2(G1961), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G11), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n720), .A2(G33), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n484), .A2(G139), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n469), .A2(G103), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  AOI22_X1  g310(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n733), .B(new_n735), .C1(new_n464), .C2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n732), .B1(new_n737), .B2(G29), .ZN(new_n738));
  INV_X1    g313(.A(G2072), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n730), .B(new_n731), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NOR4_X1   g315(.A1(new_n719), .A2(new_n724), .A3(new_n729), .A4(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(G34), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n478), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2084), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n738), .A2(new_n739), .ZN(new_n748));
  NOR2_X1   g323(.A1(G4), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n594), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1348), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n676), .A2(G20), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT97), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT23), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G299), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT93), .B(G28), .Z(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT94), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n760), .B(new_n720), .C1(new_n758), .C2(new_n757), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n756), .B(new_n761), .C1(new_n711), .C2(new_n712), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n751), .B(new_n762), .C1(G1341), .C2(new_n716), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n741), .A2(new_n747), .A3(new_n748), .A4(new_n763), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n708), .A2(new_n709), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n720), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n484), .A2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n469), .A2(G105), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n487), .A2(G129), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT26), .Z(new_n771));
  NAND4_X1  g346(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(new_n720), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT90), .Z(new_n775));
  XOR2_X1   g350(.A(KEYINPUT27), .B(G1996), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n608), .A2(G29), .A3(new_n613), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n720), .A2(G26), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n484), .A2(G140), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n487), .A2(G128), .ZN(new_n782));
  OR2_X1    g357(.A1(G104), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(new_n720), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n780), .B(new_n787), .S(KEYINPUT28), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT89), .B(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n765), .A2(new_n778), .A3(new_n779), .A4(new_n790), .ZN(G150));
  INV_X1    g366(.A(G150), .ZN(G311));
  AOI22_X1  g367(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n517), .ZN(new_n794));
  INV_X1    g369(.A(G93), .ZN(new_n795));
  INV_X1    g370(.A(G55), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n520), .A2(new_n795), .B1(new_n796), .B2(new_n523), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G860), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT98), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT37), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n548), .B(new_n798), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n594), .A2(G559), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n805), .B(new_n806), .Z(new_n807));
  OAI21_X1  g382(.A(new_n802), .B1(new_n807), .B2(G860), .ZN(G145));
  XNOR2_X1  g383(.A(new_n786), .B(new_n772), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT99), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n495), .A2(new_n496), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n495), .B2(new_n496), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n506), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(KEYINPUT100), .B1(new_n504), .B2(new_n505), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n811), .A2(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n809), .B(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n817), .A2(KEYINPUT101), .A3(new_n737), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n737), .B(KEYINPUT101), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n487), .A2(G130), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n464), .A2(G118), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT102), .Z(new_n824));
  OAI21_X1  g399(.A(new_n821), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G142), .B2(new_n484), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n701), .B(new_n826), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n820), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n491), .B(G160), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n614), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n618), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n828), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G37), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g410(.A(G290), .B(G166), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G305), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G288), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n594), .B(G299), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT41), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n602), .B(new_n803), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n841), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n844), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n840), .A2(new_n847), .A3(KEYINPUT104), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n847), .B(KEYINPUT104), .Z(new_n849));
  AOI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(new_n840), .ZN(new_n850));
  MUX2_X1   g425(.A(new_n799), .B(new_n850), .S(G868), .Z(G295));
  MUX2_X1   g426(.A(new_n799), .B(new_n850), .S(G868), .Z(G331));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n854));
  OAI21_X1  g429(.A(G286), .B1(new_n854), .B2(G171), .ZN(new_n855));
  NAND2_X1  g430(.A1(G171), .A2(new_n854), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(new_n803), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n803), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT106), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n857), .B2(new_n803), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n841), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT107), .ZN(new_n864));
  INV_X1    g439(.A(new_n838), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n858), .A2(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n843), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT107), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n860), .A2(new_n868), .A3(new_n841), .A4(new_n862), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n864), .A2(new_n865), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n842), .B1(new_n860), .B2(new_n862), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n866), .A2(new_n846), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n838), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n833), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT109), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n870), .A2(KEYINPUT109), .A3(new_n873), .A4(new_n833), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n853), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n864), .A2(new_n867), .A3(new_n869), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n838), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n833), .A3(new_n870), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(new_n853), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT44), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT43), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n881), .B2(KEYINPUT43), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n874), .A2(KEYINPUT43), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n883), .B1(new_n888), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g464(.A(G1384), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n816), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT110), .ZN(new_n894));
  INV_X1    g469(.A(G40), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n478), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n480), .A2(new_n482), .ZN(new_n897));
  INV_X1    g472(.A(G125), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n475), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n899), .A2(G2105), .B1(G137), .B2(new_n483), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n900), .A2(KEYINPUT110), .A3(G40), .A4(new_n472), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n893), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(KEYINPUT111), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(KEYINPUT111), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G1996), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n908), .A2(KEYINPUT112), .A3(new_n772), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT112), .B1(new_n908), .B2(new_n772), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G2067), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n785), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n907), .B2(new_n773), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n911), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n701), .A2(new_n703), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n704), .B1(new_n698), .B2(new_n700), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n906), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G290), .B(G1986), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n906), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(G303), .A2(G8), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT115), .ZN(new_n924));
  INV_X1    g499(.A(G8), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n507), .A2(new_n509), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n495), .A2(new_n496), .ZN(new_n927));
  AOI21_X1  g502(.A(G1384), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT50), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT113), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n508), .B1(new_n504), .B2(new_n505), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n504), .A2(new_n508), .A3(new_n505), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n890), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT113), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT50), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(KEYINPUT114), .B(G2090), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n497), .A2(KEYINPUT99), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n495), .A2(new_n496), .A3(new_n810), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n506), .B(new_n813), .ZN(new_n943));
  AOI21_X1  g518(.A(G1384), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n902), .B1(new_n944), .B2(new_n929), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n939), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n816), .A2(KEYINPUT45), .A3(new_n890), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n896), .A2(new_n901), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n892), .B1(G164), .B2(G1384), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1971), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n925), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n924), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT49), .ZN(new_n956));
  NOR2_X1   g531(.A1(G305), .A2(G1981), .ZN(new_n957));
  INV_X1    g532(.A(G1981), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n678), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n925), .B1(new_n948), .B2(new_n944), .ZN(new_n963));
  OR3_X1    g538(.A1(new_n957), .A2(new_n956), .A3(new_n959), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n961), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n967), .B2(G288), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n687), .A2(G1976), .ZN(new_n969));
  OR3_X1    g544(.A1(new_n968), .A2(KEYINPUT52), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(KEYINPUT52), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n966), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n966), .A2(new_n970), .A3(KEYINPUT117), .A4(new_n971), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n955), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n923), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n933), .A2(new_n929), .A3(new_n890), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n896), .A3(new_n901), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n929), .B1(new_n816), .B2(new_n890), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n952), .B1(new_n981), .B2(new_n938), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n982), .B2(G8), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G2084), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n937), .A2(new_n985), .A3(new_n945), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n933), .A2(KEYINPUT45), .A3(new_n890), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n948), .B(new_n987), .C1(new_n944), .C2(KEYINPUT45), .ZN(new_n988));
  INV_X1    g563(.A(new_n712), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(G286), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n976), .A2(new_n984), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT118), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT63), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n976), .A2(new_n997), .A3(new_n984), .A4(new_n993), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n954), .B(new_n993), .C1(new_n953), .C2(new_n977), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT63), .B1(new_n1000), .B2(new_n972), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT124), .B(G1961), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n935), .B1(new_n934), .B2(KEYINPUT50), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT113), .B(new_n929), .C1(new_n933), .C2(new_n890), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n948), .B1(new_n891), .B2(KEYINPUT50), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G2078), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n893), .A2(new_n948), .A3(new_n1009), .A4(new_n987), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1008), .B1(new_n950), .B2(G2078), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G171), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT125), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT125), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1015), .A3(G171), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT62), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n478), .A2(new_n895), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n893), .A2(new_n1018), .A3(new_n947), .A4(new_n1009), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1007), .A2(G301), .A3(new_n1011), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1014), .A2(new_n1022), .A3(new_n1016), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1012), .A2(G301), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1007), .A2(G171), .A3(new_n1011), .A4(new_n1019), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(KEYINPUT54), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n816), .A2(new_n890), .A3(new_n896), .A4(new_n901), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT119), .B1(new_n1028), .B2(G2067), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n948), .A2(new_n944), .A3(new_n1030), .A4(new_n912), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1348), .B1(new_n937), .B2(new_n945), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n594), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1956), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n979), .B2(new_n980), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n560), .B(KEYINPUT57), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT56), .B(G2072), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT120), .B(new_n594), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1045), .A2(new_n1039), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n947), .A2(new_n948), .A3(new_n907), .A4(new_n949), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT58), .B(G1341), .Z(new_n1048));
  NAND2_X1  g623(.A1(new_n1028), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n548), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT59), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1053), .A3(new_n548), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1042), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1038), .A2(KEYINPUT61), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n937), .A2(new_n945), .ZN(new_n1060));
  INV_X1    g635(.A(G1348), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1060), .A2(new_n1061), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT60), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n594), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1055), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n594), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(new_n1067), .B2(new_n1034), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1044), .B(new_n1046), .C1(new_n1065), .C2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n991), .A2(KEYINPUT122), .A3(G8), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G286), .A2(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT122), .B1(new_n991), .B2(G8), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n992), .A2(new_n1078), .A3(new_n1071), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1071), .B1(new_n986), .B2(new_n990), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1081), .B(KEYINPUT121), .ZN(new_n1082));
  AOI221_X4 g657(.A(new_n1017), .B1(new_n1027), .B2(new_n1069), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT62), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(new_n1085), .A3(new_n1082), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n976), .A2(new_n984), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n999), .B(new_n1001), .C1(new_n1083), .C2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n966), .A2(new_n967), .A3(new_n687), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n963), .B1(new_n1090), .B2(new_n957), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n972), .B2(new_n954), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n921), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n906), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n915), .A2(new_n916), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n786), .A2(new_n912), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1094), .A2(G1986), .A3(G290), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT48), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n919), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n908), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1101), .A2(KEYINPUT46), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(KEYINPUT46), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1094), .B1(new_n773), .B2(new_n913), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT47), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1097), .A2(new_n1100), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1093), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT126), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1093), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g687(.A1(new_n881), .A2(KEYINPUT43), .ZN(new_n1114));
  NAND2_X1  g688(.A1(new_n1114), .A2(KEYINPUT108), .ZN(new_n1115));
  INV_X1    g689(.A(new_n887), .ZN(new_n1116));
  NAND3_X1  g690(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT43), .ZN(new_n1117));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NOR4_X1   g692(.A1(G229), .A2(G227), .A3(new_n462), .A4(G401), .ZN(new_n1119));
  INV_X1    g693(.A(KEYINPUT127), .ZN(new_n1120));
  AOI22_X1  g694(.A1(new_n1119), .A2(new_n1120), .B1(new_n833), .B2(new_n832), .ZN(new_n1121));
  OR2_X1    g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1122));
  AND3_X1   g696(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .ZN(G308));
  NAND3_X1  g697(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .ZN(G225));
endmodule


