//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G232), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n201), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  AND2_X1   g0019(.A1(KEYINPUT65), .A2(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(KEYINPUT65), .A2(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n203), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n209), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n219), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n211), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  XNOR2_X1  g0048(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n223), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n206), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n255), .A2(new_n259), .B1(new_n250), .B2(new_n257), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT7), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n222), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n207), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n265), .A2(new_n271), .A3(G68), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n265), .A2(new_n271), .A3(new_n274), .A4(G68), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT72), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(new_n201), .B2(new_n202), .ZN(new_n277));
  NAND3_X1  g0077(.A1(KEYINPUT72), .A2(G58), .A3(G68), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n203), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n279), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n273), .A2(KEYINPUT16), .A3(new_n275), .A4(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(new_n253), .ZN(new_n283));
  OR2_X1    g0083(.A1(KEYINPUT65), .A2(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT65), .A2(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT7), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n263), .A2(new_n264), .A3(new_n207), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G68), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n281), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT16), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT73), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT73), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n294), .B(KEYINPUT16), .C1(new_n290), .C2(new_n281), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n260), .B1(new_n283), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  AND2_X1   g0098(.A1(G1), .A2(G13), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G274), .ZN(new_n302));
  INV_X1    g0102(.A(G41), .ZN(new_n303));
  INV_X1    g0103(.A(G45), .ZN(new_n304));
  AOI21_X1  g0104(.A(G1), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n300), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n223), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(new_n305), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n307), .B1(G232), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G1698), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n268), .B2(new_n269), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G226), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G87), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n287), .A2(new_n312), .ZN(new_n318));
  INV_X1    g0118(.A(G223), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n287), .A2(KEYINPUT74), .A3(G223), .A4(new_n312), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT68), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n299), .B2(new_n300), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n298), .B(new_n311), .C1(new_n322), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n310), .A2(G232), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n306), .B2(new_n302), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n313), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n263), .A2(G1698), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT74), .B1(new_n332), .B2(G223), .ZN(new_n333));
  INV_X1    g0133(.A(new_n321), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n330), .B1(new_n335), .B2(new_n326), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n328), .B1(new_n336), .B2(G200), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n249), .B1(new_n297), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n260), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n291), .A2(new_n292), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n294), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n291), .A2(KEYINPUT73), .A3(new_n292), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(new_n253), .A3(new_n282), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AND4_X1   g0146(.A1(new_n339), .A2(new_n343), .A3(new_n337), .A4(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n320), .A2(new_n321), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n327), .B1(new_n349), .B2(new_n331), .ZN(new_n350));
  OAI21_X1  g0150(.A(G169), .B1(new_n350), .B2(new_n330), .ZN(new_n351));
  OAI211_X1 g0151(.A(G179), .B(new_n311), .C1(new_n322), .C2(new_n327), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT18), .B1(new_n297), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n343), .A2(new_n339), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT18), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n352), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n222), .A2(G33), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n364), .A2(new_n253), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(KEYINPUT11), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(KEYINPUT11), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT12), .B1(new_n250), .B2(G68), .ZN(new_n368));
  OR3_X1    g0168(.A1(new_n250), .A2(KEYINPUT12), .A3(G68), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n368), .A2(new_n369), .B1(new_n254), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n307), .B1(G238), .B2(new_n310), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G97), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n211), .A2(G1698), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G226), .B2(G1698), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n376), .B2(new_n263), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n326), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(new_n380), .A3(new_n378), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT70), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT14), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(G169), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n379), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT13), .ZN(new_n389));
  OAI211_X1 g0189(.A(G179), .B(new_n383), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n386), .B1(new_n384), .B2(G169), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n372), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n372), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n384), .A2(G200), .ZN(new_n395));
  OAI211_X1 g0195(.A(G190), .B(new_n383), .C1(new_n388), .C2(new_n389), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n313), .A2(G238), .B1(new_n263), .B2(G107), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n211), .B2(new_n318), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n326), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n307), .B1(G244), .B2(new_n310), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G200), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT15), .B(G87), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n362), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n280), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n222), .A2(new_n363), .B1(new_n256), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n253), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n258), .A2(G77), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n254), .A2(new_n411), .B1(new_n363), .B2(new_n251), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n404), .B(new_n414), .C1(new_n298), .C2(new_n403), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n313), .A2(G223), .B1(new_n263), .B2(G77), .ZN(new_n416));
  INV_X1    g0216(.A(G222), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n318), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n326), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT67), .B(G226), .Z(new_n420));
  AOI21_X1  g0220(.A(new_n307), .B1(new_n310), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G169), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n425));
  INV_X1    g0225(.A(G150), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n425), .B1(new_n426), .B2(new_n407), .C1(new_n362), .C2(new_n256), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n253), .ZN(new_n428));
  INV_X1    g0228(.A(G50), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n206), .B2(G20), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n254), .A2(new_n430), .B1(new_n429), .B2(new_n251), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n424), .B(new_n432), .C1(G179), .C2(new_n422), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n403), .A2(new_n423), .ZN(new_n434));
  INV_X1    g0234(.A(G179), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n401), .A2(new_n435), .A3(new_n402), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n436), .A3(new_n413), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n415), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n428), .A2(new_n431), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT9), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n422), .A2(G200), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n419), .A2(G190), .A3(new_n421), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT9), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT10), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n432), .B(KEYINPUT9), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT10), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n442), .A4(new_n441), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n438), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n360), .A2(new_n398), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT76), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT76), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n360), .A2(new_n398), .A3(new_n450), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n304), .A2(G1), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n301), .A3(G274), .A4(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n456), .B2(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n301), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n462), .B2(new_n213), .ZN(new_n463));
  OAI211_X1 g0263(.A(G244), .B(new_n312), .C1(new_n261), .C2(new_n262), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT79), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT4), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT4), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n313), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n463), .B1(new_n471), .B2(new_n326), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT80), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI211_X1 g0274(.A(KEYINPUT80), .B(new_n463), .C1(new_n471), .C2(new_n326), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n423), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n288), .A2(G107), .A3(new_n289), .ZN(new_n477));
  AND2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n478), .A2(new_n479), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(KEYINPUT6), .B2(new_n212), .ZN(new_n482));
  XNOR2_X1  g0282(.A(G97), .B(G107), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n480), .B(new_n286), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n363), .B2(new_n407), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n253), .B1(new_n477), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n206), .A2(G33), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n250), .A2(new_n487), .A3(new_n223), .A4(new_n252), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n488), .A2(KEYINPUT78), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(KEYINPUT78), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n251), .A2(new_n212), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n486), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n472), .A2(new_n435), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n476), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G200), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n472), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(new_n494), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n287), .A2(G250), .A3(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n468), .B1(new_n464), .B2(new_n465), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n327), .B1(new_n505), .B2(new_n469), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT80), .B1(new_n506), .B2(new_n463), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n472), .A2(new_n473), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(G190), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G238), .B(new_n312), .C1(new_n261), .C2(new_n262), .ZN(new_n511));
  OAI211_X1 g0311(.A(G244), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n512));
  INV_X1    g0312(.A(G116), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n511), .B(new_n512), .C1(new_n267), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n326), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n301), .A2(G274), .A3(new_n459), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n206), .A2(G45), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n301), .A2(G250), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  INV_X1    g0322(.A(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n479), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT19), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n374), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n286), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n284), .A2(G33), .A3(G97), .A4(new_n285), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n525), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n222), .A2(new_n287), .A3(G68), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n253), .B1(new_n251), .B2(new_n405), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n491), .A2(G87), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n519), .B1(new_n514), .B2(new_n326), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G190), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n522), .A2(new_n532), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n521), .A2(new_n423), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(new_n253), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n405), .A2(new_n251), .ZN(new_n539));
  INV_X1    g0339(.A(new_n405), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n489), .A2(new_n540), .A3(new_n490), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n534), .A2(new_n435), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n497), .A2(new_n510), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n461), .A2(G264), .A3(new_n301), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT83), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n461), .A2(KEYINPUT83), .A3(G264), .A4(new_n301), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G257), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n553));
  OAI211_X1 g0353(.A(G250), .B(new_n312), .C1(new_n261), .C2(new_n262), .ZN(new_n554));
  INV_X1    g0354(.A(G294), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n554), .C1(new_n267), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n326), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n552), .A2(new_n460), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n498), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n552), .A2(new_n298), .A3(new_n460), .A4(new_n557), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  INV_X1    g0362(.A(G107), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n284), .B2(new_n285), .ZN(new_n565));
  NAND2_X1  g0365(.A1(KEYINPUT23), .A2(G107), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(G20), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT82), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n567), .A2(G20), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n562), .B(new_n563), .C1(new_n220), .C2(new_n221), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n566), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n222), .A2(new_n287), .A3(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT22), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n222), .A2(new_n287), .A3(new_n577), .A4(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT24), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n574), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n574), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n253), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n491), .A2(G107), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n251), .A2(new_n563), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT25), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n561), .A2(new_n583), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n574), .A2(new_n579), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT24), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n574), .A2(new_n579), .A3(new_n580), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n588), .B1(new_n594), .B2(new_n253), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n558), .A2(new_n423), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n552), .A2(new_n435), .A3(new_n460), .A4(new_n557), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n590), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n302), .A2(new_n461), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n309), .B1(new_n458), .B2(new_n459), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(G270), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n287), .A2(G264), .A3(G1698), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n287), .A2(G257), .A3(new_n312), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n263), .A2(G303), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n326), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n423), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT81), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n251), .A2(new_n513), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n488), .B2(new_n513), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n267), .A2(G97), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n284), .A2(new_n612), .A3(new_n285), .A4(new_n502), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n252), .A2(new_n223), .B1(G20), .B2(new_n513), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT20), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(KEYINPUT20), .A3(new_n614), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n609), .B(new_n611), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  INV_X1    g0420(.A(new_n611), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT81), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n608), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n618), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT20), .B1(new_n613), .B2(new_n614), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n609), .B1(new_n628), .B2(new_n611), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n620), .A2(KEYINPUT81), .A3(new_n621), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n602), .A2(new_n607), .A3(G179), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(KEYINPUT21), .B(new_n608), .C1(new_n619), .C2(new_n622), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n602), .A2(new_n607), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G200), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n602), .A2(new_n607), .A3(G190), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(new_n629), .A3(new_n630), .A4(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n625), .A2(new_n634), .A3(new_n635), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n599), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n455), .A2(new_n547), .A3(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n433), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n449), .A2(new_n446), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n397), .A2(new_n436), .A3(new_n413), .A4(new_n434), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n393), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n338), .B2(new_n347), .ZN(new_n650));
  INV_X1    g0450(.A(new_n359), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT84), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n647), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n650), .A2(KEYINPUT84), .A3(new_n651), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n643), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n544), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n497), .B2(new_n545), .ZN(new_n660));
  AOI21_X1  g0460(.A(G169), .B1(new_n507), .B2(new_n508), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n494), .A2(new_n495), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(KEYINPUT26), .A3(new_n546), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n583), .A2(new_n589), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(new_n597), .A3(new_n596), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n634), .A2(new_n635), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n625), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n476), .A2(new_n496), .B1(new_n500), .B2(new_n509), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n546), .A4(new_n590), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n657), .B1(new_n455), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT86), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n222), .A2(new_n206), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n595), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT88), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n667), .A3(new_n590), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n598), .B1(new_n583), .B2(new_n589), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n680), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n640), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT87), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n631), .A2(new_n680), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(KEYINPUT87), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n625), .A2(new_n634), .A3(new_n635), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(new_n693), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n690), .A2(new_n695), .A3(G330), .A4(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT89), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n685), .A2(new_n686), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n681), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n701), .A2(new_n703), .B1(new_n688), .B2(new_n681), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n228), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n206), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n524), .A2(G116), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n708), .A2(new_n709), .B1(new_n226), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  NAND4_X1  g0511(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT91), .A4(new_n625), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n696), .B2(new_n688), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n547), .A2(new_n712), .A3(new_n590), .A4(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n680), .B1(new_n715), .B2(new_n665), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n680), .B1(new_n665), .B2(new_n671), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n534), .A2(new_n552), .A3(new_n557), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n632), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n507), .A2(new_n723), .A3(new_n508), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n507), .A2(new_n723), .A3(new_n508), .A4(KEYINPUT30), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n558), .A2(new_n636), .A3(new_n435), .A4(new_n521), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(new_n472), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT90), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n547), .A2(new_n641), .A3(new_n681), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n680), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT90), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n730), .A2(new_n737), .A3(KEYINPUT31), .A4(new_n680), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n732), .A2(new_n733), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n718), .B(new_n721), .C1(G330), .C2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n711), .B1(new_n740), .B2(G1), .ZN(G364));
  NAND3_X1  g0541(.A1(new_n695), .A2(G330), .A3(new_n697), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n222), .A2(G13), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G45), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n708), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n695), .A2(new_n697), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n223), .B1(G20), .B2(new_n423), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n228), .A2(new_n287), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT92), .Z(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G355), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G116), .B2(new_n228), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n706), .A2(new_n287), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G45), .B2(new_n225), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(G45), .B2(new_n247), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n755), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n745), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n222), .A2(new_n435), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G200), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT93), .Z(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n201), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n298), .A2(G179), .A3(G200), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n222), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G97), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n498), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G20), .A3(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G87), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n773), .A2(new_n287), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n498), .A2(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n766), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n778), .B1(G68), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n286), .A2(new_n298), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n767), .A2(new_n498), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G50), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n286), .A2(new_n298), .A3(new_n774), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n563), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n766), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n791), .B1(new_n794), .B2(G77), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n782), .A2(new_n787), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  INV_X1    g0597(.A(new_n784), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n781), .A2(new_n797), .B1(G329), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n790), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G322), .A2(new_n768), .B1(new_n788), .B2(G326), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n287), .B1(new_n776), .B2(G303), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT94), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(new_n804), .B1(G294), .B2(new_n772), .ZN(new_n805));
  INV_X1    g0605(.A(new_n803), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(KEYINPUT94), .B1(new_n794), .B2(G311), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n802), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n770), .A2(new_n796), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n765), .B1(new_n809), .B2(new_n754), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n749), .B1(new_n753), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NOR2_X1   g0612(.A1(new_n437), .A2(new_n680), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n415), .B1(new_n414), .B2(new_n681), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n437), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT26), .B1(new_n663), .B2(new_n546), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n661), .A2(new_n545), .A3(new_n662), .A4(new_n659), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n544), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n497), .A2(new_n510), .A3(new_n546), .A4(new_n590), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n696), .A2(new_n688), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n681), .B(new_n815), .C1(new_n818), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT96), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n719), .A2(new_n815), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n823), .B(new_n824), .Z(new_n825));
  NAND2_X1  g0625(.A1(new_n739), .A2(G330), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n745), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(new_n826), .ZN(new_n829));
  INV_X1    g0629(.A(new_n754), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G159), .A2(new_n794), .B1(new_n781), .B2(G150), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  INV_X1    g0632(.A(new_n788), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n769), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(G143), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT34), .Z(new_n837));
  INV_X1    g0637(.A(KEYINPUT95), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n790), .A2(new_n202), .ZN(new_n841));
  INV_X1    g0641(.A(new_n772), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n287), .B1(new_n429), .B2(new_n775), .C1(new_n842), .C2(new_n201), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(G132), .C2(new_n798), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n839), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n773), .B(new_n263), .C1(new_n563), .C2(new_n775), .ZN(new_n846));
  INV_X1    g0646(.A(new_n790), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(G87), .B2(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n513), .A2(new_n793), .B1(new_n780), .B2(new_n800), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G311), .B2(new_n798), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n788), .A2(G303), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n768), .A2(G294), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n848), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n830), .B1(new_n845), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n754), .A2(new_n750), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n764), .B1(G77), .B2(new_n856), .C1(new_n815), .C2(new_n751), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n828), .A2(new_n829), .B1(new_n854), .B2(new_n857), .ZN(G384));
  MUX2_X1   g0658(.A(new_n482), .B(new_n481), .S(new_n483), .Z(new_n859));
  OAI211_X1 g0659(.A(G116), .B(new_n224), .C1(new_n859), .C2(KEYINPUT35), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT97), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n859), .A2(KEYINPUT35), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n226), .A2(G77), .A3(new_n277), .A4(new_n278), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n429), .A2(G68), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n206), .B(G13), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n678), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n651), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n343), .A2(new_n337), .A3(new_n339), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n273), .A2(new_n275), .A3(new_n281), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT100), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n273), .A2(KEYINPUT100), .A3(new_n275), .A4(new_n281), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n292), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n260), .B1(new_n879), .B2(new_n283), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n874), .B1(new_n880), .B2(new_n678), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n353), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n355), .A2(new_n357), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n355), .A2(new_n872), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n874), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n880), .A2(new_n678), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n348), .B2(new_n359), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT101), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n890), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT101), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n813), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n822), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n372), .A2(new_n680), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n393), .A2(KEYINPUT99), .A3(new_n397), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT99), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n393), .A2(new_n905), .A3(new_n397), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n391), .A2(new_n392), .A3(new_n903), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n903), .A2(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n873), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT102), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT102), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n909), .B1(new_n893), .B2(new_n899), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n914), .B2(new_n873), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n891), .A2(new_n892), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n874), .B1(new_n297), .B2(new_n353), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n297), .A2(new_n678), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT37), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n887), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n919), .B1(new_n348), .B2(new_n359), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n895), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT39), .B1(new_n924), .B2(new_n898), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n393), .A2(new_n680), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n917), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n912), .A2(new_n915), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n455), .B1(new_n721), .B2(new_n718), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n656), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(KEYINPUT31), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n734), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n730), .B(new_n680), .C1(new_n934), .C2(KEYINPUT31), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n733), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n908), .A2(new_n938), .A3(new_n815), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n933), .B1(new_n900), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n924), .A2(new_n898), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT40), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n938), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n452), .B2(new_n454), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n747), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n932), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n206), .B2(new_n743), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n932), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n871), .B1(new_n951), .B2(new_n952), .ZN(G367));
  NAND2_X1  g0753(.A1(new_n494), .A2(new_n680), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n670), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT106), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n663), .A2(new_n680), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n701), .A3(new_n703), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT42), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n497), .B1(new_n956), .B2(new_n667), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n681), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(KEYINPUT42), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n533), .A2(new_n532), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n680), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n546), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n544), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT105), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n698), .B(KEYINPUT89), .ZN(new_n974));
  INV_X1    g0774(.A(new_n972), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n964), .A2(new_n975), .A3(new_n969), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n958), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n974), .A2(new_n958), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n707), .B(KEYINPUT41), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n958), .A2(new_n704), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT45), .B1(new_n958), .B2(new_n704), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n958), .A2(new_n704), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT44), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(new_n988), .A3(new_n700), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n987), .A2(KEYINPUT44), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n958), .A2(new_n704), .A3(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n990), .A2(new_n992), .B1(new_n984), .B2(new_n985), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n974), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n701), .A2(new_n703), .ZN(new_n995));
  OAI211_X1 g0795(.A(KEYINPUT107), .B(new_n995), .C1(new_n690), .C2(new_n703), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(KEYINPUT107), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(KEYINPUT108), .A3(new_n742), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n742), .A2(KEYINPUT108), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n742), .A2(KEYINPUT108), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n1000), .A2(new_n996), .A3(new_n1001), .A4(new_n997), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n989), .A2(new_n994), .A3(new_n740), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n981), .B1(new_n1004), .B2(new_n740), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n744), .A2(G1), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n977), .B(new_n980), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n760), .A2(new_n240), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n755), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n706), .B2(new_n540), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n745), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n752), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n788), .A2(G143), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n768), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n202), .B2(new_n842), .C1(new_n1014), .C2(new_n426), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT111), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n287), .B1(new_n201), .B2(new_n775), .C1(new_n784), .C2(new_n832), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n847), .A2(G77), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n780), .B2(new_n785), .C1(new_n429), .C2(new_n793), .ZN(new_n1020));
  OR3_X1    g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n794), .A2(G283), .B1(G107), .B2(new_n772), .ZN(new_n1023));
  INV_X1    g0823(.A(G311), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n1024), .B2(new_n833), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n776), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT46), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n775), .B2(new_n513), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(new_n780), .C2(new_n555), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1025), .B1(KEYINPUT109), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(KEYINPUT109), .B2(new_n1029), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n790), .A2(new_n212), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n287), .B(new_n1032), .C1(G317), .C2(new_n798), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT110), .ZN(new_n1034));
  INV_X1    g0834(.A(G303), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n769), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1021), .A2(new_n1022), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT47), .Z(new_n1038));
  OAI221_X1 g0838(.A(new_n1011), .B1(new_n1012), .B2(new_n968), .C1(new_n1038), .C2(new_n830), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1007), .A2(new_n1039), .ZN(G387));
  OAI22_X1  g0840(.A1(new_n1035), .A2(new_n793), .B1(new_n780), .B2(new_n1024), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G322), .B2(new_n788), .ZN(new_n1042));
  INV_X1    g0842(.A(G317), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n769), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n772), .A2(G283), .B1(G294), .B2(new_n776), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n790), .A2(new_n513), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n287), .B(new_n1053), .C1(G326), .C2(new_n798), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n772), .A2(new_n540), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n287), .C1(new_n363), .C2(new_n775), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT112), .B(G150), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1032), .B(new_n1057), .C1(new_n798), .C2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n202), .A2(new_n793), .B1(new_n780), .B2(new_n256), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT113), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G50), .A2(new_n768), .B1(new_n788), .B2(G159), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n830), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n760), .B1(new_n237), .B2(new_n304), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n757), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n709), .B2(new_n1066), .ZN(new_n1067));
  OR3_X1    g0867(.A1(new_n256), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1068));
  OAI21_X1  g0868(.A(KEYINPUT50), .B1(new_n256), .B2(G50), .ZN(new_n1069));
  AOI21_X1  g0869(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n709), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1067), .A2(new_n1071), .B1(new_n563), .B2(new_n706), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n764), .B1(new_n1072), .B2(new_n1009), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1064), .A2(KEYINPUT114), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n690), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n752), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT114), .B1(new_n1064), .B2(new_n1073), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1006), .A2(new_n1003), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1003), .A2(new_n740), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n707), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1003), .A2(new_n740), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(G393));
  NAND2_X1  g0882(.A1(new_n989), .A2(new_n994), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n956), .A2(new_n752), .A3(new_n957), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n760), .A2(new_n244), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1086), .B(new_n755), .C1(new_n212), .C2(new_n228), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n764), .A2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT115), .Z(new_n1089));
  AOI22_X1  g0889(.A1(G150), .A2(new_n788), .B1(new_n768), .B2(G159), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n772), .A2(G77), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n263), .B1(new_n776), .B2(G68), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G87), .B2(new_n847), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n794), .A2(new_n257), .B1(G143), .B2(new_n798), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n429), .C2(new_n780), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G311), .A2(new_n768), .B1(new_n788), .B2(G317), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT52), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n287), .B(new_n791), .C1(G116), .C2(new_n772), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n798), .A2(G322), .B1(G283), .B2(new_n776), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(KEYINPUT116), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(KEYINPUT116), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G294), .A2(new_n794), .B1(new_n781), .B2(G303), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1091), .A2(new_n1097), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1089), .B1(new_n1106), .B2(new_n754), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1084), .A2(new_n1006), .B1(new_n1085), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1083), .A2(new_n1079), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n707), .A3(new_n1004), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(G390));
  NAND4_X1  g0911(.A1(new_n908), .A2(new_n938), .A3(G330), .A4(new_n815), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT38), .B1(new_n921), .B2(new_n922), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n916), .B1(new_n891), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1115), .A2(new_n1116), .B1(new_n909), .B2(new_n926), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n926), .B1(new_n891), .B2(new_n1114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n814), .A2(new_n437), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n813), .B1(new_n716), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1118), .B1(new_n1121), .B2(new_n908), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1113), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n813), .B1(new_n719), .B2(new_n815), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n908), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n926), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n917), .B2(new_n925), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n942), .B(new_n926), .C1(new_n1120), .C2(new_n1125), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n739), .A2(new_n908), .A3(G330), .A4(new_n815), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1123), .A2(new_n1006), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n750), .B1(new_n917), .B2(new_n925), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n764), .B1(new_n257), .B2(new_n856), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n212), .A2(new_n793), .B1(new_n780), .B2(new_n563), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G294), .B2(new_n798), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n788), .A2(G283), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n768), .A2(G116), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1092), .A2(new_n263), .A3(new_n777), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1138), .A2(new_n841), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n776), .A2(new_n1058), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT120), .Z(new_n1142));
  OR2_X1    g0942(.A1(new_n1142), .A2(KEYINPUT53), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(KEYINPUT53), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1144), .C1(new_n1145), .C2(new_n833), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n287), .B1(new_n842), .B2(new_n785), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G50), .B2(new_n847), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  INV_X1    g0949(.A(G125), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n793), .A2(new_n1149), .B1(new_n1150), .B2(new_n784), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G137), .B2(new_n781), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n768), .A2(G132), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1148), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1140), .B1(new_n1146), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1133), .B1(new_n1155), .B2(new_n754), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1132), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT117), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n938), .A2(new_n1158), .A3(G330), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n815), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1158), .B1(new_n938), .B2(G330), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1125), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1129), .A2(new_n1120), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n739), .A2(G330), .A3(new_n815), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1165), .A2(new_n1125), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n902), .B1(new_n1166), .B2(new_n1113), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n455), .A2(G330), .A3(new_n938), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n930), .A2(new_n656), .A3(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1123), .A2(new_n1168), .A3(new_n1130), .A4(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(new_n707), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(KEYINPUT118), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1123), .A2(new_n1130), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1171), .A2(KEYINPUT118), .A3(new_n707), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT119), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1174), .A2(new_n1175), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1131), .B(new_n1157), .C1(new_n1173), .C2(new_n1181), .ZN(G378));
  NAND2_X1  g0982(.A1(new_n646), .A2(new_n433), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n439), .A2(new_n678), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n646), .B(new_n433), .C1(new_n439), .C2(new_n678), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n944), .A2(new_n942), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(G330), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n941), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n747), .B1(new_n944), .B2(new_n942), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n939), .B1(new_n893), .B2(new_n899), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1196), .B(new_n1197), .C1(new_n1198), .C2(new_n933), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n929), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n927), .B1(new_n911), .B2(KEYINPUT102), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1195), .A2(new_n1202), .A3(new_n915), .A4(new_n1199), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1006), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n856), .A2(G50), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n793), .A2(new_n405), .B1(new_n201), .B2(new_n790), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT121), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n303), .B(new_n263), .C1(new_n775), .C2(new_n363), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G107), .A2(new_n768), .B1(new_n788), .B2(G116), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n842), .A2(new_n202), .B1(new_n780), .B2(new_n212), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1209), .A2(new_n1208), .B1(new_n800), .B2(new_n784), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1210), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n263), .A2(new_n303), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G50), .B1(new_n267), .B2(new_n303), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1215), .A2(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n781), .A2(G132), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n426), .B2(new_n842), .C1(new_n775), .C2(new_n1149), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1150), .A2(new_n833), .B1(new_n1014), .B2(new_n1145), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(G137), .C2(new_n794), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n267), .B(new_n303), .C1(new_n790), .C2(new_n785), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G124), .B2(new_n798), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT59), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1219), .B1(new_n1216), .B2(new_n1215), .C1(new_n1225), .C2(new_n1229), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n745), .B(new_n1206), .C1(new_n1230), .C2(new_n754), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1196), .B2(new_n751), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1205), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1200), .A2(new_n929), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1199), .A2(new_n1195), .B1(new_n1202), .B2(new_n915), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT122), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT122), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1204), .A2(new_n1241), .A3(new_n1236), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1201), .A2(new_n1203), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n707), .B1(new_n1244), .B2(KEYINPUT57), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1234), .B1(new_n1243), .B2(new_n1245), .ZN(G375));
  INV_X1    g1046(.A(KEYINPUT123), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1168), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1006), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1168), .A2(KEYINPUT123), .A3(new_n1006), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n563), .A2(new_n793), .B1(new_n780), .B2(new_n513), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G294), .B2(new_n788), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT124), .Z(new_n1254));
  AOI21_X1  g1054(.A(new_n287), .B1(new_n776), .B2(G97), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1019), .A2(new_n1056), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G303), .B2(new_n798), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1254), .B(new_n1257), .C1(new_n800), .C2(new_n1014), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n263), .B1(new_n776), .B2(G159), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n201), .B2(new_n790), .C1(new_n842), .C2(new_n429), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G132), .B2(new_n788), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n793), .A2(new_n426), .B1(new_n1145), .B2(new_n784), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1149), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n781), .B2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1261), .B(new_n1264), .C1(new_n769), .C2(new_n832), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n830), .B1(new_n1258), .B2(new_n1265), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n745), .B(new_n1266), .C1(new_n202), .C2(new_n855), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n908), .B2(new_n751), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1250), .A2(new_n1251), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n981), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1175), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(G381));
  OAI211_X1 g1074(.A(new_n811), .B(new_n1078), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1275), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G378), .A2(new_n1276), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g1077(.A1(new_n679), .A2(G213), .ZN(new_n1278));
  OR3_X1    g1078(.A1(G375), .A2(G378), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(G407), .A2(G213), .A3(new_n1279), .ZN(G409));
  XNOR2_X1  g1080(.A(G393), .B(new_n811), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G387), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1007), .B2(new_n1039), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G390), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1282), .B(G390), .C1(new_n1284), .C2(new_n1281), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1289), .B(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G378), .B(new_n1234), .C1(new_n1243), .C2(new_n1245), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1131), .A2(new_n1157), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1181), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1172), .A2(KEYINPUT118), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1244), .A2(new_n1272), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1233), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1292), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G384), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1301), .A2(new_n1271), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n707), .B1(new_n1301), .B2(new_n1271), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1300), .B1(new_n1304), .B2(new_n1269), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1270), .B(G384), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1299), .A2(new_n1278), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT125), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1299), .A2(KEYINPUT125), .A3(new_n1278), .A4(new_n1308), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT62), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1299), .A2(new_n1278), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n679), .A2(G213), .A3(G2897), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1307), .B(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT61), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1291), .B1(new_n1313), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1311), .A2(new_n1321), .A3(new_n1312), .ZN(new_n1322));
  OR2_X1    g1122(.A1(new_n1309), .A2(new_n1321), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1322), .A2(new_n1323), .A3(new_n1317), .A4(new_n1289), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1320), .A2(new_n1324), .ZN(G405));
  NAND2_X1  g1125(.A1(G375), .A2(new_n1296), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1292), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1308), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1326), .A2(new_n1307), .A3(new_n1292), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  XOR2_X1   g1130(.A(new_n1330), .B(new_n1289), .Z(G402));
endmodule


