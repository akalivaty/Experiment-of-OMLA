//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT67), .B(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n470), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OAI221_X1 g053(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n478), .B(new_n479), .C1(new_n480), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n469), .A2(new_n472), .A3(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n486), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(new_n482), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT4), .A2(G138), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n463), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n492), .B(new_n496), .C1(new_n470), .C2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n510), .A2(new_n511), .B1(new_n504), .B2(new_n505), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n511), .A2(new_n510), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G62), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n513), .B1(G651), .B2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n507), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n506), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n514), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G168));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n507), .A2(new_n533), .B1(new_n534), .B2(new_n512), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  OAI211_X1 g114(.A(G43), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT71), .B(G81), .Z(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n512), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n514), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n537), .B1(new_n545), .B2(KEYINPUT70), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n547), .B(new_n543), .C1(new_n514), .C2(new_n544), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n542), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NOR2_X1   g129(.A1(new_n504), .A2(new_n505), .ZN(new_n555));
  INV_X1    g130(.A(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n557), .A2(KEYINPUT72), .A3(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n514), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n512), .ZN(new_n563));
  AOI22_X1  g138(.A1(G651), .A2(new_n562), .B1(new_n563), .B2(G91), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n559), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(new_n513), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n523), .A2(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G303));
  AOI22_X1  g145(.A1(G87), .A2(new_n563), .B1(new_n557), .B2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(G288));
  INV_X1    g151(.A(G48), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n507), .A2(new_n577), .B1(new_n578), .B2(new_n512), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n537), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(G305));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  XOR2_X1   g160(.A(KEYINPUT75), .B(G85), .Z(new_n586));
  OAI22_X1  g161(.A1(new_n507), .A2(new_n585), .B1(new_n512), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n537), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n563), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n514), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n557), .B2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G297));
  XNOR2_X1  g181(.A(G297), .B(KEYINPUT76), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  AOI21_X1  g184(.A(new_n544), .B1(new_n517), .B2(new_n518), .ZN(new_n610));
  INV_X1    g185(.A(new_n543), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT70), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n612), .A2(G651), .A3(new_n548), .ZN(new_n613));
  INV_X1    g188(.A(new_n542), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n604), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n600), .A2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n477), .A2(G135), .ZN(new_n620));
  OAI221_X1 g195(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n621));
  INV_X1    g196(.A(G123), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n487), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT78), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND2_X1  g200(.A1(KEYINPUT77), .A2(G2100), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n482), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  NOR2_X1   g204(.A1(KEYINPUT77), .A2(G2100), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n625), .B(new_n631), .C1(new_n629), .C2(new_n626), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT79), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(KEYINPUT81), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n651), .B(KEYINPUT82), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n649), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n649), .A2(new_n656), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n649), .A2(new_n656), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n651), .B(KEYINPUT17), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n674), .A2(KEYINPUT83), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(KEYINPUT83), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(KEYINPUT20), .A3(new_n676), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n670), .A2(new_n671), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n669), .B2(new_n672), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n669), .A2(KEYINPUT84), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT85), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n667), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n691), .A3(new_n666), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  OAI221_X1 g275(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT87), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n477), .A2(G131), .ZN(new_n703));
  INV_X1    g278(.A(new_n487), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G119), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n700), .B1(new_n707), .B2(new_n698), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n708), .A2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G24), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n590), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1986), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G6), .B(G305), .S(G16), .Z(new_n718));
  XOR2_X1   g293(.A(KEYINPUT32), .B(G1981), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n713), .A2(G23), .ZN(new_n721));
  INV_X1    g296(.A(G288), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n713), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT33), .B(G1976), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n713), .A2(G22), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT88), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G303), .B2(G16), .ZN(new_n728));
  INV_X1    g303(.A(G1971), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n725), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n720), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n711), .B(new_n717), .C1(new_n733), .C2(KEYINPUT34), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n734), .A2(new_n735), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n738), .A2(new_n737), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n736), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n698), .A2(G32), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n477), .A2(G141), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT26), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(G105), .B2(new_n461), .ZN(new_n754));
  INV_X1    g329(.A(G129), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n749), .B(new_n754), .C1(new_n755), .C2(new_n487), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n748), .B1(new_n761), .B2(new_n698), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n762), .B(new_n763), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n713), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n713), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n713), .A2(G5), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G171), .B2(new_n713), .ZN(new_n768));
  AOI22_X1  g343(.A1(G1966), .A2(new_n766), .B1(new_n768), .B2(G1961), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G1961), .B2(new_n768), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT31), .B(G11), .Z(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT96), .B(G28), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT30), .ZN(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n772), .B2(KEYINPUT30), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT24), .ZN(new_n776));
  INV_X1    g351(.A(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(G29), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G160), .B2(new_n698), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n775), .B1(new_n780), .B2(G2084), .C1(new_n766), .C2(G1966), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n770), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G27), .A2(G29), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G164), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2078), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G2084), .B2(new_n780), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n782), .B(new_n786), .C1(new_n698), .C2(new_n624), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n764), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n698), .A2(G33), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT25), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n477), .A2(G139), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n469), .A2(new_n472), .A3(G127), .ZN(new_n797));
  INV_X1    g372(.A(G115), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n460), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(new_n486), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n795), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(KEYINPUT92), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n793), .A2(new_n794), .B1(new_n486), .B2(new_n799), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n796), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n790), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n801), .A2(KEYINPUT92), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n804), .A2(new_n803), .A3(new_n796), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT93), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n789), .B1(new_n810), .B2(new_n698), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n788), .B1(G2072), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(G2072), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  OR3_X1    g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n813), .B1(new_n812), .B2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n713), .A2(G4), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n601), .B2(new_n713), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G1348), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n698), .A2(G26), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n477), .A2(G140), .ZN(new_n824));
  OAI221_X1 g399(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n825));
  INV_X1    g400(.A(G128), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n487), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n823), .B1(new_n828), .B2(new_n698), .ZN(new_n829));
  INV_X1    g404(.A(G2067), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n713), .A2(G19), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n549), .B2(new_n713), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(G1341), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n713), .A2(G20), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT23), .Z(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G299), .B2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1956), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n820), .A2(new_n831), .A3(new_n834), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G29), .A2(G35), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G162), .B2(G29), .ZN(new_n841));
  INV_X1    g416(.A(G2090), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n816), .A2(new_n817), .A3(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n743), .A2(new_n747), .A3(new_n847), .ZN(G311));
  NOR2_X1   g423(.A1(new_n747), .A2(new_n847), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n746), .A2(new_n741), .A3(new_n736), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(G150));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  OAI211_X1 g427(.A(G55), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n512), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(G67), .B1(new_n511), .B2(new_n510), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n537), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n852), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n517), .B2(new_n518), .ZN(new_n861));
  INV_X1    g436(.A(new_n857), .ZN(new_n862));
  OAI21_X1  g437(.A(G651), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n506), .A2(G93), .A3(new_n519), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT100), .A4(new_n853), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(new_n853), .A3(new_n864), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n613), .A2(new_n869), .A3(new_n614), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n866), .B2(new_n549), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT101), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n873), .B(new_n870), .C1(new_n866), .C2(new_n549), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT102), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n600), .A2(new_n608), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n881));
  INV_X1    g456(.A(G860), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n880), .B2(KEYINPUT39), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n868), .B1(new_n881), .B2(new_n883), .ZN(G145));
  XNOR2_X1  g459(.A(new_n624), .B(G160), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G162), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n828), .A2(new_n502), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n827), .A2(G164), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n761), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n887), .B(new_n888), .C1(new_n758), .C2(new_n760), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n810), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n889), .A2(new_n756), .B1(new_n807), .B2(new_n808), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n757), .A3(new_n888), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n895), .A3(new_n706), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n706), .B1(new_n892), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n628), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n892), .A2(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n707), .ZN(new_n901));
  INV_X1    g476(.A(new_n628), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n477), .A2(G142), .ZN(new_n904));
  INV_X1    g479(.A(G130), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(new_n905), .B2(new_n487), .ZN(new_n906));
  OAI21_X1  g481(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(KEYINPUT104), .Z(new_n908));
  OAI21_X1  g483(.A(KEYINPUT103), .B1(new_n463), .B2(G118), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n463), .A2(KEYINPUT103), .A3(G118), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n899), .A2(new_n903), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n899), .B2(new_n903), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n886), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n899), .A2(new_n903), .ZN(new_n917));
  INV_X1    g492(.A(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n886), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n899), .A2(new_n903), .A3(new_n913), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n916), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g500(.A1(new_n866), .A2(new_n604), .ZN(new_n926));
  XNOR2_X1  g501(.A(G166), .B(new_n590), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G305), .A2(G288), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(G305), .A2(G288), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n927), .A3(new_n929), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n875), .B(new_n617), .ZN(new_n937));
  NAND2_X1  g512(.A1(G299), .A2(new_n600), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n559), .A2(new_n595), .A3(new_n564), .A4(new_n599), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n940), .B2(KEYINPUT41), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n940), .B2(new_n937), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n936), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n926), .B1(new_n947), .B2(new_n604), .ZN(G295));
  OAI21_X1  g523(.A(new_n926), .B1(new_n947), .B2(new_n604), .ZN(G331));
  INV_X1    g524(.A(new_n940), .ZN(new_n950));
  INV_X1    g525(.A(new_n874), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n615), .A2(new_n859), .A3(new_n865), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n873), .B1(new_n952), .B2(new_n870), .ZN(new_n953));
  OAI21_X1  g528(.A(G171), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n872), .A2(G301), .A3(new_n874), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(G168), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G168), .B1(new_n954), .B2(new_n955), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G286), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n944), .A3(new_n956), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n935), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n963), .A2(new_n923), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT41), .B1(new_n938), .B2(new_n939), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n950), .B2(new_n942), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n961), .A2(new_n967), .A3(new_n956), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n959), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n935), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT106), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n972), .B(new_n935), .C1(new_n959), .C2(new_n968), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n964), .B(new_n965), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT107), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n961), .A2(new_n956), .A3(new_n967), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n940), .B1(new_n961), .B2(new_n956), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n970), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n972), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n969), .A2(KEYINPUT106), .A3(new_n970), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n965), .A4(new_n964), .ZN(new_n983));
  INV_X1    g558(.A(new_n964), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n935), .B1(new_n959), .B2(new_n962), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n975), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n965), .B1(new_n984), .B2(new_n985), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n981), .A2(KEYINPUT43), .A3(new_n964), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n989), .A2(new_n993), .ZN(G397));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n502), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n475), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n481), .A2(G137), .A3(new_n463), .ZN(new_n1000));
  XOR2_X1   g575(.A(KEYINPUT108), .B(G40), .Z(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n999), .A2(new_n1000), .A3(new_n462), .A4(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1996), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n1006), .A3(new_n1004), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT109), .Z(new_n1008));
  XNOR2_X1  g583(.A(new_n827), .B(new_n830), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1006), .B2(new_n757), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(new_n709), .A3(new_n707), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n828), .A2(new_n830), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1005), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1005), .B1(new_n1009), .B2(new_n757), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1016), .A2(KEYINPUT46), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(KEYINPUT46), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  XNOR2_X1  g595(.A(new_n706), .B(new_n710), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1004), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1011), .A2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1005), .A2(G1986), .A3(G290), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1020), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1014), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(G166), .B2(new_n1028), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n471), .A2(new_n475), .A3(new_n1001), .ZN(new_n1034));
  OAI22_X1  g609(.A1(new_n486), .A2(new_n499), .B1(new_n497), .B2(new_n482), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n495), .B1(new_n1035), .B2(new_n481), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1384), .B1(new_n1036), .B2(new_n492), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(KEYINPUT110), .A3(new_n1038), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n842), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n998), .A2(new_n1034), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n729), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1028), .B(new_n1033), .C1(new_n1044), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1037), .A2(new_n1034), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1050), .B(G8), .C1(new_n1051), .C2(G288), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT112), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n996), .A2(new_n1003), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(new_n1028), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n722), .A2(G1976), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1053), .ZN(new_n1060));
  AOI22_X1  g635(.A1(G86), .A2(new_n563), .B1(new_n557), .B2(G48), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1061), .B(new_n1062), .C1(new_n537), .C2(new_n580), .ZN(new_n1063));
  OAI21_X1  g638(.A(G1981), .B1(new_n579), .B2(new_n581), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1063), .A2(KEYINPUT49), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT49), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1055), .A2(new_n1060), .B1(new_n1057), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1052), .A2(KEYINPUT111), .A3(KEYINPUT52), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1068), .A2(new_n1073), .A3(KEYINPUT113), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT113), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1049), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g651(.A(G1976), .B(G288), .C1(new_n1067), .C2(new_n1057), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1063), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1057), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(new_n1049), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1003), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1048), .B1(G2090), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT114), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1048), .B(new_n1088), .C1(G2090), .C2(new_n1085), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(G8), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1033), .ZN(new_n1091));
  INV_X1    g666(.A(G1966), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n502), .A2(KEYINPUT115), .A3(KEYINPUT45), .A4(new_n995), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(new_n1034), .C1(KEYINPUT45), .C2(new_n1037), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT115), .B1(new_n1037), .B2(KEYINPUT45), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT116), .B(G2084), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT110), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1098));
  AND4_X1   g673(.A1(KEYINPUT110), .A2(new_n502), .A3(new_n1038), .A4(new_n995), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1083), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1028), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G168), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1082), .A2(new_n1091), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1049), .A2(new_n1105), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1102), .B1(new_n1109), .B2(new_n1033), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1107), .B(new_n1110), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1080), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1096), .A2(G168), .A3(new_n1100), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(G8), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT121), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT51), .B1(new_n1114), .B2(G8), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1114), .A2(new_n1120), .A3(G8), .A4(new_n1115), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1101), .A2(G286), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1113), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1114), .A2(G8), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT121), .B(new_n1116), .C1(new_n1125), .C2(KEYINPUT51), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1123), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(KEYINPUT122), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1056), .A2(new_n830), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT118), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1043), .A2(G1348), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n601), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n559), .B(new_n564), .C1(KEYINPUT117), .C2(KEYINPUT57), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT57), .B1(new_n564), .B2(KEYINPUT117), .ZN(new_n1136));
  NAND2_X1  g711(.A1(G299), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1003), .B1(new_n996), .B2(new_n997), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT56), .B(G2072), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1046), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1956), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1135), .B(new_n1137), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1134), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1142), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1137), .A2(new_n1135), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(new_n1140), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1131), .B(KEYINPUT118), .Z(new_n1152));
  NOR2_X1   g727(.A1(new_n600), .A2(KEYINPUT60), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1152), .B(new_n1153), .C1(G1348), .C2(new_n1043), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1143), .A2(new_n1147), .A3(KEYINPUT61), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT119), .B(G1996), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1138), .A2(new_n1046), .A3(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT58), .B(G1341), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1050), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n615), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1152), .B(new_n600), .C1(G1348), .C2(new_n1043), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1134), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1148), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(G2078), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n998), .A2(new_n1168), .A3(new_n1046), .A4(new_n1034), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT53), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT115), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1046), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1138), .A2(new_n1173), .A3(new_n1093), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1170), .A2(G2078), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT123), .B(G1961), .ZN(new_n1177));
  OAI221_X1 g752(.A(new_n1171), .B1(new_n1174), .B2(new_n1176), .C1(new_n1043), .C2(new_n1177), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1178), .A2(G171), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1175), .A2(G40), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT124), .B1(new_n473), .B2(new_n474), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1181), .A2(new_n463), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n473), .A2(KEYINPUT124), .A3(new_n474), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1180), .B(new_n471), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n998), .A2(new_n1184), .A3(new_n1046), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1171), .B(new_n1185), .C1(new_n1043), .C2(new_n1177), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(G171), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1179), .A2(KEYINPUT125), .A3(KEYINPUT54), .A4(new_n1187), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1187), .B(KEYINPUT54), .C1(G171), .C2(new_n1178), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1178), .A2(G171), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1043), .A2(new_n1177), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(G301), .A3(new_n1171), .A4(new_n1185), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT54), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1108), .A2(G8), .A3(new_n1032), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1197), .A2(new_n1073), .A3(new_n1068), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1028), .B1(new_n1086), .B2(KEYINPUT114), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1032), .B1(new_n1199), .B2(new_n1089), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1196), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1167), .A2(new_n1192), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1112), .B1(new_n1130), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n1129), .B2(KEYINPUT62), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1124), .A2(new_n1206), .A3(new_n1128), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1198), .A2(new_n1200), .A3(new_n1193), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1129), .A2(new_n1204), .A3(KEYINPUT62), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1203), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n590), .B(G1986), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1011), .B(new_n1022), .C1(new_n1005), .C2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1027), .B1(new_n1212), .B2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g790(.A(G319), .ZN(new_n1217));
  NOR3_X1   g791(.A1(G401), .A2(G227), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g792(.A1(new_n694), .A2(new_n696), .A3(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g793(.A(new_n1219), .B(KEYINPUT127), .ZN(new_n1220));
  AND3_X1   g794(.A1(new_n1220), .A2(new_n987), .A3(new_n924), .ZN(G308));
  NAND3_X1  g795(.A1(new_n1220), .A2(new_n987), .A3(new_n924), .ZN(G225));
endmodule


