//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n206), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n203), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n202), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n212), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n215), .B(new_n220), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n232), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  OAI21_X1  g0051(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n210), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  XOR2_X1   g0059(.A(KEYINPUT8), .B(G58), .Z(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n210), .A2(G33), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n252), .B1(new_n253), .B2(new_n259), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n266), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n218), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT68), .ZN(new_n269));
  INV_X1    g0069(.A(G50), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n271), .A2(new_n210), .A3(G1), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n263), .A2(new_n269), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n268), .B(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n209), .A2(G20), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n275), .A2(G50), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n255), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G223), .A3(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G77), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G222), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n284), .B1(new_n285), .B2(new_n283), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  OAI211_X1 g0095(.A(G1), .B(G13), .C1(new_n255), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n293), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n294), .B1(G226), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n279), .B(new_n302), .C1(G179), .C2(new_n300), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n291), .B2(new_n299), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT10), .B1(new_n306), .B2(KEYINPUT71), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n279), .B(KEYINPUT9), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n306), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(new_n307), .A3(new_n311), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n255), .A2(G20), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n259), .B2(new_n270), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n269), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n269), .A2(KEYINPUT73), .A3(new_n318), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(KEYINPUT11), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(KEYINPUT11), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n276), .A2(G68), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n326));
  NAND2_X1  g0126(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n268), .A2(new_n272), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n203), .B1(new_n209), .B2(G20), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n324), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n227), .A2(G1698), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n283), .B(new_n336), .C1(G226), .C2(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n290), .ZN(new_n340));
  INV_X1    g0140(.A(G45), .ZN(new_n341));
  AOI21_X1  g0141(.A(G1), .B1(new_n295), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n296), .A2(G274), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n297), .B2(new_n222), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n335), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n296), .B1(new_n337), .B2(new_n338), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n347), .A2(KEYINPUT13), .A3(new_n344), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n334), .B(G169), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n340), .A2(new_n335), .A3(new_n345), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT13), .B1(new_n347), .B2(new_n344), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(G179), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n301), .B1(new_n350), .B2(new_n351), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(new_n334), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT75), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n349), .A2(new_n352), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n358), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n333), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(G200), .B1(new_n346), .B2(new_n348), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT72), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n325), .A2(new_n332), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n350), .A2(G190), .A3(new_n351), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n363), .A2(new_n324), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n283), .A2(G238), .A3(G1698), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n367), .B1(new_n368), .B2(new_n283), .C1(new_n287), .C2(new_n227), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n290), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n294), .B1(G244), .B2(new_n298), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n301), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G179), .B2(new_n372), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n330), .A2(G77), .A3(new_n277), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G77), .B2(new_n276), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n260), .A2(new_n258), .B1(G20), .B2(G77), .ZN(new_n377));
  XOR2_X1   g0177(.A(KEYINPUT15), .B(G87), .Z(new_n378));
  AOI22_X1  g0178(.A1(new_n377), .A2(KEYINPUT70), .B1(new_n316), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(KEYINPUT70), .B2(new_n377), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n376), .B1(new_n380), .B2(new_n268), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n372), .A2(G200), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n381), .B(new_n384), .C1(new_n309), .C2(new_n372), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n315), .A2(new_n361), .A3(new_n366), .A4(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n296), .A2(G232), .A3(new_n293), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n343), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT77), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n286), .A2(G226), .ZN(new_n392));
  OR2_X1    g0192(.A1(G223), .A2(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(KEYINPUT3), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT3), .A2(G33), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n394), .A2(new_n397), .B1(new_n255), .B2(new_n223), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n290), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n343), .A2(new_n389), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n391), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G169), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n391), .A2(new_n399), .A3(G179), .A4(new_n401), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT78), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT78), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n260), .A2(new_n277), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n275), .A2(new_n276), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n276), .B2(new_n260), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n265), .A2(new_n218), .A3(new_n267), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT7), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n283), .B2(G20), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G68), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n258), .A2(G159), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G20), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT76), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(KEYINPUT76), .A3(G20), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n418), .A2(new_n419), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT16), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n413), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n417), .A2(G68), .B1(G159), .B2(new_n258), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n428), .A2(KEYINPUT16), .A3(new_n423), .A4(new_n424), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n412), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n409), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT80), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n402), .A2(new_n305), .ZN(new_n435));
  AND2_X1   g0235(.A1(KEYINPUT79), .A2(G190), .ZN(new_n436));
  NOR2_X1   g0236(.A1(KEYINPUT79), .A2(G190), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n435), .B1(new_n402), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n430), .A2(new_n434), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n441), .B(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n388), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT87), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G116), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(G20), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n210), .A2(KEYINPUT87), .A3(G33), .A4(G116), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT23), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n210), .B2(G107), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n368), .A2(KEYINPUT23), .A3(G20), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n448), .A2(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n210), .B(G87), .C1(new_n395), .C2(new_n396), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT24), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT24), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n453), .C1(new_n455), .C2(new_n456), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n413), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT89), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n272), .A2(new_n463), .A3(new_n368), .ZN(new_n464));
  XOR2_X1   g0264(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n272), .B2(new_n368), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n255), .A2(G1), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n269), .A2(new_n272), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n462), .A2(new_n471), .A3(KEYINPUT90), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT90), .ZN(new_n473));
  INV_X1    g0273(.A(new_n467), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n466), .B(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n469), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n275), .A2(new_n276), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n477), .B2(new_n368), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n473), .B1(new_n478), .B2(new_n461), .ZN(new_n479));
  OR2_X1    g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n341), .A2(G1), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G264), .A3(new_n296), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n290), .A2(new_n292), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n209), .A2(G45), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n480), .B2(new_n481), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(G250), .A2(G1698), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n229), .B2(G1698), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(new_n283), .B1(G33), .B2(G294), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n485), .B(new_n489), .C1(new_n492), .C2(new_n296), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G169), .ZN(new_n494));
  INV_X1    g0294(.A(G179), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n493), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n472), .A2(new_n479), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n458), .A2(new_n460), .ZN(new_n498));
  INV_X1    g0298(.A(new_n492), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n488), .A2(new_n290), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n499), .A2(new_n290), .B1(G264), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n309), .A3(new_n489), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n305), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n498), .A2(new_n268), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n471), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(new_n286), .C1(new_n395), .C2(new_n396), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G250), .A2(G1698), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT4), .A2(G244), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(G1698), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n283), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT84), .B1(new_n516), .B2(new_n290), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  AOI211_X1 g0318(.A(new_n518), .B(new_n296), .C1(new_n509), .C2(new_n515), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n500), .A2(G257), .B1(new_n486), .B2(new_n488), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n275), .A2(G97), .A3(new_n276), .A4(new_n476), .ZN(new_n524));
  INV_X1    g0324(.A(new_n257), .ZN(new_n525));
  NOR3_X1   g0325(.A1(KEYINPUT69), .A2(G20), .A3(G33), .ZN(new_n526));
  OAI21_X1  g0326(.A(G77), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT81), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n258), .A2(new_n529), .A3(G77), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT7), .B1(new_n397), .B2(new_n210), .ZN(new_n532));
  NOR4_X1   g0332(.A1(new_n395), .A2(new_n396), .A3(new_n414), .A4(G20), .ZN(new_n533));
  OAI21_X1  g0333(.A(G107), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(KEYINPUT82), .A2(G97), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(KEYINPUT82), .A2(G97), .ZN(new_n538));
  OAI211_X1 g0338(.A(KEYINPUT6), .B(new_n368), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  XNOR2_X1  g0341(.A(G97), .B(G107), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n228), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n536), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(KEYINPUT83), .A3(KEYINPUT6), .A4(new_n368), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n210), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n268), .B1(new_n535), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n276), .A2(G97), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n516), .A2(new_n290), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n521), .A3(G190), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n523), .A2(new_n524), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(G169), .B1(new_n553), .B2(new_n521), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n521), .A2(new_n495), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n520), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n549), .A2(new_n524), .A3(new_n551), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n470), .A2(new_n378), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT86), .ZN(new_n563));
  AOI21_X1  g0363(.A(G20), .B1(new_n281), .B2(new_n282), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G87), .A2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n545), .A2(new_n536), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n210), .B1(new_n338), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(G68), .A2(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT85), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n262), .B1(new_n545), .B2(new_n536), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n316), .B1(new_n537), .B2(new_n538), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(KEYINPUT85), .A3(new_n567), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n268), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n276), .A2(new_n378), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n563), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  AOI211_X1 g0379(.A(KEYINPUT86), .B(new_n577), .C1(new_n575), .C2(new_n268), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n562), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n483), .A2(new_n224), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n296), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n296), .A2(G274), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n487), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n283), .A2(G244), .A3(G1698), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n586), .B(new_n447), .C1(new_n287), .C2(new_n222), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n587), .B2(new_n290), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(G169), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n495), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n581), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n309), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G200), .B2(new_n588), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n477), .A2(new_n223), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n595), .C1(new_n580), .C2(new_n579), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  INV_X1    g0398(.A(G116), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n469), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n330), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n272), .A2(new_n599), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT20), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(G20), .ZN(new_n605));
  AOI21_X1  g0405(.A(G33), .B1(new_n545), .B2(new_n536), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n510), .A2(new_n210), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n604), .B1(new_n608), .B2(new_n413), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n606), .A2(new_n607), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(KEYINPUT20), .A3(new_n268), .A4(new_n605), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n603), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(G303), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n296), .B1(new_n397), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(G257), .A2(G1698), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n286), .A2(G264), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n283), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n484), .A2(G270), .A3(new_n296), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n489), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G169), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n598), .B1(new_n612), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n611), .A2(new_n609), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n330), .A2(new_n600), .B1(new_n599), .B2(new_n272), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n625), .A2(KEYINPUT21), .A3(G169), .A4(new_n620), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n620), .A2(new_n495), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n622), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n620), .A2(new_n438), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n630), .B(new_n625), .C1(G200), .C2(new_n620), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n597), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n445), .A2(new_n506), .A3(new_n561), .A4(new_n632), .ZN(G372));
  NAND2_X1  g0433(.A1(new_n576), .A2(new_n578), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT86), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n576), .A2(new_n563), .A3(new_n578), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n594), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n593), .B1(new_n581), .B2(new_n590), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n496), .B1(new_n478), .B2(new_n461), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(new_n622), .A3(new_n628), .A4(new_n626), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n504), .A2(new_n471), .B1(new_n559), .B2(new_n558), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n638), .A2(new_n555), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n581), .A2(new_n643), .A3(new_n590), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n581), .B2(new_n590), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n558), .A2(new_n559), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT26), .B1(new_n638), .B2(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(KEYINPUT26), .A2(new_n591), .A3(new_n647), .A4(new_n596), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n642), .B(new_n646), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n445), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n425), .A2(new_n426), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n268), .A3(new_n429), .ZN(new_n653));
  INV_X1    g0453(.A(new_n412), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n405), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(new_n432), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n366), .A2(new_n382), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n361), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(new_n443), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n313), .A2(new_n314), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n304), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n651), .A2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n472), .A2(new_n479), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n506), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n497), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n670), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n612), .A2(new_n677), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n629), .A2(new_n631), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n629), .A2(new_n678), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n639), .A2(new_n670), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n629), .A2(new_n677), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n497), .A3(new_n505), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n213), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n566), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n216), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n644), .A2(new_n645), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT26), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n597), .B2(new_n560), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n638), .A2(KEYINPUT26), .A3(new_n647), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n626), .A2(new_n628), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n497), .A2(new_n622), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n555), .A3(new_n638), .A4(new_n641), .ZN(new_n702));
  AOI211_X1 g0502(.A(new_n694), .B(new_n670), .C1(new_n699), .C2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n702), .B(new_n646), .C1(new_n648), .C2(new_n649), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT93), .B1(new_n704), .B2(new_n677), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT29), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  INV_X1    g0507(.A(new_n650), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n670), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n588), .A2(new_n553), .A3(new_n521), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(KEYINPUT30), .A3(new_n501), .A4(new_n627), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n627), .A2(new_n501), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n588), .A2(new_n553), .A3(new_n521), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n587), .A2(new_n290), .ZN(new_n719));
  INV_X1    g0519(.A(new_n585), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(KEYINPUT92), .A3(new_n495), .A4(new_n620), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT92), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n620), .A2(new_n495), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n588), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n493), .A3(new_n522), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n711), .B(new_n677), .C1(new_n718), .C2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n717), .A3(new_n713), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT31), .B1(new_n729), .B2(new_n670), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n632), .A2(new_n506), .A3(new_n561), .A4(new_n677), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n676), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n710), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n693), .B1(new_n734), .B2(G1), .ZN(G364));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n679), .A2(new_n680), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n271), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n209), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n688), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n218), .B1(G20), .B2(new_n301), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n210), .A2(new_n495), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n438), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n305), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n270), .A2(new_n750), .B1(new_n753), .B2(new_n285), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n305), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G20), .A3(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n223), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n210), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n755), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n368), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n754), .A2(new_n397), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n751), .A2(new_n438), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G58), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n748), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n210), .B1(new_n767), .B2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(G68), .B1(G97), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n758), .A2(new_n767), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G159), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT32), .Z(new_n774));
  NAND4_X1  g0574(.A1(new_n761), .A2(new_n765), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n756), .A2(new_n613), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n397), .B1(new_n759), .B2(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n776), .B(new_n778), .C1(G329), .C2(new_n772), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n762), .A2(G322), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n766), .A2(new_n781), .B1(new_n752), .B2(G311), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n749), .A2(G326), .B1(G294), .B2(new_n769), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n779), .A2(new_n780), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n746), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n738), .A2(new_n745), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n213), .A2(new_n283), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(G116), .B2(new_n213), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n687), .A2(new_n283), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n216), .B2(G45), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(G45), .B2(new_n250), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n744), .B(new_n785), .C1(new_n786), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n739), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT96), .Z(new_n797));
  AND3_X1   g0597(.A1(new_n679), .A2(new_n676), .A3(new_n680), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n681), .B(new_n798), .C1(new_n689), .C2(new_n741), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  OAI21_X1  g0601(.A(new_n385), .B1(new_n381), .B2(new_n677), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n383), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n382), .A2(new_n677), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n650), .B2(new_n677), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT99), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n386), .A2(new_n670), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n650), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n650), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(KEYINPUT99), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n806), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(new_n733), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n733), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n688), .C2(new_n742), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n745), .A2(new_n736), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT97), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n744), .B1(new_n818), .B2(new_n285), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G294), .A2(new_n762), .B1(new_n752), .B2(G116), .ZN(new_n820));
  INV_X1    g0620(.A(new_n766), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n777), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n397), .B1(new_n771), .B2(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n756), .A2(new_n368), .B1(new_n759), .B2(new_n223), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n750), .A2(new_n613), .B1(new_n228), .B2(new_n768), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n756), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n397), .B1(new_n828), .B2(G50), .ZN(new_n829));
  INV_X1    g0629(.A(new_n759), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G68), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n829), .B(new_n831), .C1(new_n832), .C2(new_n771), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G58), .B2(new_n769), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT98), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G137), .A2(new_n749), .B1(new_n752), .B2(G159), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n253), .B2(new_n821), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G143), .B2(new_n764), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n827), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n819), .B1(new_n842), .B2(new_n746), .C1(new_n805), .C2(new_n737), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n815), .A2(new_n843), .ZN(G384));
  AND2_X1   g0644(.A1(new_n543), .A2(new_n547), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT35), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT35), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(G116), .A3(new_n219), .A4(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT36), .Z(new_n850));
  OAI211_X1 g0650(.A(new_n217), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n270), .A2(G68), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n209), .B(G13), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n668), .B(KEYINPUT102), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n657), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n408), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT37), .B1(new_n860), .B2(new_n655), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n653), .A2(new_n654), .A3(new_n440), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n855), .B1(new_n653), .B2(new_n654), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT103), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT103), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n409), .B2(new_n430), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n653), .A2(new_n654), .A3(new_n440), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n430), .B2(new_n855), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n652), .A2(new_n269), .A3(new_n429), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n654), .ZN(new_n874));
  INV_X1    g0674(.A(new_n668), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n869), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n874), .A2(new_n405), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT101), .B(KEYINPUT37), .C1(new_n877), .C2(new_n878), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n872), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n876), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n433), .B2(new_n443), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT38), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n867), .B1(new_n864), .B2(new_n656), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n871), .B2(new_n865), .ZN(new_n889));
  INV_X1    g0689(.A(new_n863), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n441), .B(KEYINPUT17), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n657), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n887), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT39), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n883), .B2(new_n885), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n894), .B1(new_n897), .B2(KEYINPUT39), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n361), .A2(new_n670), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n857), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n333), .A2(new_n670), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n361), .A2(new_n366), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n333), .B(new_n670), .C1(new_n357), .C2(new_n360), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n650), .A2(new_n807), .A3(new_n808), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n807), .B1(new_n650), .B2(new_n808), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n804), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT100), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(KEYINPUT100), .B(new_n804), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n895), .B2(new_n896), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n900), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n706), .A2(new_n445), .A3(new_n709), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n663), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n914), .B(new_n916), .Z(new_n917));
  NOR3_X1   g0717(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT40), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n731), .A2(new_n732), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n904), .A3(new_n805), .ZN(new_n920));
  AND2_X1   g0720(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n886), .A2(new_n893), .B1(new_n920), .B2(KEYINPUT104), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n918), .A2(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n445), .A3(new_n919), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n886), .A2(new_n893), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n920), .A2(KEYINPUT104), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n883), .A2(new_n885), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n887), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n925), .A3(new_n886), .ZN(new_n933));
  AOI22_X1  g0733(.A1(KEYINPUT40), .A2(new_n930), .B1(new_n933), .B2(new_n922), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n445), .A2(new_n919), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n927), .A2(new_n936), .A3(G330), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n917), .A2(new_n937), .B1(new_n209), .B2(new_n740), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n917), .A2(new_n937), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n854), .B1(new_n941), .B2(new_n942), .ZN(G367));
  NOR2_X1   g0743(.A1(new_n637), .A2(new_n677), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n597), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n695), .B2(new_n944), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n738), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n239), .A2(new_n687), .A3(new_n283), .ZN(new_n948));
  INV_X1    g0748(.A(new_n378), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n786), .B1(new_n213), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n743), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n756), .A2(new_n202), .B1(new_n759), .B2(new_n285), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n397), .B(new_n952), .C1(G137), .C2(new_n772), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n752), .A2(G50), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n762), .A2(G150), .B1(G68), .B2(new_n769), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G143), .A2(new_n749), .B1(new_n766), .B2(G159), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n777), .A2(new_n753), .B1(new_n750), .B2(new_n823), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G107), .B2(new_n769), .ZN(new_n959));
  INV_X1    g0759(.A(G317), .ZN(new_n960));
  INV_X1    g0760(.A(new_n546), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n397), .B1(new_n771), .B2(new_n960), .C1(new_n961), .C2(new_n759), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n959), .B(new_n963), .C1(new_n613), .C2(new_n763), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n828), .A2(KEYINPUT46), .A3(G116), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT46), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n756), .B2(new_n599), .ZN(new_n967));
  INV_X1    g0767(.A(G294), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n965), .B(new_n967), .C1(new_n821), .C2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT109), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n957), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n951), .B1(new_n972), .B2(new_n745), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n947), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n682), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n559), .A2(new_n670), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n555), .A2(new_n560), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n647), .A2(new_n670), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT106), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT108), .ZN(new_n983));
  INV_X1    g0783(.A(new_n685), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT107), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n985), .A3(new_n979), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n977), .A2(new_n978), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT107), .B1(new_n987), .B2(new_n685), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT42), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n985), .B1(new_n984), .B2(new_n979), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n987), .A2(new_n685), .A3(KEYINPUT107), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT42), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n647), .B1(new_n981), .B2(new_n673), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n990), .B(new_n993), .C1(new_n994), .C2(new_n670), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n995), .A2(new_n996), .A3(new_n946), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n946), .A2(new_n996), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n946), .A2(new_n996), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n999), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n983), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n995), .A2(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n998), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT108), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n982), .B(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n995), .A2(new_n996), .A3(new_n946), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n733), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n706), .A2(new_n709), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n685), .A2(new_n683), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n987), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT44), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(KEYINPUT44), .A3(new_n987), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1013), .B2(new_n987), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n685), .A2(new_n979), .A3(KEYINPUT45), .A4(new_n683), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n975), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1016), .A2(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n682), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n685), .B1(new_n675), .B2(new_n684), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1028), .A2(new_n681), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(new_n681), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1011), .B(new_n1012), .C1(new_n1027), .C2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n688), .B(KEYINPUT41), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n742), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n974), .B1(new_n1010), .B2(new_n1035), .ZN(G387));
  OR2_X1    g0836(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n734), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT111), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1012), .A2(new_n1037), .A3(new_n1011), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n688), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1039), .A3(new_n688), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n672), .A2(new_n674), .A3(new_n738), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n791), .B1(new_n243), .B2(new_n341), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n690), .B2(new_n787), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n261), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1048));
  AOI21_X1  g0848(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT50), .B1(new_n261), .B2(G50), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1048), .A2(new_n690), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1047), .A2(new_n1051), .B1(new_n368), .B2(new_n687), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n786), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n743), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G50), .A2(new_n762), .B1(new_n752), .B2(G68), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n261), .B2(new_n821), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n397), .B1(new_n830), .B2(G97), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n828), .A2(G77), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n253), .C2(new_n771), .ZN(new_n1059));
  INV_X1    g0859(.A(G159), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n750), .A2(new_n1060), .B1(new_n949), .B2(new_n768), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1056), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT110), .Z(new_n1063));
  AOI22_X1  g0863(.A1(G303), .A2(new_n752), .B1(new_n766), .B2(G311), .ZN(new_n1064));
  INV_X1    g0864(.A(G322), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n750), .C1(new_n763), .C2(new_n960), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n756), .A2(new_n968), .B1(new_n768), .B2(new_n777), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(KEYINPUT49), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n283), .B1(new_n772), .B2(G326), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n599), .C2(new_n759), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT49), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1054), .B1(new_n1075), .B2(new_n745), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1037), .A2(new_n742), .B1(new_n1045), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1044), .A2(new_n1077), .ZN(G393));
  OAI21_X1  g0878(.A(KEYINPUT112), .B1(new_n1025), .B2(new_n682), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1018), .A2(new_n682), .A3(new_n1022), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1023), .A2(KEYINPUT112), .A3(new_n975), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n742), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n786), .B1(new_n213), .B2(new_n961), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n791), .B2(new_n247), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n744), .A2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G294), .A2(new_n752), .B1(new_n766), .B2(G303), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n599), .B2(new_n768), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n756), .A2(new_n777), .B1(new_n771), .B2(new_n1065), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1088), .A2(new_n283), .A3(new_n760), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G311), .A2(new_n762), .B1(new_n749), .B2(G317), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT52), .Z(new_n1092));
  AOI22_X1  g0892(.A1(G150), .A2(new_n749), .B1(new_n762), .B2(G159), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT51), .Z(new_n1094));
  AOI21_X1  g0894(.A(new_n397), .B1(new_n830), .B2(G87), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G50), .A2(new_n766), .B1(new_n752), .B2(new_n260), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n828), .A2(G68), .B1(new_n772), .B2(G143), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n769), .A2(G77), .ZN(new_n1098));
  AND4_X1   g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1090), .A2(new_n1092), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n738), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1086), .B1(new_n746), .B2(new_n1100), .C1(new_n981), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1082), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1024), .A2(KEYINPUT112), .A3(new_n1026), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1040), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n688), .B1(new_n1040), .B2(new_n1027), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1083), .B(new_n1102), .C1(new_n1106), .C2(new_n1107), .ZN(G390));
  NAND2_X1  g0908(.A1(new_n445), .A2(new_n733), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n915), .A2(new_n663), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n733), .A2(new_n805), .A3(new_n904), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT113), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n904), .B1(new_n733), .B2(new_n805), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n811), .A2(new_n809), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT100), .B1(new_n1114), .B2(new_n804), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n911), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1112), .A2(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n705), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n704), .A2(KEYINPUT93), .A3(new_n677), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n1119), .A3(new_n804), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n803), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1113), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1111), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1110), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n932), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n928), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(KEYINPUT39), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n912), .B2(new_n899), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n899), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1130), .B(new_n928), .C1(new_n1121), .C2(new_n905), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1129), .A2(new_n1131), .A3(new_n1111), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1112), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1125), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1131), .A3(new_n1111), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n928), .A2(new_n1130), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n803), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n703), .A2(new_n705), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n804), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1137), .B1(new_n1140), .B2(new_n904), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n904), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1130), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1141), .B1(new_n1143), .B2(new_n1128), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1136), .B(new_n1124), .C1(new_n1144), .C2(new_n1133), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1135), .A2(new_n688), .A3(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G283), .A2(new_n749), .B1(new_n766), .B2(G107), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n961), .B2(new_n753), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n757), .A2(new_n283), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1149), .B(new_n831), .C1(new_n968), .C2(new_n771), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n762), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1098), .B1(new_n1151), .B2(new_n599), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1148), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n828), .A2(G150), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  INV_X1    g0955(.A(G128), .ZN(new_n1156));
  INV_X1    g0956(.A(G137), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1156), .A2(new_n750), .B1(new_n821), .B2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n753), .A2(new_n1159), .B1(new_n1060), .B2(new_n768), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n772), .A2(G125), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1151), .B2(new_n832), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1155), .A2(new_n1158), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n283), .B1(new_n759), .B2(new_n270), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT114), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1153), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n743), .B1(new_n260), .B2(new_n817), .C1(new_n1166), .C2(new_n746), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1128), .B2(new_n736), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1169), .B2(new_n742), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1146), .A2(new_n1170), .A3(KEYINPUT115), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT115), .B1(new_n1146), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(G378));
  NAND2_X1  g0973(.A1(new_n279), .A2(new_n875), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n315), .B(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1175), .B(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n926), .A2(G330), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n926), .B2(G330), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n914), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1178), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n934), .B2(new_n676), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n926), .A2(G330), .A3(new_n1178), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1183), .A2(new_n913), .A3(new_n900), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n742), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n736), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n743), .B1(new_n817), .B2(G50), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G125), .A2(new_n749), .B1(new_n766), .B2(G132), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n1156), .B2(new_n1151), .C1(new_n1157), .C2(new_n753), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n756), .A2(new_n1159), .B1(new_n768), .B2(new_n253), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n255), .B(new_n295), .C1(new_n759), .C2(new_n1060), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G124), .B2(new_n772), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n599), .A2(new_n750), .B1(new_n753), .B2(new_n949), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n759), .A2(new_n202), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G283), .B2(new_n772), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n766), .A2(G97), .B1(G68), .B2(new_n769), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n283), .A2(G41), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1058), .A4(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1200), .B(new_n1205), .C1(G107), .C2(new_n762), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1204), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n270), .C1(G33), .C2(G41), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1199), .A2(new_n1207), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1189), .B1(new_n1211), .B2(new_n745), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1188), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT116), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1187), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1110), .B(KEYINPUT117), .Z(new_n1217));
  NAND2_X1  g1017(.A1(new_n1145), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n688), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1218), .B2(new_n1186), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1216), .B1(new_n1222), .B2(new_n1223), .ZN(G375));
  OAI22_X1  g1024(.A1(new_n821), .A2(new_n599), .B1(new_n753), .B2(new_n368), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G283), .B2(new_n762), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n756), .A2(new_n228), .B1(new_n771), .B2(new_n613), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n283), .B(new_n1227), .C1(G77), .C2(new_n830), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n749), .A2(G294), .B1(new_n378), .B2(new_n769), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n749), .A2(G132), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT118), .Z(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n1157), .B2(new_n763), .C1(new_n821), .C2(new_n1159), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT119), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n753), .A2(new_n253), .B1(new_n270), .B2(new_n768), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n756), .A2(new_n1060), .B1(new_n771), .B2(new_n1156), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n397), .A4(new_n1201), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1230), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n745), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n744), .B1(new_n818), .B2(new_n203), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n904), .C2(new_n737), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1117), .A2(new_n1123), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n741), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT120), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(KEYINPUT120), .B(new_n1243), .C1(new_n1244), .C2(new_n741), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1110), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1034), .A3(new_n1125), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(G381));
  NAND2_X1  g1052(.A1(new_n1218), .A2(new_n1186), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1219), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n689), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1215), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT121), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1146), .A2(new_n1170), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  OR3_X1    g1059(.A1(G387), .A2(G390), .A3(G384), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1044), .A2(new_n800), .A3(new_n1077), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(G381), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1257), .A2(new_n1259), .A3(new_n1262), .ZN(G407));
  NAND2_X1  g1063(.A1(new_n669), .A2(G213), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT122), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1257), .A2(new_n1259), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(G407), .A2(new_n1266), .A3(G213), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT123), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1267), .B(new_n1268), .ZN(G409));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1250), .B1(new_n1270), .B2(new_n1124), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1244), .A2(KEYINPUT60), .A3(new_n1110), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n688), .A3(new_n1272), .ZN(new_n1273));
  XOR2_X1   g1073(.A(G384), .B(KEYINPUT124), .Z(new_n1274));
  AND3_X1   g1074(.A1(new_n1273), .A2(new_n1249), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT124), .B1(new_n815), .B2(new_n843), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1273), .B2(new_n1249), .ZN(new_n1277));
  INV_X1    g1077(.A(G2897), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1265), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n1275), .A2(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1273), .A2(new_n1249), .A3(new_n1274), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1264), .A2(new_n1278), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1273), .A2(new_n1249), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1281), .B(new_n1282), .C1(new_n1283), .C2(new_n1276), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1145), .A2(new_n1217), .B1(new_n1185), .B2(new_n1181), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1034), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1186), .A2(new_n742), .B1(new_n1188), .B2(new_n1212), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1258), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(G378), .B2(new_n1256), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1264), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1285), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1259), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT115), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1135), .A2(new_n688), .A3(new_n1145), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1168), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1136), .B1(new_n1144), .B2(new_n1133), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1298), .B2(new_n741), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1295), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1146), .A2(new_n1170), .A3(KEYINPUT115), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1294), .B1(new_n1302), .B2(G375), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1275), .A2(new_n1277), .A3(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1279), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT125), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1035), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1310), .B2(new_n974), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1083), .A2(new_n1102), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1107), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1313), .B2(new_n1105), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(G387), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1307), .B1(new_n1311), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1043), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1317), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1077), .ZN(new_n1319));
  OAI21_X1  g1119(.A(G396), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1320), .A2(new_n1261), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1316), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1310), .A2(new_n974), .A3(G390), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G387), .A2(new_n1314), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1320), .A2(new_n1261), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(new_n1327), .A3(new_n1307), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1322), .A2(new_n1323), .A3(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT126), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1322), .A2(new_n1328), .A3(KEYINPUT126), .A4(new_n1323), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1292), .A2(new_n1306), .A3(new_n1333), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1221), .B(new_n688), .C1(KEYINPUT57), .C2(new_n1286), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1335), .A2(new_n1300), .A3(new_n1301), .A4(new_n1216), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1291), .B1(new_n1336), .B2(new_n1294), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT63), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(KEYINPUT127), .B1(new_n1334), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1303), .A2(new_n1264), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1265), .B1(new_n1336), .B2(new_n1294), .ZN(new_n1342));
  AOI22_X1  g1142(.A1(new_n1341), .A2(new_n1285), .B1(new_n1342), .B2(new_n1305), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT127), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1303), .A2(new_n1264), .A3(new_n1338), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1304), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1343), .A2(new_n1344), .A3(new_n1346), .A4(new_n1333), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1340), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1322), .A2(new_n1328), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT62), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1275), .A2(new_n1277), .A3(new_n1350), .ZN(new_n1351));
  AOI22_X1  g1151(.A1(new_n1345), .A2(new_n1350), .B1(new_n1342), .B2(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1285), .B1(new_n1290), .B2(new_n1265), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1323), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1349), .B1(new_n1352), .B2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1348), .A2(new_n1355), .ZN(G405));
  XNOR2_X1  g1156(.A(new_n1349), .B(new_n1338), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1336), .B1(new_n1258), .B2(new_n1256), .ZN(new_n1358));
  XNOR2_X1  g1158(.A(new_n1357), .B(new_n1358), .ZN(G402));
endmodule


