//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT86), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G214), .A3(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT86), .B(G143), .ZN(new_n192));
  INV_X1    g006(.A(G214), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n193), .A2(G237), .A3(G953), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  OR2_X1    g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT88), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(G131), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n195), .B2(G131), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n187), .B(new_n196), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n200), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT17), .A3(new_n198), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(KEYINPUT72), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT72), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(G125), .A3(G140), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT73), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(G125), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT16), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n210), .B1(new_n206), .B2(new_n208), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(G146), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n216), .A3(G146), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n201), .A2(new_n203), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G113), .B(G122), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n195), .A2(G131), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n191), .B(new_n225), .C1(new_n192), .C2(new_n194), .ZN(new_n227));
  XNOR2_X1  g041(.A(G125), .B(G140), .ZN(new_n228));
  MUX2_X1   g042(.A(new_n228), .B(new_n209), .S(G146), .Z(new_n229));
  NAND4_X1  g043(.A1(new_n226), .A2(new_n227), .A3(new_n229), .A4(new_n196), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n220), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n196), .B1(new_n199), .B2(new_n200), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT74), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n219), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n211), .A2(new_n216), .A3(KEYINPUT74), .A4(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n209), .A2(KEYINPUT19), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT19), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n228), .A2(KEYINPUT89), .A3(new_n237), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(new_n240), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n232), .A2(new_n234), .A3(new_n235), .A4(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n230), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT90), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n223), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n230), .A3(KEYINPUT90), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n231), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(G475), .A2(G902), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT20), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT20), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n244), .A2(KEYINPUT90), .A3(new_n230), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT90), .B1(new_n244), .B2(new_n230), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n254), .A2(new_n255), .A3(new_n223), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n253), .B(new_n250), .C1(new_n256), .C2(new_n231), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G475), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n220), .A2(new_n230), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT91), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n223), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(G902), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n260), .B1(new_n262), .B2(new_n223), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(G234), .A2(G237), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(G952), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT21), .B(G898), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT94), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n269), .A2(G902), .A3(G953), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT92), .ZN(new_n278));
  INV_X1    g092(.A(G128), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(G143), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n188), .A2(KEYINPUT92), .A3(G128), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(G143), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G134), .ZN(new_n285));
  INV_X1    g099(.A(G134), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n282), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G107), .ZN(new_n289));
  INV_X1    g103(.A(G122), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G116), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n291), .B2(KEYINPUT14), .ZN(new_n292));
  INV_X1    g106(.A(G116), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G122), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n295), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n288), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT13), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n282), .A2(new_n299), .B1(new_n279), .B2(G143), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n280), .A2(KEYINPUT13), .A3(new_n281), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n286), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n291), .A2(new_n294), .A3(G107), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n295), .A2(new_n289), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n287), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT93), .B1(new_n298), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n302), .A2(new_n305), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT93), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n288), .A2(new_n296), .A3(new_n297), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  INV_X1    g126(.A(G217), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n312), .A2(new_n313), .A3(G953), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n307), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n307), .B2(new_n311), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n277), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G478), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT15), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n318), .B(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n268), .A2(new_n276), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(new_n222), .B2(G107), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n289), .A3(G104), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n222), .A2(G107), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G101), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n325), .A3(new_n329), .A4(new_n326), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT64), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n293), .B2(G119), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT64), .A3(G116), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n293), .A2(G119), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G113), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT2), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G113), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n341), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n343), .A2(new_n333), .A3(new_n335), .A4(new_n336), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n327), .A2(new_n346), .A3(G101), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n331), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G110), .B(G122), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n293), .A2(G119), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT5), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n338), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n337), .B2(new_n353), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n344), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n222), .A2(G107), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n289), .A2(G104), .ZN(new_n358));
  OAI21_X1  g172(.A(G101), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n330), .A2(new_n359), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n331), .A2(new_n345), .A3(KEYINPUT82), .A4(new_n347), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n350), .A2(new_n351), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(KEYINPUT83), .A2(KEYINPUT6), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n351), .ZN(new_n366));
  INV_X1    g180(.A(new_n350), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n362), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n366), .B(new_n364), .C1(new_n367), .C2(new_n368), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n241), .A2(G143), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n188), .A2(G146), .ZN(new_n374));
  AND2_X1   g188(.A1(KEYINPUT0), .A2(G128), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G143), .B(G146), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT0), .B(G128), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G125), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n379), .B2(G125), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n188), .A2(G146), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n241), .A2(G143), .ZN(new_n387));
  OAI211_X1 g201(.A(G128), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n373), .B(new_n374), .C1(KEYINPUT1), .C2(new_n279), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n205), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n270), .A2(G224), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n372), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n356), .B(new_n360), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n351), .B(KEYINPUT8), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n379), .A2(G125), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT84), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT85), .A3(new_n381), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n403));
  AND4_X1   g217(.A1(new_n384), .A2(new_n402), .A3(new_n391), .A4(new_n403), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n403), .A2(new_n402), .B1(new_n384), .B2(new_n391), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n363), .B(new_n399), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n277), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n409), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n394), .B1(new_n370), .B2(new_n371), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(new_n407), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G214), .B1(G237), .B2(G902), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n270), .A2(G227), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND4_X1  g233(.A1(new_n388), .A2(new_n330), .A3(new_n359), .A4(new_n389), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT10), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT11), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n286), .B2(G137), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n286), .A2(G137), .ZN(new_n424));
  INV_X1    g238(.A(G137), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT11), .A3(G134), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G131), .ZN(new_n428));
  INV_X1    g242(.A(G131), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n423), .A2(new_n426), .A3(new_n429), .A4(new_n424), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT78), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n433));
  INV_X1    g247(.A(new_n379), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(new_n347), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n435), .B2(new_n331), .ZN(new_n436));
  AND4_X1   g250(.A1(new_n433), .A2(new_n331), .A3(new_n434), .A4(new_n347), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n421), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n439));
  INV_X1    g253(.A(new_n420), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n389), .A2(new_n388), .B1(new_n330), .B2(new_n359), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n431), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT79), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT12), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI221_X1 g259(.A(new_n431), .B1(new_n443), .B2(KEYINPUT12), .C1(new_n440), .C2(new_n441), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n438), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n439), .B1(new_n438), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n419), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n421), .B1(new_n436), .B2(new_n437), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n431), .ZN(new_n452));
  INV_X1    g266(.A(new_n419), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n438), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(G469), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G469), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n438), .A2(new_n453), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n445), .B2(new_n446), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n445), .A2(new_n458), .A3(new_n446), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n453), .B1(new_n452), .B2(new_n438), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n456), .B(new_n277), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(G469), .A2(G902), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G221), .B1(new_n312), .B2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n416), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n322), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n313), .B1(G234), .B2(new_n277), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT23), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n334), .B2(G128), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n279), .A2(KEYINPUT23), .A3(G119), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n472), .B(new_n473), .C1(G119), .C2(new_n279), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n474), .A2(G110), .ZN(new_n475));
  XOR2_X1   g289(.A(G119), .B(G128), .Z(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT24), .B(G110), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n475), .A2(new_n478), .B1(new_n241), .B2(new_n228), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n234), .A2(new_n235), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n476), .A2(new_n477), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n474), .A2(G110), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT71), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n474), .A2(KEYINPUT71), .A3(G110), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n211), .A2(new_n216), .A3(G146), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n217), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT22), .B(G137), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT75), .Z(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(KEYINPUT76), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n480), .A2(new_n488), .A3(new_n492), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT76), .B1(new_n489), .B2(new_n493), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT25), .B1(new_n498), .B2(new_n277), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n489), .A2(new_n493), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT76), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n502), .A2(new_n277), .A3(new_n495), .A4(new_n494), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT25), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n470), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n470), .A2(G902), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n424), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n286), .A2(G137), .ZN(new_n511));
  OAI21_X1  g325(.A(G131), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n512), .A2(new_n388), .A3(new_n389), .A4(new_n430), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n431), .A2(KEYINPUT65), .A3(new_n434), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT65), .B1(new_n431), .B2(new_n434), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT30), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n342), .A2(new_n344), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n431), .A2(new_n434), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n513), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n513), .B(new_n517), .C1(new_n514), .C2(new_n515), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n190), .A2(G210), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n524), .B(KEYINPUT67), .Z(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT26), .B(G101), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n525), .B(new_n528), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT68), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n516), .A2(new_n521), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n523), .A4(new_n529), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(KEYINPUT31), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT65), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n518), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n431), .A2(KEYINPUT65), .A3(new_n434), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(KEYINPUT28), .A3(new_n513), .A4(new_n517), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n517), .B1(new_n518), .B2(new_n513), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n518), .A2(new_n517), .A3(new_n513), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n529), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n530), .B1(new_n516), .B2(new_n521), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT31), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n535), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(G472), .A2(G902), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT69), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n553));
  INV_X1    g367(.A(new_n550), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n535), .B2(new_n548), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT69), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n552), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n517), .B1(new_n539), .B2(new_n513), .ZN(new_n559));
  INV_X1    g373(.A(new_n523), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT28), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n543), .A2(new_n542), .ZN(new_n562));
  INV_X1    g376(.A(new_n529), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT29), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT70), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n532), .A2(new_n523), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n563), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n540), .A2(new_n544), .A3(new_n529), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT70), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n561), .A2(new_n572), .A3(new_n562), .A4(new_n565), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n567), .A2(new_n277), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n574), .A2(G472), .B1(new_n555), .B2(KEYINPUT32), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n509), .B1(new_n558), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n469), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT95), .B(G101), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G3));
  NAND2_X1  g393(.A1(new_n549), .A2(new_n277), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n552), .A2(new_n581), .A3(new_n557), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n582), .A2(new_n509), .A3(new_n467), .ZN(new_n583));
  INV_X1    g397(.A(new_n276), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n409), .B1(new_n396), .B2(new_n408), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n412), .A2(new_n407), .A3(new_n411), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n415), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n266), .B1(new_n252), .B2(new_n257), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n316), .B2(new_n317), .ZN(new_n590));
  INV_X1    g404(.A(new_n317), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT33), .A3(new_n315), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n590), .A2(new_n592), .A3(G478), .A4(new_n277), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n318), .A2(new_n319), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n587), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n583), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT34), .B(G104), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G6));
  NAND2_X1  g413(.A1(new_n588), .A2(new_n321), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT96), .B1(new_n600), .B2(new_n587), .ZN(new_n601));
  INV_X1    g415(.A(new_n415), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n602), .B(new_n276), .C1(new_n410), .C2(new_n413), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n321), .A4(new_n588), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n583), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G107), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  INV_X1    g422(.A(new_n470), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n498), .A2(KEYINPUT25), .A3(new_n277), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n503), .A2(new_n504), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n489), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n507), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n582), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n469), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT37), .B(G110), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G12));
  AOI21_X1  g435(.A(new_n617), .B1(new_n558), .B2(new_n575), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n270), .A2(G900), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(G902), .A3(new_n269), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n271), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n588), .A2(new_n321), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n588), .A2(KEYINPUT98), .A3(new_n321), .A4(new_n628), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n622), .A2(new_n468), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT99), .B(G128), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G30));
  AND2_X1   g449(.A1(new_n465), .A2(new_n466), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n628), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT40), .Z(new_n640));
  AND2_X1   g454(.A1(new_n531), .A2(new_n534), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n345), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n529), .B1(new_n643), .B2(new_n523), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n277), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n648), .A2(G472), .B1(KEYINPUT32), .B2(new_n555), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n558), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n585), .A2(new_n586), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT38), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n617), .A2(new_n415), .ZN(new_n653));
  INV_X1    g467(.A(new_n320), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n318), .B(new_n654), .ZN(new_n655));
  NOR4_X1   g469(.A1(new_n652), .A2(new_n653), .A3(new_n655), .A4(new_n588), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n640), .A2(new_n650), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  INV_X1    g472(.A(new_n628), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n588), .A2(new_n595), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n622), .A2(new_n468), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT102), .B(G146), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G48));
  NAND2_X1  g477(.A1(new_n558), .A2(new_n575), .ZN(new_n664));
  INV_X1    g478(.A(new_n509), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n461), .A2(new_n462), .ZN(new_n666));
  OAI21_X1  g480(.A(G469), .B1(new_n666), .B2(G902), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n466), .A3(new_n463), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n664), .A2(new_n596), .A3(new_n665), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT41), .B(G113), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G15));
  NAND4_X1  g486(.A1(new_n576), .A2(new_n605), .A3(new_n601), .A4(new_n669), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G116), .ZN(G18));
  NAND2_X1  g488(.A1(new_n506), .A2(new_n615), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n416), .A2(new_n668), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n664), .A2(new_n322), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  NOR3_X1   g492(.A1(new_n416), .A2(new_n655), .A3(new_n588), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT103), .B1(new_n561), .B2(new_n562), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n542), .B1(new_n643), .B2(new_n523), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n682));
  INV_X1    g496(.A(new_n562), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n680), .A2(new_n684), .A3(new_n529), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n546), .A2(new_n547), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n535), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n550), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n688), .A2(new_n581), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n668), .A2(new_n276), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n679), .A2(new_n665), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  AND4_X1   g506(.A1(new_n675), .A2(new_n660), .A3(new_n676), .A4(new_n689), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n205), .ZN(G27));
  NAND3_X1  g508(.A1(new_n551), .A2(KEYINPUT104), .A3(new_n553), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n555), .B2(KEYINPUT32), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n575), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n410), .A2(new_n413), .A3(new_n415), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n467), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n660), .A2(new_n698), .A3(new_n700), .A4(new_n665), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT42), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n593), .A2(new_n594), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n268), .A2(new_n703), .A3(new_n628), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n651), .A2(new_n415), .A3(new_n466), .A4(new_n465), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n576), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n429), .ZN(G33));
  AND3_X1   g524(.A1(new_n664), .A2(new_n665), .A3(new_n700), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n631), .A2(new_n632), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G134), .ZN(G36));
  XNOR2_X1  g529(.A(new_n268), .B(KEYINPUT105), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n595), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n717), .B1(new_n268), .B2(new_n595), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n582), .A3(new_n675), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT44), .ZN(new_n723));
  INV_X1    g537(.A(new_n699), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT45), .B1(new_n450), .B2(new_n454), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n456), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n450), .A2(KEYINPUT45), .A3(new_n454), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT46), .B1(new_n728), .B2(new_n464), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n452), .A2(new_n438), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n419), .ZN(new_n731));
  INV_X1    g545(.A(new_n459), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n445), .A2(new_n446), .A3(new_n458), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n453), .A3(new_n438), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(G902), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n729), .B1(new_n456), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n464), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n466), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(new_n638), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n723), .A2(new_n724), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G137), .ZN(G39));
  NAND2_X1  g557(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n664), .A2(new_n665), .A3(new_n699), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n660), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G140), .ZN(G42));
  NOR3_X1   g564(.A1(new_n668), .A2(new_n271), .A3(new_n699), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n721), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n698), .A2(new_n665), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT48), .ZN(new_n756));
  INV_X1    g570(.A(new_n650), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n665), .A3(new_n751), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n268), .A2(new_n703), .ZN(new_n759));
  OAI211_X1 g573(.A(G952), .B(new_n270), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n665), .A2(new_n689), .A3(new_n272), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n719), .B2(new_n720), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n760), .B1(new_n676), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n758), .A2(new_n268), .A3(new_n703), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n602), .A3(new_n652), .A4(new_n669), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT50), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n688), .B(new_n581), .C1(new_n612), .C2(new_n616), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n765), .B(new_n767), .C1(new_n769), .C2(new_n752), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n735), .B(G469), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n744), .B(new_n746), .C1(new_n466), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n724), .A3(new_n762), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n764), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n622), .A2(new_n468), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n693), .B1(new_n778), .B2(new_n713), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n636), .A2(new_n617), .A3(KEYINPUT110), .A4(new_n628), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n465), .A2(new_n466), .A3(new_n628), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n675), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(new_n784), .A3(new_n650), .A4(new_n679), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(new_n780), .A3(new_n661), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n693), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n633), .A3(new_n785), .A4(new_n661), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n768), .A2(new_n704), .A3(new_n705), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n711), .B2(new_n713), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n555), .A2(new_n556), .ZN(new_n794));
  AOI211_X1 g608(.A(KEYINPUT69), .B(new_n554), .C1(new_n535), .C2(new_n548), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT32), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n574), .A2(G472), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n553), .B2(new_n551), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n675), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n258), .A2(new_n655), .A3(new_n267), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n636), .A3(new_n628), .A4(new_n724), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT108), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n268), .A2(new_n321), .A3(new_n659), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n622), .A2(new_n803), .A3(new_n700), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n791), .B1(new_n793), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n793), .A2(new_n806), .A3(new_n791), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n670), .A2(new_n677), .A3(new_n691), .ZN(new_n811));
  AOI211_X1 g625(.A(KEYINPUT42), .B(new_n509), .C1(new_n558), .C2(new_n575), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n812), .A2(new_n706), .B1(new_n701), .B2(KEYINPUT42), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n813), .A3(new_n673), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n759), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n583), .A3(new_n603), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n583), .A2(new_n321), .A3(new_n588), .A4(new_n603), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n469), .B1(new_n618), .B2(new_n576), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n790), .A2(new_n810), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n822), .A2(KEYINPUT112), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT112), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n824), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT54), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n673), .A2(new_n670), .A3(new_n677), .A4(new_n691), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n709), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n811), .A2(new_n813), .A3(KEYINPUT113), .A4(new_n673), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n817), .A2(new_n819), .A3(KEYINPUT53), .A4(new_n818), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n793), .A2(new_n806), .A3(new_n791), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n789), .B(new_n786), .C1(new_n838), .C2(new_n807), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT114), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n835), .B1(new_n832), .B2(new_n833), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n790), .A2(new_n841), .A3(new_n810), .A4(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n814), .A2(new_n820), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n823), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n840), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n762), .A2(new_n724), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n773), .B2(KEYINPUT116), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(KEYINPUT116), .B2(new_n773), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n770), .A2(KEYINPUT51), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n777), .A2(new_n829), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(G952), .B2(G953), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n772), .A2(KEYINPUT49), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT106), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(KEYINPUT106), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n703), .A2(new_n415), .A3(new_n466), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n772), .B2(KEYINPUT49), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n665), .A3(new_n652), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n757), .A2(new_n716), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n853), .B1(new_n861), .B2(new_n862), .ZN(G75));
  NOR2_X1   g677(.A1(new_n270), .A2(G952), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT119), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n840), .A2(new_n843), .A3(new_n845), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(KEYINPUT118), .A3(G902), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT118), .B1(new_n866), .B2(G902), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n868), .A2(new_n869), .A3(new_n409), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n372), .A2(new_n395), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n412), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT55), .Z(new_n873));
  OR2_X1    g687(.A1(new_n873), .A2(KEYINPUT56), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n865), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT56), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n866), .A2(G902), .ZN(new_n877));
  INV_X1    g691(.A(G210), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n873), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(KEYINPUT117), .A3(new_n873), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(G51));
  INV_X1    g698(.A(new_n864), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n868), .A2(new_n869), .A3(new_n728), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n666), .B(KEYINPUT120), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n847), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n464), .B(KEYINPUT57), .Z(new_n890));
  AOI21_X1  g704(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n885), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(KEYINPUT121), .B(new_n885), .C1(new_n886), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(G54));
  INV_X1    g710(.A(new_n869), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(new_n867), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n898), .A2(new_n249), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n249), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n864), .ZN(G60));
  AND2_X1   g715(.A1(new_n590), .A2(new_n592), .ZN(new_n902));
  NAND2_X1  g716(.A1(G478), .A2(G902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT59), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n889), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n829), .B2(new_n847), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n865), .B1(new_n909), .B2(new_n902), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n910), .ZN(G63));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT123), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n866), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n614), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n498), .B(KEYINPUT124), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n916), .B(new_n865), .C1(new_n915), .C2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G66));
  INV_X1    g734(.A(G224), .ZN(new_n921));
  OAI21_X1  g735(.A(G953), .B1(new_n274), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n820), .A2(new_n831), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(G953), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n370), .B(new_n371), .C1(G898), .C2(new_n270), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(G69));
  NAND2_X1  g740(.A1(new_n519), .A2(new_n520), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n516), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n236), .A2(new_n240), .A3(new_n242), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n742), .A2(new_n749), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n779), .A2(new_n661), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n657), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT62), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n268), .A2(new_n655), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n711), .B(new_n638), .C1(new_n816), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n931), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n930), .B1(new_n937), .B2(new_n270), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(KEYINPUT125), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n740), .A2(new_n638), .A3(new_n679), .A4(new_n754), .ZN(new_n940));
  AND4_X1   g754(.A1(new_n813), .A2(new_n940), .A3(new_n714), .A4(new_n932), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n941), .A2(new_n742), .A3(new_n749), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n930), .B1(new_n943), .B2(new_n623), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n270), .B1(G227), .B2(G900), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G72));
  NAND2_X1  g761(.A1(G472), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT63), .Z(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n641), .B2(new_n569), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n828), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n568), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n931), .A2(new_n934), .A3(new_n923), .A4(new_n936), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n563), .B(new_n953), .C1(new_n954), .C2(new_n949), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n950), .B1(new_n942), .B2(new_n923), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(new_n563), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n885), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n885), .C1(new_n956), .C2(new_n958), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n952), .B(new_n955), .C1(new_n960), .C2(new_n962), .ZN(G57));
endmodule


