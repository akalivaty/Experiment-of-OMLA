//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985;
  XNOR2_X1  g000(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT2), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(KEYINPUT80), .A3(new_n212), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G141gat), .B(G148gat), .Z(new_n218));
  OAI211_X1 g017(.A(new_n218), .B(new_n208), .C1(KEYINPUT80), .C2(new_n214), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n225), .A2(new_n226), .B1(G211gat), .B2(G218gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n225), .B2(new_n226), .ZN(new_n228));
  XNOR2_X1  g027(.A(G197gat), .B(G204gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n230), .B(new_n231), .Z(new_n234));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n234), .B2(new_n223), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n219), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT81), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT81), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n233), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(G228gat), .A3(G233gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n233), .A2(KEYINPUT89), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n221), .B1(new_n232), .B2(KEYINPUT29), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n244), .A2(new_n236), .B1(G228gat), .B2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT89), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n224), .A2(new_n246), .A3(new_n232), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G78gat), .B(G106gat), .ZN(new_n249));
  INV_X1    g048(.A(G50gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT88), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n242), .A2(new_n248), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n242), .B2(new_n248), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n205), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n256), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(new_n204), .A3(new_n254), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT76), .ZN(new_n261));
  NAND2_X1  g060(.A1(G226gat), .A2(G233gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT65), .B(G176gat), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT23), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT24), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  INV_X1    g066(.A(G190gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n267), .A3(new_n268), .ZN(new_n271));
  NAND3_X1  g070(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G176gat), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT23), .B1(new_n264), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n264), .A2(new_n275), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n265), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT25), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n275), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT25), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n283), .A2(new_n277), .A3(new_n276), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n272), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n272), .A2(new_n285), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n267), .A2(new_n268), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n269), .A4(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n279), .A2(new_n280), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G183gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n293), .A3(new_n268), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT28), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n294), .B(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n277), .B1(KEYINPUT26), .B2(new_n281), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n281), .A2(KEYINPUT26), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n298), .A2(new_n299), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n290), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n261), .B(new_n262), .C1(new_n305), .C2(KEYINPUT29), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n279), .A2(new_n280), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n284), .A2(new_n289), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n301), .ZN(new_n310));
  INV_X1    g109(.A(new_n262), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n297), .A2(new_n303), .A3(new_n300), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n303), .B1(new_n297), .B2(new_n300), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n311), .B1(new_n316), .B2(new_n223), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(new_n261), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n232), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n305), .B2(new_n262), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(KEYINPUT78), .A3(new_n311), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT29), .B1(new_n309), .B2(new_n301), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT77), .B1(new_n323), .B2(new_n311), .ZN(new_n324));
  INV_X1    g123(.A(new_n301), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n223), .B1(new_n325), .B2(new_n290), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(new_n262), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n321), .A2(new_n322), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n234), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n333));
  XOR2_X1   g132(.A(G8gat), .B(G36gat), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT79), .ZN(new_n335));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n317), .A2(new_n261), .B1(new_n311), .B2(new_n310), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n262), .B1(new_n305), .B2(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT76), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n234), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n322), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n328), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n344), .A2(new_n234), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n339), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n319), .A2(new_n330), .A3(new_n337), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(KEYINPUT30), .A3(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n338), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n352), .A2(KEYINPUT1), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT70), .B(G120gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G113gat), .ZN(new_n355));
  INV_X1    g154(.A(G113gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G120gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(KEYINPUT71), .A3(new_n357), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n353), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G120gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G113gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n365), .A2(KEYINPUT69), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT1), .B1(new_n365), .B2(KEYINPUT69), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n351), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n238), .A2(KEYINPUT3), .A3(new_n239), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n352), .A2(KEYINPUT1), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n355), .A2(KEYINPUT71), .A3(new_n357), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT71), .B1(new_n355), .B2(new_n357), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n368), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n377), .A3(new_n222), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n220), .A3(new_n376), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n370), .A2(new_n378), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT85), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n379), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n239), .B(new_n238), .C1(new_n362), .C2(new_n368), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n380), .B1(new_n387), .B2(KEYINPUT83), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n238), .A2(new_n239), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n377), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n386), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n392), .A2(KEYINPUT84), .A3(new_n383), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n394), .B(new_n386), .C1(new_n388), .C2(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT5), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n385), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n395), .A2(KEYINPUT5), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(KEYINPUT84), .A3(new_n383), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n384), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT0), .ZN(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n397), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT39), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n370), .A2(new_n378), .ZN(new_n408));
  INV_X1    g207(.A(new_n382), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n407), .B(new_n386), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n410), .A2(new_n404), .ZN(new_n411));
  INV_X1    g210(.A(new_n391), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n390), .A2(new_n389), .A3(new_n377), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n379), .A4(new_n380), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n386), .B1(new_n408), .B2(new_n409), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT39), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n411), .A2(KEYINPUT40), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT40), .B1(new_n411), .B2(new_n416), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n350), .A2(new_n406), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n337), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n331), .B2(new_n339), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n329), .B2(new_n232), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n234), .B1(new_n313), .B2(new_n318), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT38), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT90), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT38), .B1(new_n424), .B2(new_n425), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT90), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n337), .B1(new_n319), .B2(new_n330), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n422), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n348), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n332), .A2(new_n421), .B1(new_n432), .B2(new_n422), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(KEYINPUT38), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n397), .A2(new_n400), .A3(new_n405), .A4(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n406), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n405), .B1(new_n397), .B2(new_n400), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n260), .B(new_n420), .C1(new_n438), .C2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT34), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n316), .A2(new_n369), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n377), .B(new_n309), .C1(new_n315), .C2(new_n314), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G227gat), .ZN(new_n450));
  INV_X1    g249(.A(G233gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n446), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  AOI211_X1 g253(.A(KEYINPUT34), .B(new_n452), .C1(new_n447), .C2(new_n448), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n447), .A2(new_n452), .A3(new_n448), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT32), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G15gat), .B(G43gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT72), .ZN(new_n462));
  XOR2_X1   g261(.A(G71gat), .B(G99gat), .Z(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n457), .B(KEYINPUT32), .C1(new_n459), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n456), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT74), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n456), .A2(new_n465), .A3(new_n470), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n456), .B1(new_n467), .B2(new_n465), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n449), .A2(new_n453), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT34), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n449), .A2(new_n446), .A3(new_n453), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(KEYINPUT73), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT73), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n454), .B2(new_n455), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n467), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n469), .A2(new_n471), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n476), .B1(new_n485), .B2(new_n473), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n338), .A2(new_n349), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n444), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n260), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n483), .A2(new_n484), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n472), .A2(new_n260), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n444), .A2(new_n492), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT35), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n393), .A2(new_n385), .A3(new_n396), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n384), .B1(new_n398), .B2(new_n399), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n404), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n406), .A3(new_n441), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT35), .B1(new_n498), .B2(new_n440), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n474), .B1(new_n469), .B2(new_n471), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n487), .A2(new_n500), .A3(new_n260), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n445), .A2(new_n490), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(G71gat), .A2(G78gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(G57gat), .A2(G64gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(G57gat), .A2(G64gat), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n508), .B(new_n509), .C1(new_n504), .C2(KEYINPUT9), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT99), .B1(G71gat), .B2(G78gat), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT21), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G231gat), .A2(G233gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G127gat), .B(G155gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT100), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n518), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G183gat), .B(G211gat), .Z(new_n522));
  AND2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n203), .A2(G15gat), .ZN(new_n525));
  INV_X1    g324(.A(G15gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n525), .B2(new_n527), .ZN(new_n530));
  OAI211_X1 g329(.A(KEYINPUT95), .B(G1gat), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n529), .B2(new_n530), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n526), .A2(G22gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n203), .A2(G15gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT94), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(G1gat), .B1(new_n539), .B2(KEYINPUT95), .ZN(new_n540));
  OAI21_X1  g339(.A(G8gat), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT95), .B1(new_n529), .B2(new_n530), .ZN(new_n542));
  INV_X1    g341(.A(G1gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G8gat), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n531), .A4(new_n533), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n541), .B(new_n546), .C1(new_n515), .C2(new_n514), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  OR3_X1    g348(.A1(new_n523), .A2(new_n524), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n523), .B2(new_n524), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G43gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(G50gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n250), .A2(G43gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G29gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT14), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(G36gat), .ZN(new_n560));
  INV_X1    g359(.A(G36gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT14), .A3(G29gat), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT92), .B1(new_n559), .B2(G36gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(KEYINPUT15), .B(new_n557), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n555), .B2(new_n556), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n250), .A2(G43gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n554), .A2(G50gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT15), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n560), .A2(new_n562), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n568), .A2(new_n571), .A3(new_n572), .A4(new_n564), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(new_n566), .B2(new_n573), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n576), .B(KEYINPUT17), .C1(new_n575), .C2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580));
  INV_X1    g379(.A(new_n574), .ZN(new_n581));
  OAI211_X1 g380(.A(KEYINPUT96), .B(new_n580), .C1(new_n581), .C2(new_n577), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT101), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT101), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT7), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n584), .A2(KEYINPUT101), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n588), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G99gat), .B(G106gat), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(new_n588), .A3(new_n590), .A4(new_n594), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n581), .B2(new_n600), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT102), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n608), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n601), .A2(new_n613), .A3(new_n605), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n612), .B1(new_n609), .B2(new_n614), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n553), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n597), .B(new_n599), .C1(new_n512), .C2(new_n513), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n622), .A3(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n514), .A2(new_n600), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n621), .ZN(new_n630));
  INV_X1    g429(.A(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n629), .A2(new_n632), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n620), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G113gat), .B(G141gat), .Z(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G169gat), .B(G197gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n541), .A2(new_n546), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n574), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT97), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(new_n579), .B2(new_n582), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI211_X1 g453(.A(KEYINPUT97), .B(new_n650), .C1(new_n582), .C2(new_n579), .ZN(new_n655));
  OAI211_X1 g454(.A(KEYINPUT18), .B(new_n649), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n650), .B(new_n574), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n649), .B(KEYINPUT13), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n653), .B2(new_n652), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT18), .B1(new_n663), .B2(new_n649), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n648), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT18), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n668), .A2(new_n656), .A3(new_n659), .A4(new_n647), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(KEYINPUT98), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n671), .B(new_n648), .C1(new_n660), .C2(new_n664), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n641), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT104), .B1(new_n503), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n419), .A2(new_n406), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n260), .B1(new_n679), .B2(new_n487), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n434), .A2(new_n437), .ZN(new_n681));
  INV_X1    g480(.A(new_n444), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n473), .B1(new_n472), .B2(new_n491), .ZN(new_n684));
  AOI211_X1 g483(.A(KEYINPUT36), .B(new_n474), .C1(new_n469), .C2(new_n471), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n350), .B1(new_n498), .B2(new_n440), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n687), .B2(new_n260), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n493), .A2(KEYINPUT35), .B1(new_n499), .B2(new_n501), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n677), .B(new_n678), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n676), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n444), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n543), .ZN(G1324gat));
  OAI21_X1  g493(.A(G8gat), .B1(new_n692), .B2(new_n487), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n487), .B1(new_n676), .B2(new_n691), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n698), .ZN(new_n702));
  AOI211_X1 g501(.A(new_n487), .B(new_n702), .C1(new_n676), .C2(new_n691), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(new_n696), .A3(KEYINPUT42), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT42), .B1(new_n703), .B2(new_n696), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n695), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(G1325gat));
  OAI21_X1  g509(.A(G15gat), .B1(new_n692), .B2(new_n686), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n500), .A2(new_n526), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n692), .B2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n692), .A2(new_n260), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n503), .A2(new_n619), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n673), .A2(new_n553), .A3(new_n640), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n718), .A2(new_n558), .A3(new_n682), .A4(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT45), .Z(new_n721));
  INV_X1    g520(.A(new_n719), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n490), .A2(new_n445), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n494), .A2(new_n502), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n618), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT44), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n616), .B2(new_n617), .ZN(new_n729));
  INV_X1    g528(.A(new_n617), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(KEYINPUT107), .A3(new_n615), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n503), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n722), .B1(new_n727), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n558), .B1(new_n737), .B2(new_n682), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n717), .B1(new_n721), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n738), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n720), .B(KEYINPUT45), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT108), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(G1328gat));
  NAND2_X1  g542(.A1(new_n718), .A2(new_n719), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(G36gat), .A3(new_n487), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n736), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n719), .ZN(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n748), .B2(new_n487), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n737), .A2(new_n486), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G43gat), .ZN(new_n753));
  INV_X1    g552(.A(new_n500), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n744), .A2(G43gat), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n751), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  AOI211_X1 g556(.A(KEYINPUT47), .B(new_n755), .C1(new_n752), .C2(G43gat), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(G1330gat));
  OAI21_X1  g558(.A(new_n250), .B1(new_n744), .B2(new_n260), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n489), .A2(G50gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n748), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g562(.A(new_n640), .ZN(new_n764));
  NOR4_X1   g563(.A1(new_n503), .A2(new_n674), .A3(new_n620), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n682), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n350), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT49), .B(G64gat), .Z(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(G1333gat));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n486), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n754), .A2(G71gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(G71gat), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n765), .A2(new_n489), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT109), .B(G78gat), .Z(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n674), .A2(new_n553), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n640), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT110), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n747), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n444), .ZN(new_n783));
  INV_X1    g582(.A(new_n779), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT51), .B1(new_n726), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n718), .A2(new_n786), .A3(new_n779), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n787), .A3(new_n640), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n682), .A2(new_n592), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n783), .B1(new_n788), .B2(new_n789), .ZN(G1336gat));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n487), .A2(G92gat), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n785), .A2(new_n787), .A3(new_n640), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(new_n793), .B2(KEYINPUT111), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n733), .B1(new_n725), .B2(new_n618), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n350), .B(new_n781), .C1(new_n795), .C2(new_n735), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G92gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n793), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n794), .B(new_n798), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n782), .B2(new_n686), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n754), .A2(G99gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n788), .B2(new_n801), .ZN(G1338gat));
  OAI211_X1 g601(.A(new_n489), .B(new_n781), .C1(new_n795), .C2(new_n735), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G106gat), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n804), .B2(KEYINPUT112), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n260), .A2(G106gat), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n785), .A2(new_n787), .A3(new_n640), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n804), .B(new_n807), .C1(KEYINPUT112), .C2(KEYINPUT53), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(G1339gat));
  NAND2_X1  g610(.A1(new_n627), .A2(new_n628), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT10), .B1(new_n621), .B2(new_n622), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(new_n631), .A3(new_n813), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n815));
  AOI21_X1  g614(.A(new_n636), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n631), .B1(new_n812), .B2(new_n813), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT54), .A3(new_n629), .ZN(new_n818));
  AOI211_X1 g617(.A(KEYINPUT115), .B(KEYINPUT55), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n812), .A2(new_n813), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n626), .A3(new_n815), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n637), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n823), .B2(new_n824), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n816), .A2(new_n828), .A3(KEYINPUT55), .A4(new_n818), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n639), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n670), .A3(new_n672), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n663), .A2(new_n649), .B1(new_n657), .B2(new_n658), .ZN(new_n833));
  INV_X1    g632(.A(new_n646), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n669), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n640), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n732), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n732), .A2(new_n836), .A3(new_n831), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n552), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n641), .A2(new_n673), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n444), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n501), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n356), .B1(new_n844), .B2(new_n674), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT116), .Z(new_n846));
  AND2_X1   g645(.A1(new_n843), .A2(new_n492), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(new_n487), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n356), .A3(new_n674), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(G1340gat));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n354), .A3(new_n640), .ZN(new_n851));
  INV_X1    g650(.A(new_n844), .ZN(new_n852));
  OAI21_X1  g651(.A(G120gat), .B1(new_n852), .B2(new_n764), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n848), .A2(new_n855), .A3(new_n553), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n852), .B2(new_n552), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  OAI21_X1  g657(.A(G134gat), .B1(new_n852), .B2(new_n619), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n487), .A2(new_n618), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(G134gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n847), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n862), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT117), .B1(new_n862), .B2(KEYINPUT56), .ZN(new_n864));
  OAI221_X1 g663(.A(new_n859), .B1(KEYINPUT56), .B2(new_n862), .C1(new_n863), .C2(new_n864), .ZN(G1343gat));
  NAND3_X1  g664(.A1(new_n686), .A2(new_n682), .A3(new_n487), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n674), .A2(G141gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n842), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n868), .B2(new_n489), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n489), .A2(KEYINPUT57), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n823), .A2(new_n824), .ZN(new_n871));
  AND4_X1   g670(.A1(new_n639), .A2(new_n827), .A3(new_n829), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n670), .A2(new_n672), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n618), .B1(new_n873), .B2(new_n837), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n839), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT118), .B(new_n618), .C1(new_n873), .C2(new_n837), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n552), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n870), .B1(new_n878), .B2(new_n842), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n869), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n842), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n873), .A2(new_n837), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n619), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT118), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n874), .A2(new_n875), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n839), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n882), .B1(new_n887), .B2(new_n552), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT119), .B1(new_n888), .B2(new_n870), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n866), .B(new_n867), .C1(new_n881), .C2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n843), .A2(new_n489), .A3(new_n686), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n350), .ZN(new_n893));
  AOI21_X1  g692(.A(G141gat), .B1(new_n893), .B2(new_n674), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(KEYINPUT58), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n890), .B2(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1344gat));
  NAND3_X1  g698(.A1(new_n893), .A2(new_n210), .A3(new_n640), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n868), .A2(new_n489), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n831), .A2(new_n836), .A3(new_n618), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n552), .B1(new_n874), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n842), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n260), .A2(KEYINPUT57), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n901), .A2(KEYINPUT57), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n866), .A2(new_n764), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n908), .C2(new_n210), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n210), .B1(new_n906), .B2(new_n907), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(G148gat), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n866), .B1(new_n881), .B2(new_n889), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n640), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n900), .B1(new_n914), .B2(new_n917), .ZN(G1345gat));
  NAND3_X1  g717(.A1(new_n893), .A2(new_n206), .A3(new_n553), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n916), .A2(new_n553), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n206), .ZN(G1346gat));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n207), .B1(new_n916), .B2(new_n732), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n892), .A2(G162gat), .A3(new_n860), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n924), .ZN(new_n926));
  INV_X1    g725(.A(new_n732), .ZN(new_n927));
  AOI211_X1 g726(.A(new_n927), .B(new_n866), .C1(new_n881), .C2(new_n889), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT121), .B(new_n926), .C1(new_n928), .C2(new_n207), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n929), .ZN(G1347gat));
  AOI21_X1  g729(.A(new_n487), .B1(new_n498), .B2(new_n440), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n868), .A2(new_n492), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n674), .ZN(new_n933));
  AND4_X1   g732(.A1(new_n260), .A2(new_n868), .A3(new_n500), .A4(new_n931), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n673), .A2(new_n264), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G1348gat));
  AOI21_X1  g735(.A(G176gat), .B1(new_n932), .B2(new_n640), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n764), .A2(new_n263), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n934), .B2(new_n938), .ZN(G1349gat));
  NAND4_X1  g738(.A1(new_n932), .A2(new_n291), .A3(new_n293), .A4(new_n553), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n934), .A2(new_n553), .ZN(new_n942));
  OAI221_X1 g741(.A(new_n940), .B1(KEYINPUT122), .B2(new_n941), .C1(new_n942), .C2(new_n267), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(KEYINPUT122), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1350gat));
  AOI21_X1  g744(.A(new_n268), .B1(new_n934), .B2(new_n618), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT61), .Z(new_n947));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n268), .A3(new_n732), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1351gat));
  AOI21_X1  g748(.A(new_n260), .B1(new_n841), .B2(new_n842), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(new_n686), .A3(new_n931), .ZN(new_n951));
  AOI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n674), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n904), .A2(new_n905), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n686), .A2(new_n931), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT57), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n953), .B(new_n955), .C1(new_n950), .C2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n674), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  INV_X1    g759(.A(G204gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n951), .A2(new_n961), .A3(new_n640), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT124), .ZN(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n957), .B2(new_n764), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G1353gat));
  INV_X1    g766(.A(G211gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n968), .A3(new_n553), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n906), .A2(new_n686), .A3(new_n553), .A4(new_n931), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n901), .A2(KEYINPUT57), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n975), .A2(KEYINPUT125), .A3(new_n953), .A4(new_n955), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n957), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n976), .A2(new_n978), .A3(new_n618), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G218gat), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n927), .A2(G218gat), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n951), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n974), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(new_n982), .ZN(new_n984));
  AOI211_X1 g783(.A(KEYINPUT126), .B(new_n984), .C1(new_n979), .C2(G218gat), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n983), .A2(new_n985), .ZN(G1355gat));
endmodule


