//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n203), .B1(KEYINPUT23), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT23), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n215));
  AND4_X1   g014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT68), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G183gat), .B2(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n209), .B1(new_n216), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT64), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .A4(new_n222), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n207), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n232), .A2(KEYINPUT23), .A3(new_n206), .A4(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n206), .A2(new_n207), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n224), .A2(KEYINPUT25), .B1(new_n230), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT27), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(G183gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(G183gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT69), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(G190gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n245), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n247), .A3(new_n218), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n249), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT26), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n210), .B1(new_n237), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n203), .A2(KEYINPUT26), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n204), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n252), .B1(new_n251), .B2(new_n254), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n240), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n267), .A3(new_n271), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n265), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n266), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n278), .B1(new_n262), .B2(new_n263), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n251), .A2(new_n254), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n255), .A3(new_n259), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n265), .B1(new_n286), .B2(new_n240), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT74), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n281), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n202), .B(new_n280), .C1(new_n289), .C2(new_n277), .ZN(new_n290));
  XOR2_X1   g089(.A(G8gat), .B(G36gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT75), .ZN(new_n292));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n280), .B1(new_n289), .B2(new_n277), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(KEYINPUT37), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n290), .B1(new_n297), .B2(KEYINPUT88), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT88), .ZN(new_n299));
  AOI211_X1 g098(.A(new_n299), .B(new_n295), .C1(new_n296), .C2(KEYINPUT37), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT38), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n277), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n281), .A2(new_n302), .A3(new_n287), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n262), .A2(KEYINPUT74), .A3(new_n278), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT74), .B1(new_n262), .B2(new_n278), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n266), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n303), .B1(new_n306), .B2(new_n302), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n295), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n266), .B(new_n277), .C1(new_n304), .C2(new_n305), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n302), .B1(new_n281), .B2(new_n287), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n309), .A2(KEYINPUT87), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT37), .B1(new_n309), .B2(KEYINPUT87), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n295), .A2(KEYINPUT38), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n290), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n308), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT0), .ZN(new_n319));
  XNOR2_X1  g118(.A(G57gat), .B(G85gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  INV_X1    g121(.A(G155gat), .ZN(new_n323));
  INV_X1    g122(.A(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G141gat), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n322), .B(new_n325), .C1(new_n330), .C2(KEYINPUT2), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(new_n322), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n325), .A2(new_n334), .A3(new_n322), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(KEYINPUT76), .A3(new_n329), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT2), .ZN(new_n338));
  XOR2_X1   g137(.A(G141gat), .B(G148gat), .Z(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(KEYINPUT76), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n331), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(KEYINPUT1), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G113gat), .B(G120gat), .Z(new_n345));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n346));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT79), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(KEYINPUT78), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n344), .A2(new_n348), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n355), .B(new_n331), .C1(new_n337), .C2(new_n340), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n353), .A2(new_n351), .A3(new_n354), .A4(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n354), .B(new_n331), .C1(new_n340), .C2(new_n337), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n354), .B1(new_n341), .B2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n365), .B(new_n331), .C1(new_n337), .C2(new_n340), .ZN(new_n366));
  AOI211_X1 g165(.A(KEYINPUT5), .B(new_n363), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT4), .A3(new_n354), .A4(new_n356), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(new_n349), .A3(new_n366), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n351), .B1(new_n341), .B2(new_n349), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n369), .A2(new_n371), .A3(new_n362), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n341), .A2(new_n349), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n376), .B2(new_n363), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n321), .B1(new_n368), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n317), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n361), .A2(new_n367), .B1(new_n373), .B2(new_n377), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT6), .B1(new_n383), .B2(new_n321), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n380), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n316), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n301), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G22gat), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT3), .B1(new_n277), .B2(new_n263), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n341), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n366), .A2(new_n263), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n302), .ZN(new_n395));
  NAND2_X1  g194(.A1(G228gat), .A2(G233gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(new_n394), .B2(new_n302), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT83), .B(new_n277), .C1(new_n366), .C2(new_n263), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n391), .B1(new_n353), .B2(new_n356), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n390), .B(new_n398), .C1(new_n403), .C2(new_n397), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT84), .ZN(new_n405));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT31), .B(G50gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n398), .B1(new_n403), .B2(new_n397), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G22gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n404), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n411), .A2(new_n414), .A3(new_n404), .A4(new_n408), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n296), .A2(new_n294), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n308), .A3(KEYINPUT30), .ZN(new_n418));
  OR3_X1    g217(.A1(new_n296), .A2(KEYINPUT30), .A3(new_n294), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n362), .B1(new_n361), .B2(new_n371), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n321), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT39), .B1(new_n376), .B2(new_n363), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n421), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n321), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n422), .B2(new_n423), .ZN(new_n430));
  INV_X1    g229(.A(new_n421), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n430), .B(new_n431), .C1(new_n422), .C2(new_n426), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n428), .A2(new_n432), .A3(new_n380), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n416), .B1(new_n420), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n389), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n349), .A2(KEYINPUT71), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n349), .A2(KEYINPUT71), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n262), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(G227gat), .A2(G233gat), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n286), .A2(KEYINPUT71), .A3(new_n349), .A4(new_n240), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(KEYINPUT32), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT72), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n441), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n441), .A2(new_n445), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n441), .B2(KEYINPUT32), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n449), .A2(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT73), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n454), .B2(new_n456), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n454), .A2(new_n456), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n453), .A2(new_n460), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT36), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n449), .A2(new_n450), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n452), .A2(new_n451), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  OAI22_X1  g265(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(new_n457), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n460), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n418), .A2(new_n419), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n368), .A2(new_n378), .A3(new_n321), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n381), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n383), .B2(new_n321), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n368), .A2(new_n378), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(KEYINPUT80), .A3(new_n429), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT81), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n386), .B(new_n382), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n479), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n481), .A3(new_n384), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n473), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n416), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n435), .A2(new_n472), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n415), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n405), .A2(new_n408), .B1(new_n411), .B2(new_n404), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n469), .A3(new_n467), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT35), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n467), .A2(new_n469), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n420), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n387), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n488), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT99), .ZN(new_n502));
  XNOR2_X1  g301(.A(G134gat), .B(G162gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n506));
  XOR2_X1   g305(.A(G99gat), .B(G106gat), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509));
  INV_X1    g308(.A(G85gat), .ZN(new_n510));
  INV_X1    g309(.A(G92gat), .ZN(new_n511));
  AOI22_X1  g310(.A1(KEYINPUT8), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n512), .B(KEYINPUT102), .Z(new_n513));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(G85gat), .B2(G92gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT100), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(G85gat), .A3(G92gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT101), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n508), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n513), .A2(new_n519), .A3(new_n508), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT14), .B(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G29gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G43gat), .B(G50gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT15), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT89), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n530), .A2(KEYINPUT15), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n529), .A2(new_n532), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n534), .A2(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n506), .B1(new_n523), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT103), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(KEYINPUT103), .B(new_n506), .C1(new_n523), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G190gat), .B(G218gat), .Z(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n534), .A2(new_n536), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n539), .A2(new_n540), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT94), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n541), .A2(new_n554), .A3(KEYINPUT17), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n541), .B2(KEYINPUT17), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n553), .B(new_n523), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n546), .A2(new_n548), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n548), .B1(new_n546), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n505), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G64gat), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n562), .A2(G57gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(G57gat), .ZN(new_n564));
  INV_X1    g363(.A(G71gat), .ZN(new_n565));
  INV_X1    g364(.A(G78gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI22_X1  g366(.A1(new_n563), .A2(new_n564), .B1(new_n567), .B2(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n571), .B2(new_n573), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n575), .A2(new_n576), .A3(G127gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(G127gat), .B1(new_n575), .B2(new_n576), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G127gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n576), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(new_n574), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n579), .B1(new_n585), .B2(new_n577), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n323), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(G8gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(G15gat), .B(G22gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT92), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G1gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT16), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(new_n592), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n593), .A3(G1gat), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n591), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n590), .A2(G8gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n570), .A2(KEYINPUT21), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n602), .B1(new_n601), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n589), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  INV_X1    g407(.A(new_n589), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n587), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n582), .A2(new_n607), .A3(new_n610), .A4(new_n586), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n546), .A2(new_n557), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n547), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n504), .A3(new_n558), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n561), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT104), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT104), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n561), .A2(new_n617), .A3(new_n614), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n601), .B(new_n553), .C1(new_n555), .C2(new_n556), .ZN(new_n623));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT95), .Z(new_n625));
  OR2_X1    g424(.A1(new_n601), .A2(new_n541), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n623), .A2(KEYINPUT18), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n601), .B(new_n551), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n625), .B(KEYINPUT13), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G197gat), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT11), .B(G169gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n627), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT18), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT96), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n642), .A3(new_n639), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(new_n631), .A3(new_n627), .ZN(new_n645));
  INV_X1    g444(.A(new_n636), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n521), .A2(new_n570), .A3(new_n522), .ZN(new_n650));
  INV_X1    g449(.A(new_n522), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n571), .B1(new_n651), .B2(new_n520), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT105), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n649), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n650), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n650), .A2(new_n652), .A3(new_n660), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n653), .A2(KEYINPUT105), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n658), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n657), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n663), .B2(new_n653), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n622), .A2(new_n648), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n500), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT106), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n500), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n482), .A2(new_n485), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g477(.A(KEYINPUT16), .B(G8gat), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n675), .A2(new_n420), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n680), .B2(G8gat), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  INV_X1    g483(.A(new_n674), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n673), .B1(new_n500), .B2(new_n670), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n420), .B(new_n684), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n683), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n683), .B(new_n693), .C1(new_n689), .C2(new_n690), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(G1325gat));
  INV_X1    g494(.A(G15gat), .ZN(new_n696));
  INV_X1    g495(.A(new_n494), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n675), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n472), .B1(new_n672), .B2(new_n674), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(new_n696), .ZN(G1326gat));
  NAND2_X1  g499(.A1(new_n675), .A2(new_n416), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT43), .B(G22gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n471), .B1(new_n389), .B2(new_n434), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(new_n487), .B1(new_n493), .B2(new_n498), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n561), .A2(new_n617), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n704), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n500), .A2(KEYINPUT44), .A3(new_n707), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n648), .A2(new_n614), .A3(new_n669), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT109), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n709), .A2(new_n710), .A3(new_n714), .A4(new_n711), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n676), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G29gat), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n500), .A2(new_n707), .A3(new_n711), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n527), .A3(new_n676), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT110), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n717), .A2(new_n723), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1328gat));
  NAND3_X1  g524(.A1(new_n713), .A2(new_n420), .A3(new_n715), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G36gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n718), .A2(new_n525), .A3(new_n420), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n727), .A2(KEYINPUT111), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1329gat));
  OAI21_X1  g534(.A(G43gat), .B1(new_n712), .B2(new_n472), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n494), .A2(G43gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(KEYINPUT47), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n713), .A2(new_n471), .A3(new_n715), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n740), .A2(G43gat), .B1(new_n718), .B2(new_n737), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n741), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g541(.A1(new_n713), .A2(new_n416), .A3(new_n715), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n491), .A2(G50gat), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n743), .A2(G50gat), .B1(new_n718), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(G50gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n712), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(new_n416), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n718), .A2(new_n744), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT48), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n745), .A2(KEYINPUT48), .B1(new_n748), .B2(new_n750), .ZN(G1331gat));
  INV_X1    g550(.A(new_n648), .ZN(new_n752));
  INV_X1    g551(.A(new_n669), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n622), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n500), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n676), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g557(.A1(new_n755), .A2(new_n473), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n755), .B2(new_n472), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n697), .A2(new_n565), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n755), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n755), .A2(new_n491), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n566), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n752), .A2(new_n614), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n669), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n709), .A2(new_n710), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n676), .ZN(new_n775));
  OAI21_X1  g574(.A(G85gat), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n500), .A2(new_n707), .A3(new_n771), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n676), .A2(new_n510), .A3(new_n669), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(G1336gat));
  OAI21_X1  g581(.A(G92gat), .B1(new_n774), .B2(new_n473), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n420), .A2(new_n511), .A3(new_n669), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g585(.A(G99gat), .B1(new_n774), .B2(new_n472), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n494), .A2(new_n753), .A3(G99gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n780), .B2(new_n788), .ZN(G1338gat));
  INV_X1    g588(.A(G106gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n774), .A2(new_n790), .A3(new_n491), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(KEYINPUT53), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(KEYINPUT53), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n753), .A2(new_n491), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n779), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n794), .B(new_n795), .C1(new_n797), .C2(G106gat), .ZN(new_n798));
  AOI21_X1  g597(.A(G106gat), .B1(new_n779), .B2(new_n796), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n792), .B(KEYINPUT53), .C1(new_n799), .C2(new_n791), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n622), .A2(new_n669), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n625), .B1(new_n623), .B2(new_n626), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n628), .A2(new_n630), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n635), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(KEYINPUT114), .B(new_n635), .C1(new_n803), .C2(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n663), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n661), .A2(new_n662), .A3(new_n659), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n657), .B1(new_n663), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n665), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n814), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n809), .A2(new_n817), .A3(new_n644), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n614), .B1(new_n819), .B2(new_n707), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n809), .A2(new_n644), .A3(new_n669), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n818), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n821), .B(new_n708), .C1(new_n648), .C2(new_n822), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n802), .A2(new_n648), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n775), .A3(new_n416), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n495), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n752), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n669), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(G120gat), .ZN(G1341gat));
  INV_X1    g630(.A(new_n614), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(new_n583), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n707), .A2(new_n473), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(G134gat), .A3(new_n494), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n826), .B2(new_n708), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1343gat));
  NOR3_X1   g640(.A1(new_n775), .A2(new_n471), .A3(new_n420), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n824), .B2(new_n491), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n820), .A2(new_n823), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n648), .A2(new_n619), .A3(new_n621), .A4(new_n753), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT57), .A3(new_n416), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n843), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(G141gat), .A3(new_n752), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n824), .A2(new_n491), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n775), .A2(new_n471), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n852), .A2(new_n473), .A3(new_n752), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n326), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n851), .B(new_n855), .C1(KEYINPUT116), .C2(KEYINPUT58), .ZN(new_n856));
  NAND2_X1  g655(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n856), .B(new_n857), .ZN(G1344gat));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n753), .B1(new_n843), .B2(KEYINPUT117), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n619), .A2(new_n621), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n861), .A2(KEYINPUT118), .A3(new_n648), .A4(new_n753), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n846), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n865), .B2(new_n416), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n844), .B(new_n491), .C1(new_n846), .C2(new_n847), .ZN(new_n867));
  OAI221_X1 g666(.A(new_n860), .B1(KEYINPUT117), .B2(new_n843), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n859), .B1(new_n868), .B2(G148gat), .ZN(new_n869));
  AOI211_X1 g668(.A(KEYINPUT59), .B(new_n327), .C1(new_n850), .C2(new_n669), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n852), .A2(new_n473), .A3(new_n853), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n669), .A2(new_n327), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n869), .A2(new_n870), .B1(new_n871), .B2(new_n872), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n832), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n875));
  AOI21_X1  g674(.A(G155gat), .B1(new_n874), .B2(KEYINPUT119), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n832), .A2(new_n323), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n875), .A2(new_n876), .B1(new_n850), .B2(new_n877), .ZN(G1346gat));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n848), .B2(new_n416), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n842), .B1(new_n879), .B2(new_n867), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT120), .B1(new_n880), .B2(new_n708), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n850), .A2(new_n882), .A3(new_n707), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n883), .A3(G162gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n835), .A2(G162gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n852), .A2(new_n853), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n884), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n824), .A2(new_n416), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n676), .A2(new_n473), .A3(new_n494), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(new_n206), .A3(new_n648), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n824), .A2(new_n676), .ZN(new_n896));
  INV_X1    g695(.A(new_n492), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n420), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n752), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n895), .B1(new_n900), .B2(new_n206), .ZN(G1348gat));
  AOI21_X1  g700(.A(G176gat), .B1(new_n899), .B2(new_n669), .ZN(new_n902));
  INV_X1    g701(.A(new_n894), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n753), .B1(new_n232), .B2(new_n233), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(G1349gat));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n899), .A2(new_n245), .A3(new_n248), .A4(new_n614), .ZN(new_n908));
  OAI21_X1  g707(.A(G183gat), .B1(new_n894), .B2(new_n832), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n894), .B2(new_n708), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT61), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n218), .A3(new_n707), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1351gat));
  NOR3_X1   g715(.A1(new_n471), .A2(new_n491), .A3(new_n473), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n896), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(G197gat), .A3(new_n648), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n866), .B2(new_n867), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n820), .A2(new_n823), .B1(new_n847), .B2(new_n863), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n491), .B1(new_n922), .B2(new_n862), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT123), .B(new_n849), .C1(new_n923), .C2(KEYINPUT57), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n676), .A2(new_n473), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n472), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n921), .A2(new_n752), .A3(new_n924), .A4(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n919), .B1(new_n928), .B2(G197gat), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT124), .B(new_n919), .C1(new_n928), .C2(G197gat), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(G1352gat));
  NAND4_X1  g732(.A1(new_n921), .A2(new_n669), .A3(new_n924), .A4(new_n927), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT125), .B(G204gat), .Z(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n753), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n896), .A2(new_n917), .A3(new_n937), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT62), .Z(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1353gat));
  INV_X1    g743(.A(new_n918), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n269), .A3(new_n614), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n926), .A2(new_n832), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(new_n866), .B2(new_n867), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g752(.A(KEYINPUT127), .B(new_n946), .C1(new_n949), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1354gat));
  AOI21_X1  g754(.A(G218gat), .B1(new_n945), .B2(new_n707), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n921), .A2(new_n924), .A3(new_n927), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n708), .A2(new_n270), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(G1355gat));
endmodule


