//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT10), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT64), .A2(G143), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G146), .A3(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n191), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n194), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT64), .A2(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT64), .A2(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n195), .B1(new_n202), .B2(G146), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(G146), .B1(new_n192), .B2(new_n193), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  OAI21_X1  g020(.A(G128), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n199), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G104), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT72), .B1(new_n212), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT72), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n210), .A3(G104), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(KEYINPUT73), .A3(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G101), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n210), .A3(G104), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(G107), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n219), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n189), .B1(new_n208), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n194), .A2(new_n227), .A3(new_n196), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G128), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n200), .B2(new_n201), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(G143), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT65), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n194), .A2(new_n227), .A3(new_n196), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n192), .A2(new_n193), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n232), .B1(new_n238), .B2(new_n230), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n236), .B(new_n237), .C1(new_n239), .C2(new_n229), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n219), .A2(new_n221), .A3(new_n223), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G101), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(G101), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n235), .A2(new_n240), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G137), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .A3(G134), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n249), .A2(new_n251), .A3(new_n255), .A4(new_n252), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(G128), .B1(new_n195), .B2(new_n206), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n205), .B2(new_n232), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n194), .A2(new_n196), .A3(new_n198), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n189), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n224), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n262), .B1(G101), .B2(new_n217), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n226), .A2(new_n246), .A3(new_n257), .A4(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n197), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n260), .B1(new_n268), .B2(new_n203), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n270), .A2(new_n189), .B1(new_n263), .B2(new_n261), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n271), .A2(KEYINPUT74), .A3(new_n257), .A4(new_n246), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n254), .A2(new_n256), .ZN(new_n274));
  INV_X1    g088(.A(new_n270), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n225), .A2(new_n259), .A3(new_n260), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT12), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT12), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G110), .B(G140), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G227), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n282), .B(new_n284), .Z(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n273), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n271), .A2(new_n246), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n274), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n286), .B1(new_n273), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n187), .B(new_n188), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(G469), .A2(G902), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n273), .A2(new_n289), .A3(new_n286), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n267), .A2(new_n272), .B1(new_n279), .B2(new_n280), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n285), .B(KEYINPUT71), .Z(new_n295));
  OAI211_X1 g109(.A(new_n293), .B(G469), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  OAI21_X1  g115(.A(G125), .B1(new_n228), .B2(new_n234), .ZN(new_n302));
  INV_X1    g116(.A(G125), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n259), .A2(new_n303), .A3(new_n260), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(KEYINPUT76), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n259), .A2(new_n306), .A3(new_n303), .A4(new_n260), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n283), .A2(G224), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT7), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n305), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n305), .B2(new_n307), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G113), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G119), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G116), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT5), .ZN(new_n321));
  XNOR2_X1  g135(.A(G116), .B(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(KEYINPUT2), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G113), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n317), .A2(new_n321), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n218), .A3(new_n224), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT75), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n326), .A2(new_n322), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n322), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n245), .A2(new_n332), .A3(new_n243), .ZN(new_n333));
  XOR2_X1   g147(.A(G110), .B(G122), .Z(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n327), .A2(new_n218), .A3(new_n336), .A4(new_n224), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n329), .A2(new_n333), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT77), .B(KEYINPUT8), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n334), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n328), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n327), .B1(new_n224), .B2(new_n218), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(G902), .B1(new_n312), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n329), .A2(new_n333), .A3(new_n337), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n334), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n305), .A2(new_n308), .A3(new_n307), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n308), .B1(new_n305), .B2(new_n307), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n352), .A3(new_n334), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G210), .B1(G237), .B2(G902), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n345), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(new_n345), .B2(new_n354), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n301), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n360), .B(new_n301), .C1(new_n356), .C2(new_n357), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n363), .A2(new_n283), .A3(G143), .A4(G214), .ZN(new_n364));
  INV_X1    g178(.A(G214), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n365), .A2(G237), .A3(G953), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n362), .B(new_n364), .C1(new_n238), .C2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(KEYINPUT79), .A3(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT18), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(new_n255), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n367), .A2(KEYINPUT18), .A3(G131), .A4(new_n368), .ZN(new_n372));
  INV_X1    g186(.A(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G125), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n303), .A2(G140), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n375), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(G146), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n230), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n371), .A2(new_n372), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT16), .ZN(new_n386));
  OR3_X1    g200(.A1(new_n303), .A2(KEYINPUT16), .A3(G140), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n386), .A2(G146), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(G146), .B1(new_n386), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n367), .A2(G131), .A3(new_n368), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT17), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n369), .A2(new_n255), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n392), .A3(new_n391), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n394), .A2(KEYINPUT81), .A3(new_n392), .A4(new_n391), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n385), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n212), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT83), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(G902), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n395), .A2(new_n396), .ZN(new_n406));
  INV_X1    g220(.A(new_n393), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n398), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n384), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n403), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G475), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n394), .A2(new_n391), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n386), .A2(new_n387), .A3(G146), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT19), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n377), .B2(new_n380), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n376), .A2(KEYINPUT19), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n413), .B(new_n414), .C1(G146), .C2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n402), .A3(new_n384), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT82), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n420), .B(new_n422), .C1(new_n399), .C2(new_n402), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n412), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G478), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT15), .ZN(new_n428));
  INV_X1    g242(.A(G122), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT84), .B1(new_n429), .B2(G116), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n314), .A3(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT14), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(G116), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT14), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n430), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n434), .B1(new_n433), .B2(KEYINPUT14), .ZN(new_n440));
  OAI21_X1  g254(.A(G107), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n433), .A2(new_n210), .A3(new_n436), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n192), .A2(G128), .A3(new_n193), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(G128), .B2(new_n191), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G134), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n443), .B(new_n248), .C1(G128), .C2(new_n191), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n210), .B1(new_n433), .B2(new_n436), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n446), .B1(new_n442), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G134), .B1(new_n443), .B2(KEYINPUT13), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n191), .A2(G128), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n202), .B2(G128), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(KEYINPUT13), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT85), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n449), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n433), .A2(new_n210), .A3(new_n436), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT13), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n202), .A2(new_n459), .A3(G128), .ZN(new_n460));
  OAI211_X1 g274(.A(G134), .B(new_n460), .C1(new_n444), .C2(new_n459), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n458), .A2(new_n461), .A3(new_n462), .A4(new_n446), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n448), .A2(new_n455), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G217), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n298), .A2(new_n465), .A3(G953), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n464), .A2(KEYINPUT87), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT87), .B1(new_n464), .B2(new_n467), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n448), .A2(new_n455), .A3(new_n463), .A4(new_n466), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n428), .B1(new_n472), .B2(G902), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n464), .A2(new_n467), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n464), .A2(KEYINPUT87), .A3(new_n467), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n470), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n188), .C1(KEYINPUT15), .C2(new_n427), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(G234), .A2(G237), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(G952), .A3(new_n283), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(G902), .A3(G953), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT88), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT21), .B(G898), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n426), .A2(new_n480), .A3(new_n488), .ZN(new_n489));
  AND4_X1   g303(.A1(new_n300), .A2(new_n359), .A3(new_n361), .A4(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n363), .A2(new_n283), .A3(G210), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT27), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(G101), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n235), .A2(new_n274), .A3(new_n240), .ZN(new_n496));
  INV_X1    g310(.A(new_n332), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n248), .A2(G137), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n250), .A2(G134), .ZN(new_n499));
  OAI21_X1  g313(.A(G131), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n256), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n259), .B2(new_n260), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT28), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n237), .B1(new_n239), .B2(new_n229), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n257), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n332), .B1(new_n507), .B2(new_n502), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n495), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n496), .A2(KEYINPUT30), .A3(new_n503), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n507), .B2(new_n502), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n512), .A3(new_n332), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n510), .A2(new_n512), .A3(KEYINPUT66), .A4(new_n332), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n504), .A2(new_n495), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT67), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT67), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n504), .A2(new_n520), .A3(new_n495), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT31), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(KEYINPUT31), .A3(new_n522), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n509), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G472), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n188), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n491), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n509), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n517), .A2(KEYINPUT31), .A3(new_n522), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT31), .B1(new_n517), .B2(new_n522), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(KEYINPUT32), .A3(new_n528), .A4(new_n188), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n496), .A2(new_n503), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n332), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n505), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n495), .A2(KEYINPUT29), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n495), .B1(new_n517), .B2(new_n504), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n505), .A2(new_n508), .A3(new_n495), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT29), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n540), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G472), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n530), .A2(new_n535), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT68), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT22), .B(G137), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n318), .B2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n553), .B(new_n554), .C1(G119), .C2(new_n197), .ZN(new_n555));
  XNOR2_X1  g369(.A(G119), .B(G128), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT24), .B(G110), .Z(new_n557));
  AOI22_X1  g371(.A1(new_n555), .A2(G110), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n388), .B2(new_n389), .ZN(new_n559));
  OAI22_X1  g373(.A1(new_n555), .A2(G110), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n414), .A3(new_n382), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT69), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n559), .B2(new_n561), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n551), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n551), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n559), .A2(new_n561), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(KEYINPUT69), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n188), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(KEYINPUT70), .A2(KEYINPUT25), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n570), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n565), .A2(new_n188), .A3(new_n568), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(KEYINPUT70), .A2(KEYINPUT25), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n465), .B1(G234), .B2(new_n188), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n565), .A2(new_n568), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(G902), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n547), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n490), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  NOR2_X1   g396(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n527), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n583), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n534), .A2(new_n188), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n273), .A2(new_n289), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n285), .B1(new_n267), .B2(new_n272), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n588), .A2(new_n285), .B1(new_n589), .B2(new_n281), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n590), .A2(G469), .A3(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n296), .A2(new_n292), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n579), .B(new_n299), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n478), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n474), .A2(KEYINPUT33), .A3(new_n470), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n427), .A2(G902), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n596), .A2(KEYINPUT90), .A3(new_n597), .A4(new_n598), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n427), .B1(new_n472), .B2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n426), .ZN(new_n605));
  INV_X1    g419(.A(new_n301), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n345), .A2(new_n354), .ZN(new_n607));
  INV_X1    g421(.A(new_n355), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n345), .A2(new_n354), .A3(new_n355), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n488), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n594), .A2(new_n605), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  INV_X1    g430(.A(KEYINPUT92), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT91), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n425), .A2(new_n618), .B1(new_n411), .B2(G475), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n419), .A2(new_n402), .A3(new_n384), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n409), .B2(new_n401), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT20), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n422), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(KEYINPUT91), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n480), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n617), .B1(new_n626), .B2(new_n613), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n619), .A2(new_n625), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n358), .A2(new_n488), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT92), .A4(new_n480), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n594), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NAND2_X1  g447(.A1(new_n575), .A2(new_n576), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n566), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n567), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n578), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n587), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n490), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT93), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(G12));
  NOR2_X1   g458(.A1(new_n639), .A2(new_n358), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n547), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n482), .B(KEYINPUT94), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(new_n486), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n480), .A2(new_n619), .A3(new_n625), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT95), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n647), .A2(new_n300), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  NAND2_X1  g471(.A1(new_n609), .A2(new_n610), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT38), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n639), .A2(new_n301), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n426), .A2(new_n480), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n495), .B1(new_n537), .B2(new_n504), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n517), .B2(new_n522), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n665), .B2(G902), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n530), .A2(new_n535), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT96), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n663), .A2(KEYINPUT96), .A3(new_n667), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n651), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n300), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n300), .A2(KEYINPUT40), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n670), .A2(new_n671), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n238), .ZN(G45));
  NAND2_X1  g493(.A1(new_n602), .A2(new_n603), .ZN(new_n680));
  INV_X1    g494(.A(new_n597), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n478), .B2(new_n595), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT90), .B1(new_n682), .B2(new_n598), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n426), .B(new_n652), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n547), .A3(new_n300), .A4(new_n645), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  INV_X1    g501(.A(new_n299), .ZN(new_n688));
  OAI21_X1  g502(.A(G469), .B1(new_n590), .B2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(KEYINPUT97), .A3(new_n291), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT97), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n691), .B(G469), .C1(new_n590), .C2(G902), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n580), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n605), .A2(new_n613), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND2_X1  g512(.A1(new_n630), .A2(new_n627), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  AND2_X1   g515(.A1(new_n693), .A2(new_n489), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n647), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  OAI21_X1  g518(.A(G472), .B1(new_n527), .B2(G902), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n495), .B1(new_n505), .B2(new_n537), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n525), .B2(new_n526), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT98), .B1(new_n707), .B2(new_n529), .ZN(new_n708));
  OAI22_X1  g522(.A1(new_n532), .A2(new_n533), .B1(new_n495), .B2(new_n538), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT98), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n528), .A4(new_n188), .ZN(new_n711));
  AND4_X1   g525(.A1(new_n579), .A2(new_n705), .A3(new_n708), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT99), .ZN(new_n713));
  AND4_X1   g527(.A1(new_n611), .A2(new_n426), .A3(new_n480), .A4(new_n612), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n712), .A2(new_n713), .A3(new_n693), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n690), .A2(new_n692), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n714), .A3(new_n299), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n705), .A2(new_n708), .A3(new_n711), .A4(new_n579), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT99), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND2_X1  g535(.A1(new_n693), .A2(new_n611), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n705), .A2(new_n708), .A3(new_n711), .A4(new_n638), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n723), .A3(new_n684), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n303), .ZN(G27));
  NOR3_X1   g539(.A1(new_n356), .A2(new_n357), .A3(new_n606), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n297), .A2(new_n299), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n685), .A2(new_n547), .A3(new_n579), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  NAND4_X1  g547(.A1(new_n655), .A2(new_n547), .A3(new_n579), .A4(new_n727), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT101), .B(G134), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G36));
  AOI22_X1  g550(.A1(new_n623), .A2(new_n624), .B1(new_n411), .B2(G475), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n604), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(KEYINPUT104), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n604), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n639), .B1(new_n584), .B2(new_n586), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT106), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n745), .A2(new_n749), .A3(new_n746), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n741), .A2(KEYINPUT44), .A3(new_n743), .A4(new_n744), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT105), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n752), .A2(KEYINPUT105), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n726), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT107), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n726), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n752), .A2(KEYINPUT105), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n759), .B2(new_n753), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n748), .A2(new_n750), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n273), .A2(new_n289), .A3(new_n286), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n295), .B1(new_n273), .B2(new_n281), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n293), .B(KEYINPUT45), .C1(new_n294), .C2(new_n295), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(G469), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT46), .B1(new_n769), .B2(new_n292), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT102), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n292), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n291), .B(new_n774), .C1(new_n770), .C2(new_n771), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n299), .B(new_n672), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT103), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n757), .A2(new_n763), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  OAI21_X1  g594(.A(new_n299), .B1(new_n773), .B2(new_n775), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n547), .A2(new_n684), .A3(new_n579), .A4(new_n758), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  AND2_X1   g600(.A1(new_n728), .A2(new_n729), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n728), .A2(new_n731), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n723), .A2(new_n684), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n727), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n473), .A2(new_n479), .A3(new_n652), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n628), .A2(new_n638), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n297), .A2(new_n299), .A3(new_n726), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT110), .B1(new_n796), .B2(new_n547), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n619), .A2(new_n625), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n639), .A3(new_n792), .ZN(new_n799));
  AND4_X1   g613(.A1(KEYINPUT110), .A2(new_n799), .A3(new_n547), .A4(new_n727), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n734), .B(new_n791), .C1(new_n797), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n789), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n359), .A2(new_n361), .A3(new_n612), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n587), .A2(new_n803), .A3(new_n593), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n737), .A2(new_n480), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT109), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n737), .A2(new_n480), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n605), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n647), .A2(new_n702), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n490), .B1(new_n580), .B2(new_n640), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n580), .B(new_n693), .C1(new_n695), .C2(new_n699), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n720), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n693), .A2(new_n611), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n790), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n662), .A2(new_n358), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n651), .B(KEYINPUT111), .Z(new_n817));
  NOR2_X1   g631(.A1(new_n638), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n667), .A2(new_n300), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n656), .A2(new_n815), .A3(new_n686), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n685), .A2(new_n300), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n628), .A2(new_n654), .A3(new_n480), .A4(new_n652), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n653), .A2(KEYINPUT95), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n300), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n646), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n724), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n819), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n802), .A2(new_n813), .A3(new_n821), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n799), .A2(new_n547), .A3(new_n727), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n547), .A2(new_n727), .A3(new_n579), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n836), .A2(new_n655), .B1(new_n790), .B2(new_n727), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n732), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n720), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n821), .A4(new_n829), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n830), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(KEYINPUT112), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n830), .A2(new_n831), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT112), .B1(new_n830), .B2(new_n845), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n741), .A2(new_n649), .A3(new_n743), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(KEYINPUT114), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(KEYINPUT114), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n718), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n693), .A2(new_n606), .A3(new_n660), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n861), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n862), .A2(new_n863), .B1(new_n859), .B2(new_n860), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n716), .A2(new_n688), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n726), .B(new_n856), .C1(new_n783), .C2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT51), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n693), .A2(new_n726), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n854), .B2(new_n855), .ZN(new_n871));
  INV_X1    g685(.A(new_n723), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n579), .A2(new_n483), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n870), .A2(new_n667), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n604), .A2(new_n426), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n871), .A2(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n867), .A2(new_n876), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n864), .A2(new_n869), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n867), .A2(new_n868), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n879), .B(new_n880), .C1(new_n864), .C2(new_n877), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(new_n426), .A3(new_n604), .ZN(new_n882));
  INV_X1    g696(.A(G952), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT117), .B1(new_n883), .B2(G953), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n882), .B(new_n884), .C1(KEYINPUT117), .C2(G953), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n814), .B2(new_n856), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n871), .A2(new_n580), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT118), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n888), .B2(KEYINPUT48), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n887), .A2(KEYINPUT118), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n890), .A2(KEYINPUT48), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n889), .B1(new_n891), .B2(new_n888), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n878), .A2(new_n881), .A3(new_n892), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n852), .A2(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n579), .A2(new_n299), .A3(new_n301), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n660), .B1(KEYINPUT108), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n738), .B(new_n896), .C1(KEYINPUT108), .C2(new_n895), .ZN(new_n897));
  INV_X1    g711(.A(new_n667), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n716), .B(KEYINPUT49), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n894), .A2(new_n900), .ZN(G75));
  INV_X1    g715(.A(new_n842), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n188), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(G210), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n348), .A2(new_n353), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(new_n351), .Z(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n909), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n904), .B2(new_n905), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n283), .A2(G952), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(G51));
  XOR2_X1   g728(.A(new_n292), .B(KEYINPUT57), .Z(new_n915));
  NOR2_X1   g729(.A1(new_n902), .A2(new_n851), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n843), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n290), .B2(new_n287), .ZN(new_n918));
  OR3_X1    g732(.A1(new_n902), .A2(new_n188), .A3(new_n769), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n913), .B1(new_n918), .B2(new_n919), .ZN(G54));
  INV_X1    g734(.A(new_n913), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(new_n621), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(G60));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT59), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n682), .B1(new_n852), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n682), .B(new_n927), .C1(new_n916), .C2(new_n843), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n921), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G63));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  AND4_X1   g749(.A1(new_n932), .A2(new_n842), .A3(new_n636), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n832), .B2(new_n841), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n932), .B1(new_n937), .B2(new_n636), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT120), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n842), .A2(new_n636), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT119), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n932), .A3(new_n636), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n937), .A2(new_n577), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n913), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n936), .A2(new_n938), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT61), .B(new_n921), .C1(new_n937), .C2(new_n577), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT121), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n951), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT121), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n953), .B(new_n954), .C1(new_n936), .C2(new_n938), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n949), .A2(new_n956), .ZN(G66));
  INV_X1    g771(.A(G224), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n487), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n813), .B2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n907), .B1(G898), .B2(new_n283), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G69));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n778), .A2(new_n580), .A3(new_n816), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n827), .A2(new_n732), .A3(new_n734), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n964), .A2(new_n785), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(G953), .B1(new_n966), .B2(new_n779), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n283), .A2(G900), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n968), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n964), .A2(new_n785), .A3(new_n965), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n763), .A2(new_n778), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n757), .ZN(new_n973));
  OAI211_X1 g787(.A(KEYINPUT125), .B(new_n970), .C1(new_n973), .C2(G953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n510), .A2(new_n512), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(new_n418), .Z(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n969), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n678), .A2(new_n827), .ZN(new_n979));
  XOR2_X1   g793(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n678), .B(new_n827), .C1(KEYINPUT122), .C2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n836), .A2(new_n672), .A3(new_n809), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT123), .ZN(new_n985));
  AND4_X1   g799(.A1(new_n785), .A2(new_n981), .A3(new_n983), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(G953), .B1(new_n779), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT124), .B1(new_n987), .B2(new_n977), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n779), .A2(new_n986), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n283), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n991), .A3(new_n976), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n978), .A2(new_n988), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n992), .A2(new_n988), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n993), .B1(new_n995), .B2(new_n978), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n994), .A2(new_n996), .ZN(G72));
  INV_X1    g811(.A(new_n850), .ZN(new_n998));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n541), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n523), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n913), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1000), .B1(new_n989), .B2(new_n839), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n517), .A2(new_n504), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1007), .A2(new_n495), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1008), .A2(new_n495), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n973), .A2(new_n813), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n1000), .ZN(new_n1014));
  AOI211_X1 g828(.A(KEYINPUT127), .B(new_n1001), .C1(new_n973), .C2(new_n813), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1004), .A2(new_n1010), .A3(new_n1016), .ZN(G57));
endmodule


