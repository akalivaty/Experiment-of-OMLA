//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT17), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT92), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n206), .ZN(new_n208));
  OR2_X1    g007(.A1(G15gat), .A2(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G15gat), .A2(G22gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n205), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI211_X1 g011(.A(G8gat), .B(new_n207), .C1(new_n212), .C2(KEYINPUT92), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(KEYINPUT91), .A3(new_n211), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n211), .A2(KEYINPUT91), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n214), .A2(new_n215), .A3(G8gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n203), .B1(new_n217), .B2(KEYINPUT93), .ZN(new_n218));
  OR3_X1    g017(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n219), .A2(new_n220), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT15), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G50gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G43gat), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT15), .B1(new_n227), .B2(KEYINPUT89), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(new_n223), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT89), .ZN(new_n230));
  INV_X1    g029(.A(G43gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G50gat), .ZN(new_n232));
  AND4_X1   g031(.A1(new_n230), .A2(new_n227), .A3(new_n232), .A4(new_n222), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n221), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT90), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n221), .C1(new_n229), .C2(new_n233), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n225), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n218), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT93), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n238), .B2(KEYINPUT17), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n241), .A2(new_n217), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT18), .B(new_n202), .C1(new_n239), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n238), .A2(new_n218), .B1(new_n241), .B2(new_n217), .ZN(new_n245));
  INV_X1    g044(.A(new_n202), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n217), .B(new_n238), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n202), .B(KEYINPUT13), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n243), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  INV_X1    g052(.A(G197gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT11), .B(G169gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT12), .Z(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n251), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n251), .B2(new_n252), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT95), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G57gat), .B(G64gat), .Z(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G71gat), .A2(G78gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT94), .ZN(new_n270));
  NOR2_X1   g069(.A1(G71gat), .A2(G78gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT96), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n268), .A2(KEYINPUT96), .A3(new_n270), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n269), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n266), .A2(new_n267), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT97), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT21), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n217), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G183gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n286), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n277), .A2(new_n280), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT21), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n287), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n287), .B2(new_n288), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G155gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G231gat), .A2(G233gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  OR3_X1    g097(.A1(new_n293), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n293), .B2(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G85gat), .A2(G92gat), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n302), .A2(KEYINPUT99), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT7), .B1(new_n302), .B2(KEYINPUT99), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  NAND2_X1  g105(.A1(G99gat), .A2(G106gat), .ZN(new_n307));
  INV_X1    g106(.A(G85gat), .ZN(new_n308));
  INV_X1    g107(.A(G92gat), .ZN(new_n309));
  AOI22_X1  g108(.A1(KEYINPUT8), .A2(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT100), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n305), .B(new_n306), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G99gat), .B(G106gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT101), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n310), .B(new_n311), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n302), .A2(KEYINPUT99), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n304), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT101), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .A4(new_n315), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n317), .A2(new_n322), .B1(new_n316), .B2(new_n314), .ZN(new_n323));
  INV_X1    g122(.A(new_n238), .ZN(new_n324));
  OR3_X1    g123(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT17), .ZN(new_n325));
  XOR2_X1   g124(.A(G190gat), .B(G218gat), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(G232gat), .A2(G233gat), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n327), .A2(KEYINPUT102), .B1(KEYINPUT41), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n324), .B1(new_n323), .B2(KEYINPUT17), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n325), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n328), .A2(KEYINPUT41), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT98), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n333), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n325), .A2(new_n335), .A3(new_n329), .A4(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n327), .A2(KEYINPUT102), .ZN(new_n338));
  XOR2_X1   g137(.A(G134gat), .B(G162gat), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n337), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n317), .A2(new_n322), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT103), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n314), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n318), .A2(KEYINPUT103), .A3(new_n320), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n316), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n344), .A2(new_n277), .A3(new_n348), .A4(new_n280), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n349), .B(new_n350), .C1(new_n289), .C2(new_n323), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n289), .A2(KEYINPUT10), .A3(new_n323), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G230gat), .ZN(new_n354));
  INV_X1    g153(.A(G233gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n349), .B1(new_n289), .B2(new_n323), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n356), .ZN(new_n360));
  XNOR2_X1  g159(.A(G120gat), .B(G148gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G176gat), .B(G204gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n358), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n358), .B2(new_n360), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n301), .A2(new_n343), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G141gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(G148gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(G141gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT77), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  INV_X1    g175(.A(G155gat), .ZN(new_n377));
  INV_X1    g176(.A(G162gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n376), .B1(new_n379), .B2(KEYINPUT2), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(G141gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n371), .A2(G148gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n375), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  XNOR2_X1  g185(.A(G141gat), .B(G148gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n376), .B(new_n379), .C1(new_n387), .C2(KEYINPUT2), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n386), .B1(new_n385), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392));
  XNOR2_X1  g191(.A(G127gat), .B(G134gat), .ZN(new_n393));
  INV_X1    g192(.A(G120gat), .ZN(new_n394));
  INV_X1    g193(.A(G113gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT69), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G113gat), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n394), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n395), .A2(G120gat), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n392), .B(new_n393), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(G134gat), .A3(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(G127gat), .A2(G134gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G113gat), .B(G120gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n404), .B(new_n405), .C1(KEYINPUT1), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n370), .B1(new_n391), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(KEYINPUT70), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n401), .A2(new_n412), .A3(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n385), .A2(new_n388), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n408), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT78), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n417), .A2(new_n415), .A3(new_n418), .A4(new_n410), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n401), .A2(new_n385), .A3(new_n407), .A4(new_n388), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT78), .B1(new_n420), .B2(KEYINPUT4), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n409), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n415), .B(new_n408), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n424), .A2(new_n369), .ZN(new_n425));
  XOR2_X1   g224(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n414), .A2(new_n410), .A3(new_n415), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT80), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n420), .A2(new_n429), .A3(KEYINPUT4), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n420), .A2(KEYINPUT4), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT80), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n426), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n391), .A2(new_n408), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n433), .A2(new_n369), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(new_n308), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT0), .B(G57gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n427), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT81), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n427), .B2(new_n436), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n448), .A3(new_n443), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT82), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(KEYINPUT6), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n445), .A2(new_n453), .A3(new_n447), .A4(new_n449), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G211gat), .B(G218gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT74), .ZN(new_n457));
  INV_X1    g256(.A(G218gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n291), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G204gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n254), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(G197gat), .A2(G204gat), .ZN(new_n462));
  OAI22_X1  g261(.A1(KEYINPUT22), .A2(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n457), .A2(new_n463), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT75), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n457), .A2(new_n463), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n386), .B1(new_n470), .B2(KEYINPUT29), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n385), .A2(new_n388), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n474));
  INV_X1    g273(.A(G228gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(new_n355), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n466), .B(new_n469), .C1(KEYINPUT29), .C2(new_n389), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n473), .A2(new_n474), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n466), .A2(new_n469), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT29), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT3), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n476), .B(new_n477), .C1(new_n481), .C2(new_n415), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT83), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n464), .A2(new_n465), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n386), .B1(new_n484), .B2(KEYINPUT29), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n472), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n477), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n475), .B2(new_n355), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n478), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G50gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(G22gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n493), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n496), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n478), .A2(new_n488), .A3(new_n483), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT64), .ZN(new_n501));
  INV_X1    g300(.A(G190gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n284), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G183gat), .A2(G190gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT24), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n503), .A2(new_n506), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G169gat), .A2(G176gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT23), .ZN(new_n511));
  INV_X1    g310(.A(G169gat), .ZN(new_n512));
  INV_X1    g311(.A(G176gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT23), .B(new_n512), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n509), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n284), .A2(new_n502), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT23), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n523), .A2(new_n515), .A3(KEYINPUT25), .A4(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n512), .A2(KEYINPUT23), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n513), .A2(new_n528), .B1(new_n511), .B2(new_n514), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(KEYINPUT66), .A3(KEYINPUT25), .A4(new_n523), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n521), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  OR4_X1    g330(.A1(KEYINPUT67), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT67), .B1(new_n514), .B2(KEYINPUT26), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n514), .A2(KEYINPUT26), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n510), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G183gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT28), .A3(new_n502), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT28), .B1(new_n536), .B2(new_n502), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n535), .B(new_n504), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n414), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n531), .A2(new_n411), .A3(new_n540), .A4(new_n413), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G227gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n355), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT34), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT34), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G15gat), .B(G43gat), .Z(new_n554));
  XOR2_X1   g353(.A(G71gat), .B(G99gat), .Z(new_n555));
  XOR2_X1   g354(.A(new_n554), .B(new_n555), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n546), .A3(new_n543), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT33), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n560), .A2(KEYINPUT71), .B1(KEYINPUT32), .B2(new_n558), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n557), .A2(new_n559), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n553), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n558), .A2(new_n559), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(KEYINPUT71), .A3(new_n556), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n564), .A3(new_n556), .ZN(new_n571));
  INV_X1    g370(.A(new_n563), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n573), .A3(new_n552), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n500), .A2(new_n566), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n541), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n531), .A2(new_n540), .A3(KEYINPUT76), .ZN(new_n578));
  AND2_X1   g377(.A1(G226gat), .A2(G233gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(KEYINPUT29), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n531), .A2(new_n540), .A3(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n479), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n577), .A2(new_n578), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n579), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n541), .A2(new_n580), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n470), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G8gat), .B(G36gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(G64gat), .B(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT30), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n592), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT30), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n589), .B2(new_n592), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n455), .A2(new_n575), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT73), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n566), .A2(new_n574), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n570), .A2(new_n573), .A3(KEYINPUT73), .A4(new_n552), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n500), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  MUX2_X1   g407(.A(new_n444), .B(new_n443), .S(new_n446), .Z(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(KEYINPUT35), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n599), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n455), .A2(new_n599), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n603), .A2(new_n604), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n566), .A2(new_n574), .A3(KEYINPUT36), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n589), .A2(KEYINPUT37), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n588), .A2(new_n584), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n592), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n593), .B1(new_n622), .B2(KEYINPUT38), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n586), .A2(new_n479), .A3(new_n587), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n583), .A2(new_n470), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT37), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n626), .A3(new_n592), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n623), .B(new_n609), .C1(KEYINPUT38), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n433), .A2(new_n435), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n370), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT85), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(KEYINPUT85), .A3(new_n370), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n440), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n424), .B2(new_n369), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT86), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n598), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n633), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT85), .B1(new_n629), .B2(new_n370), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n635), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(new_n441), .A3(new_n638), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT86), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n640), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n447), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n500), .B(new_n628), .C1(new_n641), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n614), .A2(new_n618), .A3(new_n649), .ZN(new_n650));
  AOI211_X1 g449(.A(new_n263), .B(new_n368), .C1(new_n612), .C2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n455), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g453(.A(KEYINPUT16), .B(G8gat), .Z(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n598), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT104), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n651), .A2(new_n598), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(G8gat), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n659), .B(new_n661), .C1(new_n657), .C2(new_n656), .ZN(G1325gat));
  AOI21_X1  g461(.A(G15gat), .B1(new_n651), .B2(new_n605), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n618), .A2(KEYINPUT105), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n616), .A2(new_n665), .A3(new_n617), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT106), .Z(new_n670));
  AOI21_X1  g469(.A(new_n663), .B1(new_n651), .B2(new_n670), .ZN(G1326gat));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n607), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT43), .B(G22gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  AOI21_X1  g473(.A(new_n343), .B1(new_n612), .B2(new_n650), .ZN(new_n675));
  INV_X1    g474(.A(new_n367), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n301), .A2(new_n263), .A3(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(G29gat), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n678), .A2(KEYINPUT108), .A3(new_n679), .A4(new_n652), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n675), .A2(new_n679), .A3(new_n677), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n455), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n614), .A2(new_n649), .A3(new_n667), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n612), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n690), .A3(new_n342), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n690), .B2(new_n675), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n677), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n455), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n680), .A2(new_n685), .A3(new_n683), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n687), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT109), .ZN(G1328gat));
  INV_X1    g496(.A(new_n678), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(G36gat), .A3(new_n599), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  OAI21_X1  g499(.A(G36gat), .B1(new_n693), .B2(new_n599), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(G1329gat));
  OAI21_X1  g501(.A(new_n231), .B1(new_n698), .B2(new_n606), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n692), .A2(G43gat), .A3(new_n668), .A4(new_n677), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g505(.A(new_n226), .B1(new_n698), .B2(new_n500), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n607), .A2(G50gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n693), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g509(.A(new_n301), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n711), .B(new_n342), .C1(new_n612), .C2(new_n688), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n262), .A2(new_n367), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n455), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT110), .B(G57gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1332gat));
  NOR2_X1   g516(.A1(new_n714), .A2(new_n599), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  AND2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n718), .B2(new_n719), .ZN(G1333gat));
  INV_X1    g521(.A(new_n714), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n723), .A2(G71gat), .A3(new_n668), .ZN(new_n724));
  AOI21_X1  g523(.A(G71gat), .B1(new_n723), .B2(new_n605), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n607), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  AOI211_X1 g528(.A(new_n262), .B(new_n343), .C1(new_n612), .C2(new_n688), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT51), .B1(new_n730), .B2(new_n711), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(KEYINPUT51), .A3(new_n711), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n733), .B2(new_n732), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n455), .A2(G85gat), .A3(new_n367), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT113), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n612), .A2(new_n650), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n690), .B1(new_n739), .B2(new_n342), .ZN(new_n740));
  AOI211_X1 g539(.A(KEYINPUT44), .B(new_n343), .C1(new_n612), .C2(new_n688), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n711), .B(new_n713), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT111), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n692), .A2(new_n744), .A3(new_n711), .A4(new_n713), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n455), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n736), .A2(new_n738), .B1(new_n746), .B2(new_n308), .ZN(G1336gat));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n745), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n309), .B1(new_n748), .B2(new_n598), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n676), .A2(new_n309), .A3(new_n598), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT114), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n689), .A2(new_n263), .A3(new_n342), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n752), .A2(new_n753), .A3(new_n301), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n751), .B1(new_n731), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT115), .B(new_n751), .C1(new_n731), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n735), .B(new_n751), .C1(new_n733), .C2(new_n732), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  OAI21_X1  g561(.A(G92gat), .B1(new_n742), .B2(new_n599), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(G1337gat));
  INV_X1    g564(.A(G99gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n676), .A2(new_n605), .A3(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT116), .Z(new_n768));
  AOI21_X1  g567(.A(new_n667), .B1(new_n743), .B2(new_n745), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n736), .A2(new_n768), .B1(new_n769), .B2(new_n766), .ZN(G1338gat));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  OAI21_X1  g570(.A(G106gat), .B1(new_n742), .B2(new_n500), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n500), .A2(new_n367), .A3(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n771), .B(new_n772), .C1(new_n736), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n732), .B2(new_n734), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n748), .A2(new_n607), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(G106gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n778), .B2(new_n771), .ZN(G1339gat));
  NAND3_X1  g578(.A1(new_n351), .A2(new_n356), .A3(new_n352), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n351), .A2(KEYINPUT117), .A3(new_n356), .A4(new_n352), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n782), .A2(new_n358), .A3(KEYINPUT54), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n356), .B1(new_n351), .B2(new_n352), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n364), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n365), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n784), .A2(KEYINPUT55), .A3(new_n787), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n784), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n787), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n790), .A2(new_n793), .A3(new_n262), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n245), .A2(new_n246), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n249), .B2(new_n248), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n257), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n251), .B2(new_n258), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n367), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n343), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n790), .A2(new_n793), .A3(new_n342), .A4(new_n794), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n804), .A2(new_n799), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n342), .B1(new_n795), .B2(new_n800), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n804), .A2(new_n799), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT119), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n711), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n301), .A2(new_n263), .A3(new_n343), .A4(new_n367), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n455), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n599), .A3(new_n608), .ZN(new_n813));
  OAI21_X1  g612(.A(G113gat), .B1(new_n813), .B2(new_n263), .ZN(new_n814));
  INV_X1    g613(.A(new_n811), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n807), .A2(new_n808), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n301), .B1(new_n816), .B2(new_n803), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n817), .B2(new_n809), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n818), .A2(new_n455), .A3(new_n598), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n575), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n820), .A2(KEYINPUT120), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n396), .A2(new_n398), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(KEYINPUT120), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n814), .B1(new_n824), .B2(new_n263), .ZN(G1340gat));
  OAI21_X1  g624(.A(G120gat), .B1(new_n813), .B2(new_n367), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n676), .A2(new_n394), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(G1341gat));
  NOR2_X1   g628(.A1(new_n820), .A2(new_n711), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n402), .B2(new_n403), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n301), .A2(new_n402), .A3(new_n403), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n813), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT121), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n831), .A2(new_n834), .ZN(G1342gat));
  NOR3_X1   g634(.A1(new_n820), .A2(G134gat), .A3(new_n343), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n813), .B2(new_n343), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  NOR2_X1   g640(.A1(new_n668), .A2(new_n500), .ZN(new_n842));
  AND4_X1   g641(.A1(new_n371), .A2(new_n812), .A3(new_n599), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n810), .A2(new_n811), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n607), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n667), .A2(new_n652), .A3(new_n599), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n811), .B1(new_n816), .B2(new_n301), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n607), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(KEYINPUT57), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(new_n850), .A3(new_n262), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n262), .A2(new_n843), .B1(new_n851), .B2(G141gat), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT122), .B1(new_n851), .B2(G141gat), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n852), .A2(KEYINPUT58), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n843), .A2(new_n262), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(G141gat), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(KEYINPUT58), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n854), .A2(new_n859), .ZN(G1344gat));
  NAND4_X1  g659(.A1(new_n819), .A2(new_n373), .A3(new_n676), .A4(new_n842), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT57), .B1(new_n818), .B2(new_n500), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n847), .B(KEYINPUT123), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n799), .B1(new_n804), .B2(KEYINPUT124), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(KEYINPUT124), .B2(new_n804), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n301), .B1(new_n866), .B2(new_n802), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n845), .B(new_n607), .C1(new_n867), .C2(new_n815), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n863), .A2(new_n676), .A3(new_n864), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n373), .B1(new_n869), .B2(KEYINPUT125), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n844), .A2(new_n607), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n802), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n711), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n873), .B2(new_n811), .ZN(new_n874));
  AOI22_X1  g673(.A1(KEYINPUT57), .A2(new_n871), .B1(new_n874), .B2(new_n607), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n676), .A4(new_n864), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n862), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n846), .A2(new_n850), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n373), .C1(new_n879), .C2(new_n676), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n861), .B1(new_n878), .B2(new_n880), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n819), .A2(new_n842), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT126), .B1(new_n882), .B2(new_n711), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n819), .A2(new_n884), .A3(new_n301), .A4(new_n842), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n377), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n879), .A2(G155gat), .A3(new_n301), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(G1346gat));
  OAI21_X1  g687(.A(new_n378), .B1(new_n882), .B2(new_n343), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n879), .A2(G162gat), .A3(new_n342), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n818), .A2(new_n652), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n598), .A3(new_n575), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n512), .A3(new_n262), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n652), .A2(new_n599), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n844), .A2(new_n608), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n897), .A2(new_n262), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n512), .B2(new_n898), .ZN(G1348gat));
  AOI21_X1  g698(.A(G176gat), .B1(new_n894), .B2(new_n676), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n367), .A2(new_n517), .A3(new_n516), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n897), .B2(new_n901), .ZN(G1349gat));
  INV_X1    g701(.A(new_n536), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n893), .A2(new_n903), .A3(new_n711), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n284), .B1(new_n897), .B2(new_n301), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n904), .A2(KEYINPUT60), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT60), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1350gat));
  AOI21_X1  g707(.A(new_n502), .B1(new_n897), .B2(new_n342), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT61), .Z(new_n910));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n502), .A3(new_n342), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1351gat));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n667), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n875), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n916), .B2(new_n263), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n875), .A2(KEYINPUT127), .A3(new_n262), .A4(new_n915), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(G197gat), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n892), .A2(new_n842), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n920), .A2(new_n598), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n254), .A3(new_n262), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(G1352gat));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n460), .A3(new_n598), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n924), .A2(KEYINPUT62), .A3(new_n367), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n875), .A2(new_n676), .A3(new_n915), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G204gat), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT62), .B1(new_n924), .B2(new_n367), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n921), .A2(new_n291), .A3(new_n301), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n875), .A2(new_n301), .A3(new_n915), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n931), .B2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1354gat));
  NAND3_X1  g734(.A1(new_n921), .A2(new_n458), .A3(new_n342), .ZN(new_n936));
  OAI21_X1  g735(.A(G218gat), .B1(new_n916), .B2(new_n343), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


