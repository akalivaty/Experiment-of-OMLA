//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT66), .Z(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n212));
  AND3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n207), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT67), .ZN(new_n217));
  INV_X1    g0017(.A(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n207), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G20), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n203), .A2(G50), .ZN(new_n227));
  OAI22_X1  g0027(.A1(new_n214), .A2(new_n215), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n217), .A2(new_n222), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n241), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  AND2_X1   g0050(.A1(new_n250), .A2(G274), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n250), .A2(new_n253), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n258), .A2(G226), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G222), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n266), .B1(new_n267), .B2(new_n264), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n250), .ZN(new_n271));
  AOI211_X1 g0071(.A(new_n256), .B(new_n259), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n272), .A2(G169), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n223), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n277), .B1(new_n252), .B2(G20), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n278), .B2(G50), .ZN(new_n279));
  OAI21_X1  g0079(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT68), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT8), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT69), .B1(new_n201), .B2(KEYINPUT8), .ZN(new_n287));
  OR3_X1    g0087(.A1(new_n201), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n284), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n277), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n279), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n272), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n273), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n278), .A2(G77), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT8), .B(G58), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n300), .A2(new_n283), .B1(new_n290), .B2(new_n267), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT15), .B(G87), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n292), .B2(new_n303), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n299), .B1(G77), .B2(new_n274), .C1(new_n304), .C2(new_n294), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT70), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n256), .B1(G244), .B2(new_n258), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n264), .A2(G232), .A3(new_n265), .ZN(new_n308));
  INV_X1    g0108(.A(G107), .ZN(new_n309));
  INV_X1    g0109(.A(G238), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n308), .B1(new_n309), .B2(new_n264), .C1(new_n268), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n271), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n306), .B(new_n314), .C1(new_n315), .C2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n305), .C1(G179), .C2(new_n313), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g0120(.A(new_n295), .B(KEYINPUT71), .Z(new_n321));
  INV_X1    g0121(.A(KEYINPUT72), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT9), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n295), .B(KEYINPUT71), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT9), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT72), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n272), .A2(G190), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n272), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n325), .B2(new_n324), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT10), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n327), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n327), .B2(new_n331), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n298), .B(new_n320), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n203), .B1(new_n285), .B2(new_n202), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT78), .A3(G20), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n282), .A2(G159), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT16), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT78), .B1(new_n336), .B2(G20), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT76), .ZN(new_n343));
  AND2_X1   g0143(.A1(KEYINPUT3), .A2(G33), .ZN(new_n344));
  NOR2_X1   g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n262), .A2(KEYINPUT76), .A3(new_n263), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n290), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR4_X1   g0150(.A1(new_n344), .A2(new_n345), .A3(new_n349), .A4(G20), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT77), .B1(new_n353), .B2(G68), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n348), .B2(new_n349), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT77), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n355), .A2(new_n356), .A3(new_n202), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n342), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n341), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(new_n338), .A3(new_n337), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n344), .A2(new_n345), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT7), .B1(new_n361), .B2(new_n290), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n202), .B1(new_n363), .B2(new_n352), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n340), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(new_n365), .A3(new_n277), .ZN(new_n366));
  INV_X1    g0166(.A(new_n274), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n289), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n278), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n289), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n255), .B1(new_n231), .B2(new_n257), .ZN(new_n372));
  MUX2_X1   g0172(.A(G223), .B(G226), .S(G1698), .Z(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n264), .B1(G33), .B2(G87), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n250), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(KEYINPUT79), .A3(new_n315), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT79), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n255), .B1(new_n231), .B2(new_n257), .C1(new_n374), .C2(new_n250), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n329), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(G190), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n377), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n366), .A2(new_n371), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT17), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n353), .A2(KEYINPUT77), .A3(G68), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n356), .B1(new_n355), .B2(new_n202), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n294), .B1(new_n387), .B2(new_n342), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n370), .B1(new_n388), .B2(new_n365), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n376), .A2(G179), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n379), .A2(G169), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT18), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n366), .B2(new_n371), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n366), .A2(new_n371), .A3(new_n382), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n384), .A2(new_n394), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT75), .ZN(new_n402));
  OAI21_X1  g0202(.A(G238), .B1(new_n257), .B2(KEYINPUT74), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT74), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n250), .B2(new_n253), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n255), .B(new_n402), .C1(new_n403), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n231), .A2(G1698), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n407), .B1(G226), .B2(G1698), .C1(new_n344), .C2(new_n345), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n250), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(KEYINPUT73), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT73), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n412), .B(new_n250), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n406), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n255), .B1(new_n403), .B2(new_n405), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n415), .A2(KEYINPUT75), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT13), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n410), .B(KEYINPUT73), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(KEYINPUT75), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .A4(new_n406), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT14), .B1(new_n422), .B2(new_n317), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(G179), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n417), .A2(new_n421), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(G169), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT12), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n367), .B2(new_n202), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n274), .A2(KEYINPUT12), .A3(G68), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n369), .A2(new_n202), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n267), .B2(new_n291), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n434), .A2(KEYINPUT11), .A3(new_n277), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT11), .B1(new_n434), .B2(new_n277), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n432), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n417), .A2(new_n421), .A3(G190), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n437), .B(new_n440), .C1(new_n422), .C2(new_n329), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n335), .A2(new_n401), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G264), .A3(new_n250), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G250), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G1698), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n344), .B2(new_n345), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT85), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G294), .ZN(new_n456));
  OAI211_X1 g0256(.A(G257), .B(G1698), .C1(new_n344), .C2(new_n345), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT85), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n453), .B(new_n458), .C1(new_n345), .C2(new_n344), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n455), .A2(new_n456), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n451), .B1(new_n460), .B2(new_n271), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(G274), .A3(new_n250), .A4(new_n446), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n461), .A2(new_n315), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(G200), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n290), .B2(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n309), .A2(KEYINPUT23), .A3(G20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n261), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n290), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n290), .B(G87), .C1(new_n344), .C2(new_n345), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT22), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n264), .A2(new_n477), .A3(new_n290), .A4(G87), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT24), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI211_X1 g0281(.A(KEYINPUT24), .B(new_n474), .C1(new_n476), .C2(new_n478), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n277), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n252), .A2(G33), .ZN(new_n484));
  AND4_X1   g0284(.A1(new_n223), .A2(new_n274), .A3(new_n276), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n367), .A2(KEYINPUT25), .A3(new_n309), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT25), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n274), .B2(G107), .ZN(new_n488));
  AOI22_X1  g0288(.A1(G107), .A2(new_n485), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT87), .B1(new_n466), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n461), .A2(new_n315), .A3(new_n463), .ZN(new_n492));
  INV_X1    g0292(.A(new_n463), .ZN(new_n493));
  AOI211_X1 g0293(.A(new_n493), .B(new_n451), .C1(new_n460), .C2(new_n271), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n494), .B2(G200), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT87), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n483), .A4(new_n489), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT86), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n460), .A2(new_n271), .ZN(new_n500));
  AND4_X1   g0300(.A1(G179), .A2(new_n500), .A3(new_n450), .A4(new_n463), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n317), .B1(new_n461), .B2(new_n463), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n461), .A2(G179), .A3(new_n463), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(KEYINPUT86), .C1(new_n494), .C2(new_n317), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n490), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT81), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT6), .ZN(new_n509));
  AND2_X1   g0309(.A1(G97), .A2(G107), .ZN(new_n510));
  NOR2_X1   g0310(.A1(G97), .A2(G107), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT6), .A2(G97), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT80), .B1(new_n513), .B2(G107), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(new_n309), .A3(KEYINPUT6), .A4(G97), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n518));
  OAI21_X1  g0318(.A(G107), .B1(new_n362), .B2(new_n351), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n277), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n274), .A2(G97), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n485), .B2(G97), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n508), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n294), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  INV_X1    g0325(.A(new_n523), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n525), .A2(KEYINPUT81), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G250), .A2(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(KEYINPUT4), .A2(G244), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(G1698), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n264), .A2(new_n531), .B1(G33), .B2(G283), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(new_n265), .C1(new_n344), .C2(new_n345), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n271), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT82), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n449), .A2(G257), .A3(new_n250), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n463), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n250), .B1(new_n532), .B2(new_n535), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT82), .B1(new_n543), .B2(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(G190), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(G200), .B1(new_n543), .B2(new_n540), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n544), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n543), .A2(new_n540), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n548), .A2(new_n317), .B1(new_n296), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n521), .A2(new_n523), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n528), .A2(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n274), .A2(G116), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n485), .B2(G116), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n294), .B1(G20), .B2(new_n471), .ZN(new_n555));
  AOI21_X1  g0355(.A(G20), .B1(G33), .B2(G283), .ZN(new_n556));
  INV_X1    g0356(.A(G97), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(G33), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT83), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n555), .B(KEYINPUT20), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n558), .B(new_n559), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT20), .B1(new_n564), .B2(new_n555), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n554), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n449), .A2(G270), .A3(new_n250), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n567), .A2(new_n463), .ZN(new_n568));
  OAI211_X1 g0368(.A(G264), .B(G1698), .C1(new_n344), .C2(new_n345), .ZN(new_n569));
  OAI211_X1 g0369(.A(G257), .B(new_n265), .C1(new_n344), .C2(new_n345), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n264), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n271), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n317), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT21), .B1(new_n566), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n567), .A2(new_n463), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n271), .B2(new_n572), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n574), .A2(KEYINPUT21), .B1(new_n577), .B2(G179), .ZN(new_n578));
  INV_X1    g0378(.A(new_n554), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n564), .A2(new_n555), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n579), .B1(new_n582), .B2(new_n562), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT84), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT84), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n577), .A2(new_n586), .A3(new_n317), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n568), .A2(new_n573), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(new_n296), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n585), .B(new_n566), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n575), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n566), .B1(G200), .B2(new_n588), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n315), .B2(new_n588), .ZN(new_n593));
  OAI211_X1 g0393(.A(G244), .B(G1698), .C1(new_n344), .C2(new_n345), .ZN(new_n594));
  OAI211_X1 g0394(.A(G238), .B(new_n265), .C1(new_n344), .C2(new_n345), .ZN(new_n595));
  INV_X1    g0395(.A(new_n472), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n271), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n252), .A2(G45), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G250), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n251), .A2(new_n446), .B1(new_n601), .B2(new_n250), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n290), .B1(new_n409), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(G87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n511), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n290), .B(G68), .C1(new_n344), .C2(new_n345), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n605), .B1(new_n291), .B2(new_n557), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n277), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n302), .A2(new_n367), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n485), .A2(G87), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n598), .A2(G190), .A3(new_n602), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n604), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n485), .A2(new_n303), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n598), .A2(new_n296), .A3(new_n602), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n250), .A2(G274), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n622), .A2(new_n599), .B1(new_n271), .B2(new_n600), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n271), .B2(new_n597), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n620), .B(new_n621), .C1(new_n624), .C2(G169), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n552), .A2(new_n591), .A3(new_n593), .A4(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n444), .A2(new_n507), .A3(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n298), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n398), .B(KEYINPUT17), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n441), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n439), .B1(new_n632), .B2(new_n319), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT91), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT90), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n366), .A2(new_n371), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n396), .B1(new_n638), .B2(new_n392), .ZN(new_n639));
  AOI211_X1 g0439(.A(KEYINPUT18), .B(new_n393), .C1(new_n366), .C2(new_n371), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n397), .A2(new_n394), .A3(KEYINPUT90), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n333), .A2(new_n334), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n629), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n578), .A2(new_n583), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n575), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n490), .B1(new_n502), .B2(new_n501), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n618), .A2(KEYINPUT88), .A3(new_n625), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT88), .B1(new_n618), .B2(new_n625), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n650), .A2(new_n498), .A3(new_n552), .A4(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n538), .B1(new_n537), .B2(new_n541), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n543), .A2(new_n540), .A3(KEYINPUT82), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n317), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n549), .A2(new_n296), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT89), .B1(new_n528), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n521), .A2(new_n508), .A3(new_n523), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT81), .B1(new_n525), .B2(new_n526), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n550), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n660), .A2(new_n653), .A3(new_n661), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n626), .A2(new_n550), .A3(new_n551), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT26), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n654), .A2(new_n625), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n443), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n646), .A2(new_n671), .ZN(G369));
  AND2_X1   g0472(.A1(new_n591), .A2(new_n593), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n252), .A2(new_n290), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n566), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n648), .B2(new_n680), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n490), .A2(new_n679), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT92), .Z(new_n685));
  INV_X1    g0485(.A(new_n679), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n685), .A2(new_n507), .B1(new_n506), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n685), .A2(new_n507), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n591), .A2(new_n679), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n679), .B(KEYINPUT93), .Z(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n649), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n688), .A2(new_n695), .ZN(G399));
  NOR2_X1   g0496(.A1(new_n219), .A2(G41), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n511), .A2(new_n607), .A3(new_n471), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n697), .A2(new_n252), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n227), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n697), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  NAND4_X1  g0502(.A1(new_n660), .A2(new_n653), .A3(KEYINPUT26), .A4(new_n666), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n668), .A2(new_n661), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n584), .A2(new_n590), .ZN(new_n706));
  INV_X1    g0506(.A(new_n575), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n506), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n498), .A3(new_n552), .A4(new_n653), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n709), .A3(new_n625), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n710), .A2(KEYINPUT98), .A3(new_n686), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT98), .B1(new_n710), .B2(new_n686), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT29), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n670), .A2(new_n692), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n461), .A2(new_n624), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n588), .B2(new_n296), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n577), .A2(KEYINPUT94), .A3(G179), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n548), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT30), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n494), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n549), .A2(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n588), .A3(new_n603), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n717), .B1(new_n724), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n723), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n729), .B2(new_n548), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n732), .A2(new_n734), .A3(KEYINPUT96), .A4(new_n727), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n731), .A2(new_n679), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n503), .A2(new_n490), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n739), .A2(new_n505), .B1(new_n491), .B2(new_n497), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n528), .A2(new_n547), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n550), .A2(new_n551), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n741), .A2(new_n742), .A3(new_n626), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n673), .A2(new_n740), .A3(new_n743), .A4(new_n692), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n692), .A2(new_n737), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n724), .B2(new_n730), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(KEYINPUT95), .B(new_n745), .C1(new_n724), .C2(new_n730), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n738), .A2(new_n744), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n713), .A2(new_n716), .B1(G330), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n702), .B1(new_n751), .B2(G1), .ZN(G364));
  AOI21_X1  g0552(.A(new_n223), .B1(G20), .B2(new_n317), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n290), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n315), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n309), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n290), .A2(new_n296), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(G190), .A3(new_n329), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n202), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n755), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G159), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT103), .B(KEYINPUT32), .Z(new_n767));
  AOI211_X1 g0567(.A(new_n757), .B(new_n762), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n758), .A2(new_n763), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n329), .A2(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n759), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n264), .B1(new_n267), .B2(new_n769), .C1(new_n772), .C2(new_n285), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n607), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n766), .A2(new_n767), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(KEYINPUT102), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(KEYINPUT102), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(G20), .B1(new_n770), .B2(G179), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT104), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n782), .A2(G50), .B1(new_n788), .B2(G97), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n768), .A2(new_n777), .A3(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n782), .A2(G326), .B1(new_n788), .B2(G294), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  INV_X1    g0592(.A(G329), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n769), .A2(new_n792), .B1(new_n764), .B2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n264), .B(new_n794), .C1(G322), .C2(new_n771), .ZN(new_n795));
  INV_X1    g0595(.A(new_n774), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G303), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  INV_X1    g0598(.A(new_n756), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n760), .A2(new_n798), .B1(G283), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n791), .A2(new_n795), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n754), .B1(new_n790), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n753), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n220), .A2(new_n264), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT100), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n809), .A2(G355), .B1(new_n471), .B2(new_n219), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n346), .A2(new_n347), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n219), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT101), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n700), .A2(new_n445), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n445), .C2(new_n247), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n807), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n218), .A2(G20), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n252), .B1(new_n817), .B2(G45), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n697), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n802), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n805), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n682), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT105), .Z(new_n825));
  OR2_X1    g0625(.A1(new_n682), .A2(G330), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n683), .A2(new_n820), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n305), .A2(new_n679), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n316), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n319), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n319), .A2(new_n679), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n714), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n750), .A2(G330), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n820), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n753), .A2(new_n803), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n821), .B1(new_n267), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT106), .B(G143), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n769), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n771), .A2(new_n843), .B1(new_n844), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n281), .B2(new_n761), .C1(new_n781), .C2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT34), .ZN(new_n848));
  INV_X1    g0648(.A(new_n811), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G132), .B2(new_n765), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n850), .B1(new_n242), .B2(new_n774), .C1(new_n202), .C2(new_n756), .ZN(new_n851));
  INV_X1    g0651(.A(new_n285), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(new_n852), .B2(new_n788), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n799), .A2(G87), .ZN(new_n854));
  INV_X1    g0654(.A(G283), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n854), .B1(new_n309), .B2(new_n774), .C1(new_n761), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n361), .B1(new_n764), .B2(new_n792), .ZN(new_n857));
  INV_X1    g0657(.A(G294), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n772), .A2(new_n858), .B1(new_n769), .B2(new_n471), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n782), .A2(G303), .B1(new_n788), .B2(G97), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n848), .A2(new_n853), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n835), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n841), .B1(new_n754), .B2(new_n862), .C1(new_n863), .C2(new_n804), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n839), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n817), .A2(new_n252), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n713), .A2(new_n443), .A3(new_n716), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT110), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT110), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n713), .A2(new_n870), .A3(new_n443), .A4(new_n716), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n872), .A2(new_n646), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n354), .A2(new_n357), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n340), .B1(new_n874), .B2(new_n360), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n370), .B1(new_n875), .B2(new_n388), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n398), .B1(new_n876), .B2(new_n677), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n393), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n677), .B1(new_n366), .B2(new_n371), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n383), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(new_n395), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n876), .A2(new_n677), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n401), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n885), .A2(new_n887), .A3(KEYINPUT38), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n885), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n428), .A2(new_n438), .A3(new_n686), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n641), .A2(new_n630), .A3(new_n642), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n880), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n398), .B(KEYINPUT90), .C1(new_n389), .C2(new_n677), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n883), .A2(new_n881), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n398), .B1(new_n389), .B2(new_n677), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n898), .A2(KEYINPUT90), .A3(new_n882), .A4(new_n395), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(new_n888), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n891), .B(new_n893), .C1(KEYINPUT39), .C2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n834), .B1(new_n714), .B2(new_n835), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n441), .A2(new_n423), .A3(new_n424), .A4(new_n427), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n437), .A2(new_n686), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT109), .ZN(new_n908));
  INV_X1    g0708(.A(new_n906), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n439), .A2(new_n441), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT109), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(new_n911), .A3(new_n906), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(new_n890), .ZN(new_n915));
  INV_X1    g0715(.A(new_n677), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n643), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n903), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n873), .B(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(G330), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n731), .A2(new_n735), .A3(KEYINPUT31), .A4(new_n679), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n738), .A2(new_n744), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n913), .A2(new_n923), .A3(new_n863), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n924), .B(KEYINPUT40), .C1(new_n888), .C2(new_n901), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n913), .A2(new_n923), .A3(new_n863), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n890), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n443), .A2(new_n923), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n921), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n867), .B1(new_n920), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n920), .B2(new_n933), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n267), .B(new_n227), .C1(new_n852), .C2(G68), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n243), .B(KEYINPUT107), .ZN(new_n937));
  OAI211_X1 g0737(.A(G1), .B(new_n218), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT108), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT36), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n941), .A2(new_n471), .A3(new_n226), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(KEYINPUT35), .B2(new_n517), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n939), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n940), .B2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n935), .A2(new_n945), .ZN(G367));
  NAND2_X1  g0746(.A1(new_n813), .A2(new_n237), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n807), .B1(new_n219), .B2(new_n303), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n821), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n616), .A2(new_n686), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n653), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n625), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n787), .A2(new_n202), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n782), .B2(new_n843), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n769), .A2(new_n242), .B1(new_n764), .B2(new_n846), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n361), .B(new_n956), .C1(G150), .C2(new_n771), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n799), .A2(G77), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n285), .B2(new_n774), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G159), .B2(new_n760), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n955), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n756), .A2(new_n557), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n811), .B(new_n962), .C1(G294), .C2(new_n760), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n309), .B2(new_n787), .C1(new_n792), .C2(new_n781), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n771), .A2(G303), .B1(new_n765), .B2(G317), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n796), .A2(KEYINPUT46), .A3(G116), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT46), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n774), .B2(new_n471), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n844), .A2(G283), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n965), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n961), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT47), .Z(new_n972));
  OAI221_X1 g0772(.A(new_n949), .B1(new_n953), .B2(new_n823), .C1(new_n972), .C2(new_n754), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n552), .B1(new_n528), .B2(new_n692), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT111), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n550), .A2(new_n693), .A3(new_n664), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n695), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT45), .B1(new_n695), .B2(new_n978), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n976), .A2(new_n977), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n981), .A2(KEYINPUT44), .A3(new_n694), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT44), .B1(new_n981), .B2(new_n694), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n979), .A2(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(new_n683), .A3(new_n687), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n688), .B1(new_n982), .B2(new_n983), .C1(new_n979), .C2(new_n980), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n691), .B1(new_n687), .B2(new_n690), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n683), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n751), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n751), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n697), .B(KEYINPUT41), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n819), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n742), .B1(new_n981), .B2(new_n506), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n692), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT42), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n981), .B2(new_n691), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n978), .A2(KEYINPUT42), .A3(new_n689), .A4(new_n690), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n1000), .A2(KEYINPUT43), .A3(new_n953), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n953), .B(KEYINPUT43), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT112), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1000), .A2(KEYINPUT112), .A3(new_n1002), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n688), .A2(new_n981), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1001), .A2(new_n1005), .A3(new_n1008), .A4(new_n1006), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n973), .B1(new_n993), .B2(new_n1012), .ZN(G387));
  OR2_X1    g0813(.A1(new_n687), .A2(new_n823), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G317), .A2(new_n771), .B1(new_n844), .B2(G303), .ZN(new_n1015));
  INV_X1    g0815(.A(G322), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n792), .B2(new_n761), .C1(new_n781), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n788), .A2(G283), .B1(G294), .B2(new_n796), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT49), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n756), .A2(new_n471), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n811), .B(new_n1026), .C1(G326), .C2(new_n765), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G68), .A2(new_n844), .B1(new_n765), .B2(G150), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n242), .B2(new_n772), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n289), .B2(new_n760), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n774), .A2(new_n267), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n849), .A2(new_n962), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n788), .A2(new_n303), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n782), .A2(G159), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n754), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n809), .A2(new_n698), .B1(new_n309), .B2(new_n219), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT113), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n445), .B1(new_n202), .B2(new_n267), .C1(new_n698), .C2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1039), .B2(new_n698), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n300), .A2(G50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n813), .B(new_n1044), .C1(new_n234), .C2(new_n445), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1047), .A2(new_n1048), .A3(new_n807), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1037), .A2(new_n821), .A3(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n989), .A2(new_n819), .B1(new_n1014), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n990), .A2(new_n697), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n751), .A2(new_n989), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(G393));
  NAND2_X1  g0854(.A1(new_n813), .A2(new_n241), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n807), .B1(new_n219), .B2(G97), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n821), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(G159), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n781), .A2(new_n281), .B1(new_n1058), .B2(new_n772), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT115), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT51), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n788), .A2(G77), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n854), .B1(new_n202), .B2(new_n774), .C1(new_n761), .C2(new_n242), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n769), .A2(new_n300), .B1(new_n764), .B2(new_n842), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1063), .A2(new_n849), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1060), .A2(KEYINPUT51), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n782), .A2(G317), .B1(G311), .B2(new_n771), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  OAI221_X1 g0870(.A(new_n361), .B1(new_n764), .B2(new_n1016), .C1(new_n858), .C2(new_n769), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n757), .B1(G283), .B2(new_n796), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n571), .B2(new_n761), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G116), .C2(new_n788), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1068), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1057), .B1(new_n754), .B2(new_n1075), .C1(new_n978), .C2(new_n823), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n987), .B2(new_n818), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n697), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n987), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n990), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n987), .A2(new_n990), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1077), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G390));
  OAI21_X1  g0884(.A(new_n891), .B1(new_n902), .B2(KEYINPUT39), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n914), .A2(new_n892), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n913), .A2(new_n750), .A3(G330), .A4(new_n863), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n895), .A2(new_n900), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT38), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n888), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n893), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n710), .A2(new_n686), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT98), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n710), .A2(KEYINPUT98), .A3(new_n686), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n834), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n832), .A3(new_n913), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1093), .A2(new_n1099), .A3(KEYINPUT116), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT116), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1087), .B(new_n1088), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT116), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1098), .A2(new_n832), .A3(new_n913), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n892), .B1(new_n901), .B2(new_n888), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1093), .A2(new_n1099), .A3(KEYINPUT116), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1106), .A2(new_n1107), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n913), .A2(new_n923), .A3(G330), .A4(new_n863), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1102), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n736), .A2(new_n737), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n498), .A2(new_n506), .A3(new_n692), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n748), .B(new_n749), .C1(new_n627), .C2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n863), .B(G330), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n908), .A2(new_n910), .A3(new_n912), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1109), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n904), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n923), .A2(G330), .A3(new_n863), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1115), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n711), .A2(new_n712), .A3(new_n833), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n832), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1088), .B(new_n1120), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n931), .A2(G330), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n872), .A2(new_n1124), .A3(new_n646), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1110), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1087), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1109), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AND4_X1   g0930(.A1(new_n646), .A2(new_n872), .A3(new_n1125), .A4(new_n1124), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n1102), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(new_n697), .A3(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n819), .B(new_n1102), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1085), .A2(new_n803), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n840), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n820), .B1(new_n289), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT117), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n772), .A2(new_n471), .B1(new_n764), .B2(new_n858), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n264), .B(new_n1139), .C1(G97), .C2(new_n844), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n782), .A2(G283), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n756), .A2(new_n202), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n775), .B(new_n1142), .C1(G107), .C2(new_n760), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1062), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n264), .B1(new_n756), .B2(new_n242), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT118), .ZN(new_n1146));
  INV_X1    g0946(.A(G128), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n781), .C1(new_n1058), .C2(new_n787), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n771), .A2(G132), .ZN(new_n1149));
  INV_X1    g0949(.A(G125), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1149), .B1(new_n764), .B2(new_n1150), .C1(new_n769), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n774), .A2(new_n281), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(new_n846), .C2(new_n761), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1144), .B1(new_n1148), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1138), .B1(new_n1157), .B2(new_n753), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1135), .A2(new_n1158), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1134), .A2(KEYINPUT119), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT119), .B1(new_n1134), .B2(new_n1159), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1133), .B1(new_n1160), .B2(new_n1161), .ZN(G378));
  NAND3_X1  g0962(.A1(new_n872), .A2(new_n646), .A3(new_n1125), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1132), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n744), .A2(new_n922), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n835), .B1(new_n1166), .B2(new_n738), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(new_n913), .C1(new_n888), .C2(new_n889), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n921), .B1(new_n1168), .B2(new_n926), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n321), .A2(new_n677), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n645), .A2(new_n298), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n298), .B1(new_n333), .B2(new_n334), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1170), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1169), .A2(new_n925), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1169), .B2(new_n925), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n919), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n925), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n928), .A2(G330), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1182), .A2(new_n1183), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n903), .A2(new_n918), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1169), .A2(new_n925), .A3(new_n1178), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1181), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1184), .A2(new_n1185), .A3(KEYINPUT121), .A4(new_n1186), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(KEYINPUT57), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n697), .B1(new_n1165), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1132), .A2(new_n1164), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1181), .A2(new_n1187), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT57), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1176), .A2(new_n1177), .A3(new_n804), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n756), .A2(new_n285), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1032), .B(new_n1198), .C1(G97), .C2(new_n760), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n811), .A2(G41), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n765), .A2(G283), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G107), .A2(new_n771), .B1(new_n844), .B2(new_n303), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n954), .B(new_n1203), .C1(G116), .C2(new_n782), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT58), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n242), .B1(G33), .B2(G41), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1200), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT120), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n774), .A2(new_n1151), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n772), .A2(new_n1147), .B1(new_n769), .B2(new_n846), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(G132), .C2(new_n760), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n1150), .B2(new_n781), .C1(new_n281), .C2(new_n787), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n799), .A2(G159), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n765), .C2(G124), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1209), .B1(KEYINPUT58), .B2(new_n1204), .C1(new_n1214), .C2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n753), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n820), .C1(G50), .C2(new_n1136), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1197), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1194), .B2(new_n819), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1196), .A2(new_n1223), .ZN(G375));
  INV_X1    g1024(.A(new_n1124), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1163), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n992), .A3(new_n1126), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1115), .A2(new_n803), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n820), .B1(G68), .B2(new_n1136), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1034), .B1(new_n858), .B2(new_n781), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G107), .A2(new_n844), .B1(new_n765), .B2(G303), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1231), .B(new_n361), .C1(new_n855), .C2(new_n772), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n958), .B1(new_n557), .B2(new_n774), .C1(new_n761), .C2(new_n471), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1235), .A2(KEYINPUT122), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n761), .A2(new_n1151), .B1(new_n1058), .B2(new_n774), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n771), .A2(G137), .B1(new_n765), .B2(G128), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n281), .B2(new_n769), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(G132), .C2(new_n782), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n849), .A2(new_n1198), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT123), .Z(new_n1242));
  OAI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(new_n242), .C2(new_n787), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1235), .A2(KEYINPUT122), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1236), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1229), .B1(new_n1245), .B2(new_n753), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1124), .A2(new_n819), .B1(new_n1228), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1227), .A2(new_n1247), .ZN(G381));
  NOR2_X1   g1048(.A1(G375), .A2(G378), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1083), .B(new_n973), .C1(new_n993), .C2(new_n1012), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  OR3_X1    g1052(.A1(G381), .A2(G384), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT124), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1251), .A2(KEYINPUT124), .A3(new_n1254), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1249), .B1(new_n1255), .B2(new_n1256), .ZN(G407));
  NAND2_X1  g1057(.A1(new_n678), .A2(G213), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1249), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G407), .A2(G213), .A3(new_n1260), .ZN(G409));
  OAI211_X1 g1061(.A(G378), .B(new_n1223), .C1(new_n1192), .C2(new_n1195), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1161), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1134), .A2(KEYINPUT119), .A3(new_n1159), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1193), .A2(new_n992), .A3(new_n1194), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1189), .A2(new_n819), .A3(new_n1190), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1197), .B2(new_n1221), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1265), .B(new_n1133), .C1(new_n1266), .C2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1258), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1226), .B1(new_n1131), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n1225), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n697), .A3(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(G384), .A3(new_n1247), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1275), .B2(new_n1247), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G2897), .B(new_n1259), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1278), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1259), .A2(G2897), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1276), .A3(new_n1281), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1271), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G387), .A2(G390), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1250), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1252), .A2(KEYINPUT125), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT125), .B1(new_n1252), .B2(new_n1291), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(KEYINPUT126), .B1(new_n1290), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1295), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1250), .A4(new_n1289), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1252), .A2(new_n1291), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1290), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1296), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1259), .B1(new_n1262), .B2(new_n1269), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1286), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1284), .A2(new_n1288), .A3(new_n1302), .A4(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT62), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1303), .A2(new_n1306), .A3(new_n1286), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1303), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1306), .B1(new_n1303), .B2(new_n1286), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1307), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1305), .B1(new_n1312), .B2(new_n1302), .ZN(G405));
  INV_X1    g1113(.A(G378), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G375), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(new_n1287), .A3(new_n1262), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1302), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G378), .B1(new_n1196), .B2(new_n1223), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1262), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1286), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1316), .A2(new_n1317), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1317), .B1(new_n1320), .B2(new_n1316), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(G402));
endmodule


