//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(new_n202), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G87), .B2(G250), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT65), .B(G77), .Z(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n221), .B(new_n222), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n213), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n216), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n209), .ZN(new_n248));
  INV_X1    g0048(.A(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT67), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G58), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT8), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT8), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT8), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n257), .A3(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n210), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT69), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n259), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n267));
  INV_X1    g0067(.A(G150), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n248), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G50), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT70), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n277), .A2(new_n274), .A3(G13), .A4(G20), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n248), .B1(new_n276), .B2(new_n278), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n210), .A2(G1), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n273), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n273), .A2(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n272), .A2(KEYINPUT9), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT73), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n272), .A2(new_n283), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT9), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n293), .A3(G274), .ZN(new_n294));
  INV_X1    g0094(.A(G226), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT3), .B(G33), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(G223), .A3(G1698), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT66), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT66), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G1698), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n301), .A2(new_n303), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G222), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n300), .B1(new_n308), .B2(new_n309), .C1(new_n224), .C2(new_n299), .ZN(new_n310));
  INV_X1    g0110(.A(new_n293), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n298), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(G190), .B2(new_n312), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n285), .A2(new_n288), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT10), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n285), .A2(new_n318), .A3(new_n288), .A4(new_n315), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n293), .A2(G238), .A3(new_n296), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n294), .A2(new_n321), .A3(KEYINPUT74), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT74), .B1(new_n294), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G232), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(new_n304), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n299), .A2(new_n326), .B1(G33), .B2(G97), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT66), .B(G1698), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n299), .A2(new_n328), .A3(G226), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n293), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT13), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n329), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n311), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(new_n323), .C2(new_n322), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n331), .B2(new_n335), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n338), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n339), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT12), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n279), .A2(new_n346), .A3(new_n218), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n276), .A2(new_n278), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT12), .B1(new_n348), .B2(G68), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n280), .B(G68), .C1(G1), .C2(new_n210), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n265), .A2(G77), .A3(new_n261), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT11), .B1(new_n355), .B2(new_n248), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT75), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT11), .ZN(new_n361));
  INV_X1    g0161(.A(new_n248), .ZN(new_n362));
  AOI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(new_n353), .C2(new_n354), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT75), .B1(new_n356), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n352), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n345), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n286), .B1(G169), .B2(new_n312), .ZN(new_n368));
  AND2_X1   g0168(.A1(KEYINPUT71), .A2(G179), .ZN(new_n369));
  NOR2_X1   g0169(.A1(KEYINPUT71), .A2(G179), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n312), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n308), .A2(new_n325), .B1(new_n376), .B2(new_n299), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n301), .A2(new_n303), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n378), .A2(new_n219), .A3(new_n304), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n311), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n294), .ZN(new_n381));
  INV_X1    g0181(.A(new_n297), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(G244), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n340), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT15), .B(G87), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT72), .B1(new_n386), .B2(new_n260), .ZN(new_n387));
  XOR2_X1   g0187(.A(KEYINPUT8), .B(G58), .Z(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n387), .B1(new_n224), .B2(new_n210), .C1(new_n270), .C2(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n386), .A2(KEYINPUT72), .A3(new_n260), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n248), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G77), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n281), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n224), .A2(new_n279), .B1(new_n280), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n385), .B(new_n396), .C1(new_n371), .C2(new_n384), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n384), .A2(G200), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n380), .A2(G190), .A3(new_n383), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(new_n392), .A4(new_n395), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n320), .A2(new_n367), .A3(new_n375), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G190), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n331), .A2(new_n335), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(G200), .B1(new_n331), .B2(new_n335), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n365), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT76), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n365), .B(KEYINPUT76), .C1(new_n404), .C2(new_n405), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(KEYINPUT77), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT77), .B1(new_n408), .B2(new_n409), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n250), .A2(new_n252), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n201), .B1(new_n415), .B2(G68), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT78), .B1(new_n416), .B2(new_n210), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n269), .A2(G159), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT78), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n218), .B1(new_n250), .B2(new_n252), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(G20), .C1(new_n420), .C2(new_n201), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT7), .B1(new_n378), .B2(new_n210), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT7), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n424), .B(G20), .C1(new_n301), .C2(new_n303), .ZN(new_n425));
  OAI21_X1  g0225(.A(G68), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n414), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(KEYINPUT16), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(new_n248), .C1(new_n422), .C2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT67), .B(G58), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n249), .B1(KEYINPUT68), .B2(new_n256), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n431), .A2(KEYINPUT8), .B1(new_n432), .B2(new_n255), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n279), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n281), .B1(new_n253), .B2(new_n258), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n280), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n433), .A2(KEYINPUT79), .A3(new_n281), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT80), .B(new_n434), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT79), .B1(new_n433), .B2(new_n281), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(new_n436), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n280), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT80), .B1(new_n443), .B2(new_n434), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n299), .A2(new_n328), .A3(G223), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G226), .A2(G1698), .ZN(new_n447));
  INV_X1    g0247(.A(G87), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n378), .A2(new_n447), .B1(new_n262), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n311), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n451));
  INV_X1    g0251(.A(new_n447), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n299), .A2(new_n452), .B1(G33), .B2(G87), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n299), .A2(new_n328), .A3(G223), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n293), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n294), .B(new_n403), .C1(new_n325), .C2(new_n297), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n451), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n294), .B1(new_n325), .B2(new_n297), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n450), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n313), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n460), .A2(KEYINPUT82), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT82), .B1(new_n460), .B2(new_n464), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n430), .B(new_n445), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n421), .A2(new_n418), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n202), .B1(new_n431), .B2(new_n218), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n419), .B1(new_n472), .B2(G20), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT16), .B1(new_n474), .B2(new_n426), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n248), .B1(new_n422), .B2(new_n429), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n439), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n453), .A2(new_n454), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n456), .B1(new_n484), .B2(new_n311), .ZN(new_n485));
  AOI211_X1 g0285(.A(KEYINPUT81), .B(new_n293), .C1(new_n453), .C2(new_n454), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n485), .A2(new_n486), .A3(new_n458), .ZN(new_n487));
  AOI21_X1  g0287(.A(G200), .B1(new_n450), .B2(new_n462), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n460), .A2(KEYINPUT82), .A3(new_n464), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT17), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(KEYINPUT83), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n482), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n470), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n480), .B(new_n439), .C1(new_n475), .C2(new_n476), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT18), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n485), .A2(new_n486), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n461), .A2(new_n371), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n499), .A2(new_n500), .B1(new_n340), .B2(new_n463), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n498), .B1(new_n497), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n402), .A2(new_n413), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n301), .A2(new_n303), .A3(G257), .A4(G1698), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G294), .ZN(new_n509));
  INV_X1    g0309(.A(G250), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n508), .B(new_n509), .C1(new_n308), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n274), .A2(G45), .ZN(new_n512));
  OR2_X1    g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  NAND2_X1  g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n311), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n511), .A2(new_n311), .B1(G264), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n514), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n290), .A2(G1), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(G274), .A3(new_n293), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT89), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT89), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n517), .A2(new_n523), .A3(new_n520), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(G169), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n521), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G179), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n348), .B2(G107), .ZN(new_n530));
  INV_X1    g0330(.A(new_n529), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n276), .A2(new_n376), .A3(new_n278), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n274), .A2(G33), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT84), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n280), .A2(new_n537), .A3(G107), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT88), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT88), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n534), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n210), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n545), .A2(new_n546), .B1(new_n263), .B2(G116), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n301), .A2(new_n303), .A3(new_n210), .A4(G87), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n548), .A2(KEYINPUT22), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(KEYINPUT22), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT24), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n362), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n543), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n528), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n540), .A2(new_n542), .B1(new_n553), .B2(new_n554), .ZN(new_n558));
  AOI21_X1  g0358(.A(G190), .B1(new_n522), .B2(new_n524), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n526), .A2(G200), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n299), .A2(new_n328), .A3(KEYINPUT4), .A4(G244), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G283), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n299), .A2(G250), .A3(G1698), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT4), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n308), .B2(new_n225), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n293), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(KEYINPUT5), .A2(G41), .ZN(new_n570));
  NOR2_X1   g0370(.A1(KEYINPUT5), .A2(G41), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n519), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(G257), .A3(new_n293), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n520), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT85), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n520), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT6), .ZN(new_n580));
  INV_X1    g0380(.A(G97), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n580), .A2(new_n581), .A3(G107), .ZN(new_n582));
  XNOR2_X1  g0382(.A(G97), .B(G107), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n584), .A2(new_n210), .B1(new_n393), .B2(new_n270), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n424), .B1(new_n299), .B2(G20), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n378), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n376), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n248), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n280), .A2(new_n537), .A3(G97), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n279), .A2(new_n581), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n568), .A2(new_n564), .A3(new_n563), .A4(new_n565), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n574), .B1(new_n594), .B2(new_n311), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G190), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n579), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n301), .A2(new_n303), .A3(new_n305), .A4(new_n307), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT4), .B1(new_n599), .B2(G244), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n311), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n574), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n340), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n601), .A2(new_n372), .A3(new_n575), .A4(new_n577), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n589), .A2(new_n591), .A3(new_n590), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n597), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n299), .A2(new_n328), .A3(G257), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n299), .A2(G264), .A3(G1698), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n378), .A2(G303), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n311), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n572), .A2(G270), .A3(new_n293), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n520), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n280), .A2(new_n537), .A3(G116), .ZN(new_n618));
  INV_X1    g0418(.A(G116), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n279), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n247), .A2(new_n209), .B1(G20), .B2(new_n619), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n564), .B(new_n210), .C1(G33), .C2(new_n581), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT20), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n621), .A2(KEYINPUT20), .A3(new_n622), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n618), .B(new_n620), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n617), .A2(new_n625), .A3(G169), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n625), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n613), .A2(new_n616), .A3(G190), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n615), .B1(new_n612), .B2(new_n311), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n629), .B(new_n630), .C1(new_n313), .C2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n613), .A2(new_n616), .A3(G179), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n625), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n617), .A2(new_n625), .A3(KEYINPUT21), .A4(G169), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n628), .A2(new_n632), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n301), .A2(new_n303), .A3(G244), .A4(G1698), .ZN(new_n637));
  NAND2_X1  g0437(.A1(G33), .A2(G116), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n637), .B(new_n638), .C1(new_n308), .C2(new_n219), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n311), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n293), .A2(G274), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n512), .A2(G250), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n641), .A2(new_n512), .B1(new_n311), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n639), .B2(new_n311), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G190), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n301), .A2(new_n303), .A3(new_n210), .A4(G68), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT19), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n260), .B2(new_n581), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n210), .A2(new_n653), .B1(new_n204), .B2(new_n448), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n248), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n280), .A2(new_n537), .A3(G87), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n279), .A2(new_n386), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n646), .A2(new_n648), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n647), .A2(new_n372), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n280), .A2(new_n537), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n655), .B(new_n657), .C1(new_n386), .C2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n660), .B(new_n662), .C1(G169), .C2(new_n647), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT86), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n659), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n659), .A2(new_n663), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n608), .A2(new_n636), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n507), .A2(new_n562), .A3(new_n668), .ZN(G372));
  NOR2_X1   g0469(.A1(new_n647), .A2(new_n313), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT90), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n648), .B(new_n658), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n646), .A2(KEYINPUT90), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n663), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n608), .A2(new_n675), .A3(new_n561), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n558), .B1(new_n525), .B2(new_n527), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n628), .A2(new_n634), .A3(new_n635), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT91), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n678), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT91), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n557), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n676), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n675), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n659), .A2(new_n663), .A3(new_n664), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n664), .B1(new_n659), .B2(new_n663), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n687), .A2(new_n688), .A3(new_n607), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n686), .B(new_n663), .C1(new_n689), .C2(new_n684), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n506), .B1(new_n683), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT92), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n397), .B1(new_n408), .B2(new_n409), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n366), .B2(new_n345), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n465), .A2(new_n466), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n695), .A2(new_n497), .A3(new_n493), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n468), .B1(new_n482), .B2(new_n491), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n504), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n374), .B1(new_n699), .B2(new_n320), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n692), .A2(new_n700), .ZN(G369));
  NAND3_X1  g0501(.A1(new_n274), .A2(new_n210), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n625), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT93), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n678), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT94), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT94), .ZN(new_n712));
  INV_X1    g0512(.A(new_n636), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n709), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n556), .A2(new_n707), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT95), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n557), .A2(new_n561), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n677), .B2(new_n707), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n707), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n677), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n717), .A2(new_n718), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n678), .A2(new_n722), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n721), .A2(new_n723), .A3(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n214), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G41), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G1), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n207), .B2(new_n730), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n722), .B1(new_n683), .B2(new_n690), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT98), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n677), .A2(new_n678), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n676), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n667), .A2(new_n684), .A3(new_n665), .A4(new_n685), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT26), .B1(new_n674), .B2(new_n607), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n741), .A2(new_n663), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n557), .A2(new_n680), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n597), .A2(new_n607), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n674), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n744), .A2(new_n746), .A3(KEYINPUT98), .A4(new_n561), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n740), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(KEYINPUT29), .A3(new_n722), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n745), .A2(new_n687), .A3(new_n688), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n718), .A2(new_n636), .A3(new_n750), .A4(new_n722), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT96), .B(KEYINPUT30), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n631), .A2(G179), .A3(new_n517), .A4(new_n647), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n753), .B2(new_n603), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n601), .A2(new_n575), .A3(new_n577), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n647), .A2(new_n371), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n521), .A3(new_n617), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT97), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n517), .A2(new_n647), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n760), .A2(new_n633), .A3(KEYINPUT30), .A4(new_n595), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT97), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n754), .A2(new_n762), .A3(new_n757), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n722), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n754), .A2(new_n761), .A3(new_n757), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n707), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n764), .A2(new_n766), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n751), .A2(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n737), .A2(new_n749), .B1(G330), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n734), .B1(new_n771), .B2(G1), .ZN(G364));
  INV_X1    g0572(.A(new_n715), .ZN(new_n773));
  INV_X1    g0573(.A(G13), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n274), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n729), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G330), .B2(new_n714), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n209), .B1(G20), .B2(new_n340), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n299), .A2(new_n214), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT99), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(G116), .B2(new_n214), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n728), .A2(new_n299), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G45), .B2(new_n207), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n245), .B2(G45), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n785), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n778), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n210), .A2(new_n313), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n371), .A2(G190), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G179), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G190), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n797), .A2(G326), .B1(G294), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n210), .A2(G190), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n371), .A2(new_n313), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT100), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n371), .A2(new_n403), .A3(new_n795), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT33), .B(G317), .Z(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n313), .A2(G179), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n803), .A2(new_n798), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G283), .A2(new_n812), .B1(new_n814), .B2(G329), .ZN(new_n815));
  INV_X1    g0615(.A(G303), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n210), .A2(new_n403), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n810), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n815), .B(new_n378), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n371), .A2(new_n313), .A3(new_n817), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n809), .B(new_n819), .C1(G322), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n806), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT101), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n273), .A2(new_n796), .B1(new_n807), .B2(new_n218), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n415), .B2(new_n821), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n299), .B1(new_n811), .B2(new_n376), .C1(new_n448), .C2(new_n818), .ZN(new_n827));
  INV_X1    g0627(.A(new_n804), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(new_n223), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G159), .ZN(new_n830));
  OAI21_X1  g0630(.A(KEYINPUT32), .B1(new_n813), .B2(new_n830), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n813), .A2(KEYINPUT32), .A3(new_n830), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G97), .B2(new_n800), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n826), .A2(new_n829), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n823), .A2(KEYINPUT101), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n824), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n794), .B1(new_n836), .B2(new_n784), .ZN(new_n837));
  INV_X1    g0637(.A(new_n783), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n714), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n780), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  NOR2_X1   g0641(.A1(new_n397), .A2(new_n707), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n396), .A2(new_n707), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n400), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n842), .B1(new_n397), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n735), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n722), .B(new_n845), .C1(new_n683), .C2(new_n690), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n770), .A2(G330), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n778), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  INV_X1    g0652(.A(new_n818), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n378), .B1(new_n853), .B2(G50), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n812), .A2(G68), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n813), .ZN(new_n857));
  INV_X1    g0657(.A(new_n807), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G137), .A2(new_n797), .B1(new_n858), .B2(G150), .ZN(new_n859));
  INV_X1    g0659(.A(G143), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n860), .B2(new_n820), .C1(new_n830), .C2(new_n804), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT34), .Z(new_n862));
  AOI211_X1 g0662(.A(new_n857), .B(new_n862), .C1(new_n415), .C2(new_n800), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n378), .B1(new_n813), .B2(new_n802), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n818), .A2(new_n376), .B1(new_n811), .B2(new_n448), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(G97), .C2(new_n800), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G294), .A2(new_n821), .B1(new_n797), .B2(G303), .ZN(new_n867));
  INV_X1    g0667(.A(G283), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n619), .A2(new_n804), .B1(new_n807), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n866), .B(new_n867), .C1(KEYINPUT103), .C2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(KEYINPUT103), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n784), .B1(new_n863), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n778), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n784), .A2(new_n781), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT102), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n876), .B2(new_n393), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n872), .B(new_n877), .C1(new_n782), .C2(new_n845), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n852), .A2(new_n878), .ZN(G384));
  NOR2_X1   g0679(.A1(new_n775), .A2(new_n274), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n506), .A2(new_n737), .A3(new_n749), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n700), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT109), .ZN(new_n883));
  INV_X1    g0683(.A(new_n503), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n499), .A2(new_n500), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n463), .A2(new_n340), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n445), .B2(new_n430), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n498), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n705), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n842), .B(KEYINPUT105), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n848), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n408), .A2(new_n409), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n365), .A2(new_n722), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n367), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT77), .ZN(new_n898));
  INV_X1    g0698(.A(new_n405), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n331), .A2(new_n335), .A3(new_n403), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT76), .B1(new_n901), .B2(new_n365), .ZN(new_n902));
  INV_X1    g0702(.A(new_n409), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n345), .B1(new_n904), .B2(new_n410), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n897), .B1(new_n905), .B2(new_n896), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n893), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n497), .A2(KEYINPUT106), .A3(new_n501), .ZN(new_n909));
  INV_X1    g0709(.A(new_n705), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n497), .A2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n909), .A2(new_n467), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n497), .A2(new_n501), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT106), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n910), .B1(new_n477), .B2(new_n478), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n501), .B1(new_n477), .B2(new_n478), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n467), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n912), .A2(new_n915), .B1(KEYINPUT37), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n916), .B1(new_n496), .B2(new_n504), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n908), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n916), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n698), .B2(new_n890), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n924));
  INV_X1    g0724(.A(new_n915), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n909), .A2(new_n467), .A3(new_n911), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(KEYINPUT38), .A3(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n891), .B1(new_n907), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n921), .A2(new_n928), .A3(KEYINPUT39), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n467), .A2(new_n913), .A3(new_n911), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n912), .A2(new_n915), .B1(KEYINPUT37), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT108), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n696), .B2(new_n697), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n470), .A2(KEYINPUT108), .A3(new_n495), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n504), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n911), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n941));
  OAI21_X1  g0741(.A(new_n928), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n931), .B1(new_n932), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n345), .A2(new_n366), .A3(new_n722), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n930), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n883), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(G330), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n767), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT110), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n768), .A2(new_n765), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT110), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n767), .A2(new_n954), .A3(KEYINPUT31), .A4(new_n707), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n846), .B1(new_n956), .B2(new_n751), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n906), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n950), .B1(new_n929), .B2(new_n958), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n668), .A2(new_n562), .A3(new_n707), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n845), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n345), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n411), .B2(new_n412), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n895), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n962), .B1(new_n965), .B2(new_n897), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n942), .A2(KEYINPUT40), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n959), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n956), .A2(new_n751), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n506), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n949), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n970), .B2(new_n968), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n880), .B1(new_n948), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n948), .B2(new_n972), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n583), .A2(new_n580), .ZN(new_n975));
  INV_X1    g0775(.A(new_n582), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT35), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT35), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n978), .A2(G116), .A3(new_n211), .A4(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(KEYINPUT104), .B(KEYINPUT36), .Z(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n224), .A2(new_n207), .A3(new_n420), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n218), .A2(G50), .ZN(new_n984));
  OAI211_X1 g0784(.A(G1), .B(new_n774), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n974), .A2(new_n982), .A3(new_n985), .ZN(G367));
  NOR2_X1   g0786(.A1(new_n724), .A2(new_n725), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n608), .B1(new_n593), .B2(new_n722), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n607), .B2(new_n722), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n607), .B1(new_n988), .B2(new_n557), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n990), .A2(KEYINPUT42), .B1(new_n722), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(KEYINPUT42), .B2(new_n990), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n658), .A2(new_n722), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n674), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n663), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n994), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n720), .A2(new_n989), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n729), .B(KEYINPUT41), .Z(new_n1005));
  NAND3_X1  g0805(.A1(new_n726), .A2(new_n723), .A3(new_n989), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n726), .A2(new_n723), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT111), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT44), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n989), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1009), .B(new_n1012), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1008), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n720), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1008), .A2(new_n721), .A3(new_n1016), .A4(new_n1013), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n715), .A2(KEYINPUT112), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n715), .A2(KEYINPUT112), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n719), .A2(new_n725), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n726), .A3(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1021), .B(new_n1024), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1018), .A2(new_n1019), .A3(new_n771), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1005), .B1(new_n1026), .B2(new_n771), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1004), .B1(new_n1027), .B2(new_n777), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n790), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n785), .B1(new_n214), .B2(new_n386), .C1(new_n238), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n778), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G150), .A2(new_n821), .B1(new_n858), .B2(G159), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n273), .B2(new_n804), .C1(new_n860), .C2(new_n796), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n800), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(new_n218), .ZN(new_n1035));
  INV_X1    g0835(.A(G137), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n299), .B1(new_n813), .B2(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n224), .A2(new_n811), .B1(new_n431), .B2(new_n818), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G294), .A2(new_n858), .B1(new_n828), .B2(G283), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n802), .B2(new_n796), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n853), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT46), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n818), .B2(new_n619), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(new_n376), .C2(new_n1034), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n820), .A2(new_n816), .ZN(new_n1046));
  INV_X1    g0846(.A(G317), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n378), .B1(new_n813), .B2(new_n1047), .C1(new_n581), .C2(new_n811), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1041), .A2(new_n1045), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1039), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT47), .Z(new_n1051));
  AOI21_X1  g0851(.A(new_n1031), .B1(new_n1051), .B2(new_n784), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n995), .A2(new_n783), .A3(new_n997), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1028), .A2(new_n1054), .ZN(G387));
  OAI21_X1  g0855(.A(new_n790), .B1(new_n235), .B2(new_n290), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n731), .B2(new_n787), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n389), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1058));
  OAI21_X1  g0858(.A(KEYINPUT50), .B1(new_n389), .B2(G50), .ZN(new_n1059));
  AOI21_X1  g0859(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1058), .A2(new_n731), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1057), .A2(new_n1061), .B1(new_n376), .B2(new_n728), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n785), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n778), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n224), .A2(new_n818), .B1(new_n268), .B2(new_n813), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1034), .A2(new_n386), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n299), .B1(new_n811), .B2(new_n581), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G50), .A2(new_n821), .B1(new_n797), .B2(G159), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n858), .A2(new_n259), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n828), .A2(G68), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n299), .B1(new_n814), .B2(G326), .ZN(new_n1073));
  INV_X1    g0873(.A(G294), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1034), .A2(new_n868), .B1(new_n818), .B2(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G311), .A2(new_n858), .B1(new_n797), .B2(G322), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n816), .B2(new_n804), .C1(new_n1047), .C2(new_n820), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1073), .B1(new_n619), .B2(new_n811), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1072), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1064), .B1(new_n1084), .B2(new_n784), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n719), .A2(new_n783), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT113), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1025), .B2(new_n777), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1025), .A2(new_n771), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n729), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1025), .A2(new_n771), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(G393));
  NAND2_X1  g0893(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1090), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n729), .A3(new_n1026), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1018), .A2(new_n777), .A3(new_n1019), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n242), .A2(new_n790), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1098), .B(new_n785), .C1(new_n581), .C2(new_n214), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1074), .A2(new_n804), .B1(new_n807), .B2(new_n816), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G283), .A2(new_n853), .B1(new_n814), .B2(G322), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1101), .B(new_n378), .C1(new_n376), .C2(new_n811), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G116), .C2(new_n800), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n802), .A2(new_n820), .B1(new_n796), .B2(new_n1047), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n268), .A2(new_n796), .B1(new_n820), .B2(new_n830), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT51), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n800), .A2(G77), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G50), .A2(new_n858), .B1(new_n828), .B2(new_n388), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n378), .B1(new_n812), .B2(G87), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G68), .A2(new_n853), .B1(new_n814), .B2(G143), .ZN(new_n1111));
  AND4_X1   g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1103), .A2(new_n1105), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n784), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n778), .B(new_n1099), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT114), .Z(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n838), .B2(new_n989), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n1097), .A3(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(new_n897), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n895), .B2(new_n964), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n969), .A2(G330), .A3(new_n845), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n945), .B1(new_n893), .B2(new_n906), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n937), .A2(new_n504), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT108), .B1(new_n470), .B2(new_n495), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n939), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n934), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n941), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n928), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n932), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n921), .A2(new_n928), .A3(KEYINPUT39), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1123), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n944), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n748), .A2(new_n722), .A3(new_n845), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1134), .A2(new_n892), .B1(new_n965), .B2(new_n897), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1122), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1134), .A2(new_n892), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n944), .B(new_n942), .C1(new_n1138), .C2(new_n1120), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n949), .B(new_n846), .C1(new_n751), .C2(new_n769), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n906), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n943), .C2(new_n1123), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1142), .A3(new_n777), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n778), .B1(new_n875), .B2(new_n259), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G107), .A2(new_n858), .B1(new_n821), .B2(G116), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n581), .B2(new_n804), .C1(new_n868), .C2(new_n796), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n299), .B1(new_n853), .B2(G87), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n814), .A2(G294), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1147), .A2(new_n855), .A3(new_n1108), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n853), .A2(G150), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1150), .A2(KEYINPUT53), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1150), .A2(KEYINPUT53), .B1(G159), .B2(new_n800), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n797), .A2(G128), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n299), .B1(new_n811), .B2(new_n273), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G125), .B2(new_n814), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT54), .B(G143), .Z(new_n1157));
  AOI22_X1  g0957(.A1(G132), .A2(new_n821), .B1(new_n828), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1036), .B2(new_n807), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1146), .A2(new_n1149), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1144), .B1(new_n1160), .B2(new_n784), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n943), .B2(new_n782), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1143), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n506), .A2(G330), .A3(new_n969), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n881), .A2(new_n1164), .A3(new_n700), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1140), .A2(new_n906), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n893), .B1(new_n1122), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1138), .A2(new_n1168), .A3(new_n1141), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1165), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1137), .A2(new_n1142), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1171), .A2(KEYINPUT115), .A3(new_n729), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1165), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT115), .B1(new_n1171), .B2(new_n729), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1163), .B1(new_n1178), .B2(new_n1179), .ZN(G378));
  INV_X1    g0980(.A(KEYINPUT117), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n959), .A2(new_n967), .A3(G330), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n320), .A2(new_n375), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n705), .B1(new_n272), .B2(new_n283), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OR3_X1    g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1182), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n959), .A3(new_n967), .A4(G330), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT116), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n946), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n946), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(new_n1196), .A3(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1198), .A2(new_n1200), .B1(new_n1175), .B2(new_n1171), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1181), .B1(new_n1201), .B2(KEYINPUT57), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1203));
  AOI211_X1 g1003(.A(KEYINPUT116), .B(new_n946), .C1(new_n1194), .C2(new_n1193), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1199), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(KEYINPUT117), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1203), .A2(KEYINPUT57), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1193), .A2(new_n946), .A3(new_n1194), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n946), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n729), .B1(new_n1209), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1202), .A2(new_n1208), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1191), .A2(new_n782), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G125), .A2(new_n797), .B1(new_n821), .B2(G128), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1036), .B2(new_n804), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n853), .A2(new_n1157), .B1(new_n800), .B2(G150), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n856), .B2(new_n807), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n262), .B(new_n289), .C1(new_n811), .C2(new_n830), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G124), .B2(new_n814), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G97), .A2(new_n858), .B1(new_n821), .B2(G107), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n619), .B2(new_n796), .C1(new_n386), .C2(new_n804), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n224), .A2(new_n818), .B1(new_n868), .B2(new_n813), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n289), .B(new_n378), .C1(new_n811), .C2(new_n431), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1230), .A2(new_n1035), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT58), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT58), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G50), .B1(new_n262), .B2(new_n289), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n299), .B2(G41), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n1228), .A2(new_n1234), .A3(new_n1235), .A4(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n778), .B1(G50), .B2(new_n875), .C1(new_n1238), .C2(new_n1114), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1217), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n777), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1216), .A2(new_n1242), .ZN(G375));
  NAND2_X1  g1043(.A1(new_n1174), .A2(new_n777), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n873), .B1(new_n876), .B2(new_n218), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n299), .B1(new_n814), .B2(G303), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n393), .B2(new_n811), .C1(new_n581), .C2(new_n818), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n868), .A2(new_n820), .B1(new_n796), .B2(new_n1074), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n376), .A2(new_n804), .B1(new_n807), .B2(new_n619), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1066), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G159), .A2(new_n853), .B1(new_n814), .B2(G128), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n273), .B2(new_n1034), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n299), .B1(new_n811), .B2(new_n431), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT118), .Z(new_n1254));
  AOI211_X1 g1054(.A(new_n1252), .B(new_n1254), .C1(G137), .C2(new_n821), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n856), .A2(new_n796), .B1(new_n804), .B2(new_n268), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n858), .B2(new_n1157), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1250), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1245), .B1(new_n1114), .B2(new_n1258), .C1(new_n906), .C2(new_n782), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1244), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1170), .A2(new_n1005), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1167), .A2(new_n1169), .A3(new_n1165), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1262), .B2(new_n1264), .ZN(G381));
  INV_X1    g1065(.A(new_n1054), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1026), .A2(new_n771), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n776), .B1(new_n1267), .B2(new_n1005), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1266), .B1(new_n1268), .B2(new_n1004), .ZN(new_n1269));
  INV_X1    g1069(.A(G390), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1242), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1214), .B1(new_n1274), .B2(new_n1181), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1275), .B2(new_n1208), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT119), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G378), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(KEYINPUT119), .B(new_n1163), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n840), .B(new_n1089), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(G381), .A2(G384), .A3(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1272), .A2(new_n1276), .A3(new_n1280), .A4(new_n1282), .ZN(G407));
  NAND2_X1  g1083(.A1(new_n706), .A2(G213), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1276), .A2(new_n1280), .A3(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(G407), .A2(G213), .A3(new_n1286), .ZN(new_n1287));
  XOR2_X1   g1087(.A(new_n1287), .B(KEYINPUT120), .Z(G409));
  OAI21_X1  g1088(.A(G390), .B1(new_n1269), .B2(KEYINPUT126), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G387), .A2(new_n1290), .A3(new_n1270), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G393), .A2(G396), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT124), .B1(new_n1292), .B2(new_n1281), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(KEYINPUT124), .A3(new_n1281), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1289), .A2(new_n1291), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(G390), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT125), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1294), .A2(new_n1299), .A3(new_n1295), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1295), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT125), .B1(new_n1301), .B2(new_n1293), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1271), .A2(new_n1298), .A3(new_n1300), .A4(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(G384), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1167), .A2(new_n1165), .A3(new_n1169), .A4(KEYINPUT60), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n729), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1176), .A2(KEYINPUT60), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n1263), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1306), .B1(new_n1310), .B2(new_n1260), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1264), .B1(KEYINPUT60), .B2(new_n1176), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G384), .B(new_n1261), .C1(new_n1312), .C2(new_n1308), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1285), .A2(KEYINPUT122), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1311), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT123), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1285), .A2(G2897), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT123), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1311), .A2(new_n1313), .A3(new_n1318), .A4(new_n1314), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1316), .B2(new_n1319), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1210), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1240), .B1(new_n1324), .B2(new_n777), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n1206), .B2(new_n1005), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1278), .A2(new_n1279), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(new_n1276), .B2(G378), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1322), .B1(new_n1328), .B2(new_n1285), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1216), .A2(G378), .A3(new_n1242), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1278), .A2(new_n1279), .A3(new_n1326), .ZN(new_n1333));
  AOI211_X1 g1133(.A(new_n1285), .B(new_n1331), .C1(new_n1332), .C2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT121), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1335), .B1(new_n1336), .B2(KEYINPUT62), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1329), .B(new_n1330), .C1(new_n1334), .C2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1331), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1339), .A2(KEYINPUT121), .A3(new_n1284), .A4(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT62), .B1(new_n1341), .B2(new_n1336), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1305), .B1(new_n1338), .B2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1285), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1344));
  OR2_X1    g1144(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1304), .B(new_n1330), .C1(new_n1344), .C2(new_n1345), .ZN(new_n1346));
  AND4_X1   g1146(.A1(KEYINPUT63), .A2(new_n1339), .A3(new_n1284), .A4(new_n1340), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1339), .A2(new_n1284), .A3(new_n1340), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1335), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT63), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1350), .A2(new_n1351), .A3(new_n1341), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1348), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1343), .A2(new_n1353), .ZN(G405));
  NAND2_X1  g1154(.A1(G375), .A2(new_n1280), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1332), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1340), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1355), .A2(new_n1332), .A3(new_n1331), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1359), .B(new_n1305), .ZN(G402));
endmodule


