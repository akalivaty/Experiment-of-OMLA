

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587;

  XNOR2_X2 U320 ( .A(n307), .B(G218GAT), .ZN(n362) );
  XNOR2_X2 U321 ( .A(G36GAT), .B(G190GAT), .ZN(n307) );
  XNOR2_X2 U322 ( .A(n354), .B(n353), .ZN(n533) );
  NOR2_X2 U323 ( .A1(n485), .A2(n477), .ZN(n567) );
  NOR2_X1 U324 ( .A1(n531), .A2(n500), .ZN(n450) );
  XOR2_X1 U325 ( .A(n314), .B(n421), .Z(n288) );
  XOR2_X1 U326 ( .A(n384), .B(n383), .Z(n289) );
  XNOR2_X1 U327 ( .A(KEYINPUT25), .B(KEYINPUT95), .ZN(n400) );
  XNOR2_X1 U328 ( .A(n401), .B(n400), .ZN(n405) );
  XNOR2_X1 U329 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U330 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U331 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n468) );
  XNOR2_X1 U332 ( .A(n469), .B(n468), .ZN(n483) );
  XOR2_X1 U333 ( .A(KEYINPUT36), .B(n557), .Z(n585) );
  INV_X1 U334 ( .A(G190GAT), .ZN(n478) );
  XOR2_X1 U335 ( .A(n325), .B(n324), .Z(n557) );
  XOR2_X1 U336 ( .A(KEYINPUT101), .B(n451), .Z(n515) );
  XNOR2_X1 U337 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U338 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U339 ( .A(n481), .B(n480), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n291) );
  XNOR2_X1 U342 ( .A(G127GAT), .B(G211GAT), .ZN(n290) );
  XNOR2_X1 U343 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U344 ( .A(G8GAT), .B(G183GAT), .Z(n355) );
  XOR2_X1 U345 ( .A(n292), .B(n355), .Z(n297) );
  XOR2_X1 U346 ( .A(G15GAT), .B(G1GAT), .Z(n435) );
  XOR2_X1 U347 ( .A(KEYINPUT68), .B(KEYINPUT13), .Z(n294) );
  XNOR2_X1 U348 ( .A(G71GAT), .B(G78GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U350 ( .A(G57GAT), .B(n295), .Z(n429) );
  XNOR2_X1 U351 ( .A(n435), .B(n429), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U353 ( .A(G64GAT), .B(KEYINPUT76), .Z(n299) );
  NAND2_X1 U354 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U356 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U357 ( .A(G22GAT), .B(G155GAT), .Z(n389) );
  XOR2_X1 U358 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n303) );
  XNOR2_X1 U359 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n389), .B(n304), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n555) );
  NAND2_X1 U363 ( .A1(n362), .A2(G92GAT), .ZN(n311) );
  INV_X1 U364 ( .A(n362), .ZN(n309) );
  INV_X1 U365 ( .A(G92GAT), .ZN(n308) );
  NAND2_X1 U366 ( .A1(n309), .A2(n308), .ZN(n310) );
  NAND2_X1 U367 ( .A1(n311), .A2(n310), .ZN(n313) );
  AND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U370 ( .A(G99GAT), .B(G85GAT), .Z(n421) );
  XOR2_X1 U371 ( .A(G29GAT), .B(G43GAT), .Z(n316) );
  XNOR2_X1 U372 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n434) );
  XOR2_X1 U374 ( .A(G50GAT), .B(G162GAT), .Z(n383) );
  XNOR2_X1 U375 ( .A(n434), .B(n383), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n288), .B(n317), .ZN(n325) );
  XOR2_X1 U377 ( .A(KEYINPUT9), .B(KEYINPUT72), .Z(n319) );
  XNOR2_X1 U378 ( .A(KEYINPUT74), .B(KEYINPUT10), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U380 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n321) );
  XNOR2_X1 U381 ( .A(G134GAT), .B(G106GAT), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U383 ( .A(n323), .B(n322), .Z(n324) );
  XOR2_X1 U384 ( .A(KEYINPUT91), .B(G148GAT), .Z(n327) );
  XNOR2_X1 U385 ( .A(G29GAT), .B(G155GAT), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U387 ( .A(G162GAT), .B(G85GAT), .Z(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n352) );
  XOR2_X1 U389 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n331) );
  XNOR2_X1 U390 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U392 ( .A(n332), .B(G127GAT), .Z(n334) );
  XNOR2_X1 U393 ( .A(G113GAT), .B(G120GAT), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n378) );
  XOR2_X1 U395 ( .A(G57GAT), .B(KEYINPUT88), .Z(n336) );
  XNOR2_X1 U396 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n378), .B(n337), .ZN(n341) );
  XOR2_X1 U399 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n339) );
  XNOR2_X1 U400 ( .A(KEYINPUT5), .B(KEYINPUT87), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U403 ( .A(n342), .B(KEYINPUT4), .Z(n350) );
  INV_X1 U404 ( .A(KEYINPUT3), .ZN(n343) );
  NAND2_X1 U405 ( .A1(KEYINPUT84), .A2(n343), .ZN(n346) );
  INV_X1 U406 ( .A(KEYINPUT84), .ZN(n344) );
  NAND2_X1 U407 ( .A1(n344), .A2(KEYINPUT3), .ZN(n345) );
  NAND2_X1 U408 ( .A1(n346), .A2(n345), .ZN(n348) );
  XNOR2_X1 U409 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n384) );
  XNOR2_X1 U411 ( .A(G1GAT), .B(n384), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n354) );
  NAND2_X1 U414 ( .A1(G225GAT), .A2(G233GAT), .ZN(n353) );
  XOR2_X1 U415 ( .A(KEYINPUT92), .B(n355), .Z(n357) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n360) );
  XOR2_X1 U418 ( .A(G64GAT), .B(G92GAT), .Z(n359) );
  XNOR2_X1 U419 ( .A(G176GAT), .B(G204GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n420) );
  XOR2_X1 U421 ( .A(n360), .B(n420), .Z(n364) );
  XNOR2_X1 U422 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n361), .B(G211GAT), .ZN(n394) );
  XNOR2_X1 U424 ( .A(n394), .B(n362), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U426 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n366) );
  XNOR2_X1 U427 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(n367), .ZN(n379) );
  XNOR2_X1 U430 ( .A(n368), .B(n379), .ZN(n535) );
  XOR2_X1 U431 ( .A(KEYINPUT20), .B(G71GAT), .Z(n370) );
  XNOR2_X1 U432 ( .A(G43GAT), .B(G15GAT), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U434 ( .A(G190GAT), .B(G99GAT), .Z(n372) );
  XNOR2_X1 U435 ( .A(G183GAT), .B(G176GAT), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U437 ( .A(n374), .B(n373), .Z(n376) );
  NAND2_X1 U438 ( .A1(G227GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n485) );
  INV_X1 U442 ( .A(n485), .ZN(n537) );
  NAND2_X1 U443 ( .A1(n535), .A2(n537), .ZN(n399) );
  XOR2_X1 U444 ( .A(KEYINPUT82), .B(G204GAT), .Z(n382) );
  XNOR2_X1 U445 ( .A(KEYINPUT85), .B(G78GAT), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n398) );
  NAND2_X1 U447 ( .A1(G228GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n289), .B(n385), .ZN(n392) );
  XOR2_X1 U449 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n387) );
  XNOR2_X1 U450 ( .A(G218GAT), .B(KEYINPUT86), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U452 ( .A(G106GAT), .B(G148GAT), .Z(n422) );
  XOR2_X1 U453 ( .A(n388), .B(n422), .Z(n390) );
  XOR2_X1 U454 ( .A(KEYINPUT83), .B(n393), .Z(n396) );
  XNOR2_X1 U455 ( .A(n394), .B(KEYINPUT24), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n474) );
  NAND2_X1 U458 ( .A1(n399), .A2(n474), .ZN(n401) );
  NOR2_X1 U459 ( .A1(n537), .A2(n474), .ZN(n403) );
  XNOR2_X1 U460 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n571) );
  XNOR2_X1 U462 ( .A(n535), .B(KEYINPUT27), .ZN(n408) );
  NAND2_X1 U463 ( .A1(n571), .A2(n408), .ZN(n404) );
  NAND2_X1 U464 ( .A1(n405), .A2(n404), .ZN(n406) );
  XOR2_X1 U465 ( .A(n406), .B(KEYINPUT96), .Z(n407) );
  NOR2_X1 U466 ( .A1(n533), .A2(n407), .ZN(n413) );
  NAND2_X1 U467 ( .A1(n533), .A2(n408), .ZN(n482) );
  XNOR2_X1 U468 ( .A(KEYINPUT28), .B(KEYINPUT64), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n409), .B(n474), .ZN(n507) );
  NAND2_X1 U470 ( .A1(n485), .A2(n507), .ZN(n410) );
  NOR2_X1 U471 ( .A1(n482), .A2(n410), .ZN(n411) );
  XOR2_X1 U472 ( .A(KEYINPUT93), .B(n411), .Z(n412) );
  NOR2_X1 U473 ( .A1(n413), .A2(n412), .ZN(n497) );
  NOR2_X1 U474 ( .A1(n585), .A2(n497), .ZN(n414) );
  NAND2_X1 U475 ( .A1(n555), .A2(n414), .ZN(n416) );
  XNOR2_X1 U476 ( .A(KEYINPUT37), .B(KEYINPUT99), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n531) );
  XOR2_X1 U478 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n418) );
  XNOR2_X1 U479 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U484 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n426) );
  NAND2_X1 U485 ( .A1(G230GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U487 ( .A(n428), .B(n427), .Z(n431) );
  XNOR2_X1 U488 ( .A(n429), .B(KEYINPUT32), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n577) );
  XOR2_X1 U490 ( .A(G22GAT), .B(G197GAT), .Z(n433) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(G113GAT), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n448) );
  XOR2_X1 U493 ( .A(n435), .B(n434), .Z(n437) );
  XNOR2_X1 U494 ( .A(G36GAT), .B(G50GAT), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U496 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n439) );
  NAND2_X1 U497 ( .A1(G229GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U499 ( .A(n441), .B(n440), .Z(n446) );
  XOR2_X1 U500 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n443) );
  XNOR2_X1 U501 ( .A(G141GAT), .B(G8GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n444), .B(KEYINPUT30), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n573) );
  NAND2_X1 U506 ( .A1(n577), .A2(n573), .ZN(n500) );
  XNOR2_X1 U507 ( .A(KEYINPUT38), .B(KEYINPUT100), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U509 ( .A1(n515), .A2(n537), .ZN(n455) );
  XOR2_X1 U510 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n453) );
  XNOR2_X1 U511 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n452) );
  NOR2_X1 U512 ( .A1(n555), .A2(n585), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n456), .B(KEYINPUT45), .ZN(n457) );
  NAND2_X1 U514 ( .A1(n457), .A2(n577), .ZN(n458) );
  NOR2_X1 U515 ( .A1(n573), .A2(n458), .ZN(n459) );
  XOR2_X1 U516 ( .A(n459), .B(KEYINPUT115), .Z(n467) );
  XOR2_X1 U517 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n461) );
  XNOR2_X1 U518 ( .A(n577), .B(KEYINPUT41), .ZN(n562) );
  NAND2_X1 U519 ( .A1(n562), .A2(n573), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(n463) );
  XOR2_X1 U521 ( .A(n555), .B(KEYINPUT112), .Z(n566) );
  NOR2_X1 U522 ( .A1(n557), .A2(n566), .ZN(n462) );
  NAND2_X1 U523 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U524 ( .A(KEYINPUT47), .B(n464), .ZN(n465) );
  XNOR2_X1 U525 ( .A(KEYINPUT114), .B(n465), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n535), .B(KEYINPUT123), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n483), .A2(n470), .ZN(n473) );
  XNOR2_X1 U529 ( .A(KEYINPUT54), .B(KEYINPUT124), .ZN(n471) );
  XOR2_X1 U530 ( .A(n471), .B(KEYINPUT125), .Z(n472) );
  XNOR2_X1 U531 ( .A(n473), .B(n472), .ZN(n569) );
  INV_X1 U532 ( .A(n533), .ZN(n570) );
  AND2_X1 U533 ( .A1(n570), .A2(n474), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n569), .A2(n475), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT55), .B(n476), .Z(n477) );
  NAND2_X1 U536 ( .A1(n567), .A2(n557), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n479) );
  INV_X1 U538 ( .A(G120GAT), .ZN(n491) );
  XNOR2_X1 U539 ( .A(KEYINPUT119), .B(KEYINPUT49), .ZN(n489) );
  NOR2_X1 U540 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U541 ( .A(n484), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U542 ( .A1(n549), .A2(n507), .ZN(n486) );
  NOR2_X1 U543 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U544 ( .A(n487), .B(KEYINPUT118), .ZN(n546) );
  AND2_X1 U545 ( .A1(n546), .A2(n562), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n491), .B(n490), .ZN(G1341GAT) );
  INV_X1 U548 ( .A(G127GAT), .ZN(n495) );
  XNOR2_X1 U549 ( .A(KEYINPUT50), .B(KEYINPUT120), .ZN(n493) );
  AND2_X1 U550 ( .A1(n566), .A2(n546), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n495), .B(n494), .ZN(G1342GAT) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n503) );
  NOR2_X1 U554 ( .A1(n557), .A2(n555), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(KEYINPUT16), .ZN(n499) );
  INV_X1 U556 ( .A(n497), .ZN(n498) );
  NAND2_X1 U557 ( .A1(n499), .A2(n498), .ZN(n519) );
  NOR2_X1 U558 ( .A1(n500), .A2(n519), .ZN(n501) );
  XOR2_X1 U559 ( .A(KEYINPUT97), .B(n501), .Z(n508) );
  NAND2_X1 U560 ( .A1(n533), .A2(n508), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(G1324GAT) );
  NAND2_X1 U562 ( .A1(n508), .A2(n535), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U564 ( .A(G15GAT), .B(KEYINPUT35), .Z(n506) );
  NAND2_X1 U565 ( .A1(n508), .A2(n537), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1326GAT) );
  INV_X1 U567 ( .A(n507), .ZN(n540) );
  NAND2_X1 U568 ( .A1(n508), .A2(n540), .ZN(n509) );
  XNOR2_X1 U569 ( .A(n509), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U570 ( .A1(n515), .A2(n533), .ZN(n511) );
  XOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT39), .Z(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U573 ( .A(KEYINPUT98), .B(n512), .ZN(G1328GAT) );
  NAND2_X1 U574 ( .A1(n515), .A2(n535), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n513), .B(KEYINPUT102), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G36GAT), .B(n514), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n540), .A2(n515), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G50GAT), .B(n516), .ZN(G1331GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT42), .B(KEYINPUT106), .Z(n521) );
  INV_X1 U580 ( .A(n573), .ZN(n517) );
  NAND2_X1 U581 ( .A1(n562), .A2(n517), .ZN(n518) );
  XOR2_X1 U582 ( .A(KEYINPUT105), .B(n518), .Z(n530) );
  NOR2_X1 U583 ( .A1(n530), .A2(n519), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n526), .A2(n533), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U586 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  XOR2_X1 U587 ( .A(G64GAT), .B(KEYINPUT107), .Z(n524) );
  NAND2_X1 U588 ( .A1(n526), .A2(n535), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1333GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n537), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U593 ( .A1(n526), .A2(n540), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G78GAT), .B(n529), .ZN(G1335GAT) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT109), .B(n532), .Z(n541) );
  NAND2_X1 U598 ( .A1(n533), .A2(n541), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n534), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n541), .A2(n535), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n541), .A2(n537), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(KEYINPUT110), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G99GAT), .B(n539), .ZN(G1338GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n543) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n544), .ZN(G1339GAT) );
  NAND2_X1 U609 ( .A1(n546), .A2(n573), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n545), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U612 ( .A1(n557), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  AND2_X1 U614 ( .A1(n549), .A2(n571), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n558), .A2(n573), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n552) );
  NAND2_X1 U618 ( .A1(n558), .A2(n562), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT53), .Z(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  INV_X1 U622 ( .A(n555), .ZN(n581) );
  NAND2_X1 U623 ( .A1(n581), .A2(n558), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT122), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n567), .A2(n573), .ZN(n561) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n561), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  NAND2_X1 U631 ( .A1(n567), .A2(n562), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  AND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n584) );
  INV_X1 U639 ( .A(n584), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n582), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n579) );
  OR2_X1 U644 ( .A1(n584), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n580), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

