//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT87), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT15), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT88), .ZN(new_n214));
  INV_X1    g013(.A(new_n212), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT15), .A3(new_n202), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT90), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(KEYINPUT17), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT17), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n214), .A2(new_n216), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n218), .A3(KEYINPUT17), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G15gat), .B(G22gat), .Z(new_n225));
  INV_X1    g024(.A(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228));
  AOI21_X1  g027(.A(G8gat), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(G1gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n231), .B2(new_n225), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n229), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n224), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n217), .A2(new_n233), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT18), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n235), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n217), .B(new_n233), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n237), .B(KEYINPUT92), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT13), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT91), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n239), .A2(new_n246), .A3(new_n243), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT11), .B(G169gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XOR2_X1   g048(.A(G113gat), .B(G141gat), .Z(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT86), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n252), .B(KEYINPUT12), .Z(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n247), .B(new_n254), .C1(new_n238), .C2(new_n244), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT22), .ZN(new_n262));
  NAND2_X1  g061(.A1(G211gat), .A2(G218gat), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n263), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n260), .B1(new_n272), .B2(KEYINPUT29), .ZN(new_n273));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  INV_X1    g073(.A(G155gat), .ZN(new_n275));
  INV_X1    g074(.A(G162gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G141gat), .B(G148gat), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n274), .B(new_n277), .C1(new_n278), .C2(KEYINPUT2), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT78), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n274), .B1(new_n277), .B2(KEYINPUT2), .ZN(new_n281));
  INV_X1    g080(.A(G141gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G148gat), .ZN(new_n283));
  INV_X1    g082(.A(G148gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G141gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n283), .B2(new_n285), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n274), .A4(new_n277), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n280), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n280), .A2(new_n260), .A3(new_n290), .A4(new_n286), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n272), .ZN(new_n296));
  AND2_X1   g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n295), .A2(KEYINPUT81), .A3(new_n272), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT81), .B1(new_n295), .B2(new_n272), .ZN(new_n300));
  INV_X1    g099(.A(new_n291), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT80), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n269), .A2(new_n302), .A3(new_n261), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(new_n294), .C1(new_n271), .C2(new_n302), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n304), .B2(new_n260), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n299), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n298), .B1(new_n306), .B2(new_n297), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT82), .B1(new_n307), .B2(G22gat), .ZN(new_n308));
  XOR2_X1   g107(.A(G78gat), .B(G106gat), .Z(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT31), .ZN(new_n310));
  INV_X1    g109(.A(G50gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G22gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n314), .B(new_n298), .C1(new_n306), .C2(new_n297), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n308), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n307), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n314), .C1(KEYINPUT82), .C2(new_n312), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n307), .A2(G22gat), .A3(new_n312), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT37), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n323));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G169gat), .ZN(new_n326));
  INV_X1    g125(.A(G176gat), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n327), .A2(KEYINPUT64), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(KEYINPUT64), .ZN(new_n329));
  OAI211_X1 g128(.A(KEYINPUT23), .B(new_n326), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT65), .B1(new_n331), .B2(KEYINPUT23), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT65), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n333), .B(new_n334), .C1(G169gat), .C2(G176gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  INV_X1    g140(.A(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n330), .A2(new_n336), .A3(new_n337), .A4(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT25), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(KEYINPUT67), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n340), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n338), .A2(KEYINPUT67), .A3(new_n339), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT69), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G183gat), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n353), .B1(new_n357), .B2(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n356), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(KEYINPUT69), .A3(new_n342), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n352), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n347), .B1(new_n332), .B2(new_n335), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT66), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT23), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n337), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n364), .A2(new_n363), .A3(new_n337), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n348), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n359), .A2(KEYINPUT27), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n341), .A2(KEYINPUT71), .A3(KEYINPUT27), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(KEYINPUT28), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT71), .B1(new_n341), .B2(KEYINPUT27), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n369), .A2(new_n371), .A3(new_n342), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n331), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n374), .A2(KEYINPUT26), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(KEYINPUT26), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n337), .A3(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(KEYINPUT27), .B(G183gat), .Z(new_n378));
  OAI21_X1  g177(.A(KEYINPUT28), .B1(new_n378), .B2(G190gat), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n373), .A2(new_n377), .A3(new_n338), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n368), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n325), .B1(new_n381), .B2(new_n294), .ZN(new_n382));
  INV_X1    g181(.A(new_n380), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(KEYINPUT67), .B2(new_n344), .ZN(new_n386));
  INV_X1    g185(.A(new_n351), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT69), .B1(new_n359), .B2(new_n342), .ZN(new_n389));
  AOI211_X1 g188(.A(new_n353), .B(G190gat), .C1(new_n354), .C2(new_n356), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n366), .A2(new_n365), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n362), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT70), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n348), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n383), .B1(new_n384), .B2(new_n395), .ZN(new_n396));
  OAI22_X1  g195(.A1(new_n323), .A2(new_n382), .B1(new_n396), .B2(new_n324), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n366), .A2(new_n365), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n336), .A2(KEYINPUT25), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI221_X4 g199(.A(KEYINPUT70), .B1(new_n346), .B2(new_n347), .C1(new_n400), .C2(new_n391), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n393), .B2(new_n348), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n380), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(KEYINPUT77), .A3(new_n325), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n272), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n324), .A2(new_n294), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n396), .A2(new_n406), .B1(new_n324), .B2(new_n381), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n272), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n322), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n397), .A2(new_n272), .A3(new_n404), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n411), .B(KEYINPUT37), .C1(new_n272), .C2(new_n407), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT38), .ZN(new_n413));
  XOR2_X1   g212(.A(G8gat), .B(G36gat), .Z(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G64gat), .ZN(new_n415));
  INV_X1    g214(.A(G92gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n410), .A2(new_n412), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT0), .B(G57gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(G85gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(G127gat), .B(G134gat), .Z(new_n424));
  OR2_X1    g223(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT1), .ZN(new_n427));
  XOR2_X1   g226(.A(G113gat), .B(G120gat), .Z(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n427), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n425), .A3(new_n424), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n301), .A2(new_n433), .A3(KEYINPUT4), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n291), .B2(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n432), .A3(new_n293), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT79), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n438), .A2(KEYINPUT79), .A3(new_n432), .A4(new_n293), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g243(.A1(G225gat), .A2(G233gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n291), .B(new_n432), .ZN(new_n448));
  INV_X1    g247(.A(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n445), .A2(new_n435), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n451), .B1(new_n443), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT6), .B(new_n423), .C1(new_n447), .C2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n423), .B1(new_n447), .B2(new_n454), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n442), .ZN(new_n457));
  INV_X1    g256(.A(new_n437), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(new_n452), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n422), .B(new_n446), .C1(new_n460), .C2(new_n451), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n417), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n405), .B2(new_n409), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n418), .A2(new_n455), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n397), .A2(new_n404), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n271), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n408), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n464), .B1(new_n469), .B2(new_n322), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(KEYINPUT37), .A3(new_n408), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n413), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n459), .A2(new_n473), .A3(new_n449), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT83), .B1(new_n443), .B2(new_n445), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(KEYINPUT84), .B(KEYINPUT39), .Z(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n448), .A2(new_n449), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT39), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n422), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n485), .A3(new_n464), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n408), .A3(new_n417), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(new_n465), .A3(KEYINPUT30), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n423), .B1(new_n476), .B2(new_n477), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT85), .B1(new_n490), .B2(new_n480), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n456), .B1(new_n491), .B2(new_n483), .ZN(new_n492));
  OAI221_X1 g291(.A(new_n321), .B1(new_n466), .B2(new_n472), .C1(new_n489), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(new_n486), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n463), .A2(new_n455), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n320), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT73), .ZN(new_n498));
  INV_X1    g297(.A(G227gat), .ZN(new_n499));
  INV_X1    g298(.A(G233gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n403), .A2(new_n432), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n384), .A2(new_n395), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(new_n433), .A3(new_n380), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n502), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n498), .B1(new_n506), .B2(KEYINPUT33), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n433), .B1(new_n504), .B2(new_n380), .ZN(new_n508));
  AOI211_X1 g307(.A(new_n432), .B(new_n383), .C1(new_n384), .C2(new_n395), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT33), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(KEYINPUT73), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(KEYINPUT32), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G43gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(G71gat), .ZN(new_n515));
  INV_X1    g314(.A(G99gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n507), .A2(new_n512), .A3(new_n513), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n517), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n511), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n502), .A3(new_n505), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n522), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n518), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT75), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n518), .A2(new_n521), .A3(KEYINPUT75), .A4(new_n525), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n518), .A2(new_n521), .ZN(new_n531));
  INV_X1    g330(.A(new_n525), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT76), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n534));
  AOI211_X1 g333(.A(new_n534), .B(new_n525), .C1(new_n518), .C2(new_n521), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT36), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n532), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n538), .A2(KEYINPUT36), .A3(new_n526), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n493), .B(new_n497), .C1(new_n537), .C2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n538), .A2(new_n494), .A3(new_n321), .A4(new_n526), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542));
  INV_X1    g341(.A(new_n495), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n496), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n530), .A2(new_n536), .A3(new_n545), .A4(new_n321), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n546), .B2(new_n542), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n259), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n549));
  INV_X1    g348(.A(G85gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(new_n416), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT8), .ZN(new_n552));
  AND2_X1   g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  OAI221_X1 g352(.A(new_n551), .B1(G85gat), .B2(G92gat), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n555));
  NOR4_X1   g354(.A1(new_n555), .A2(new_n549), .A3(new_n550), .A4(new_n416), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT97), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(KEYINPUT97), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  OR2_X1    g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G57gat), .B(G64gat), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n564), .A3(new_n565), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT94), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n563), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT10), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n563), .A2(new_n574), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n553), .A2(new_n558), .A3(KEYINPUT101), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n557), .B(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n570), .A3(new_n572), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT102), .B(KEYINPUT10), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n576), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(G230gat), .A2(G233gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n577), .B2(new_n580), .ZN(new_n588));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n327), .ZN(new_n590));
  INV_X1    g389(.A(G204gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OR3_X1    g391(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n587), .B2(new_n588), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n548), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n574), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n233), .B1(new_n574), .B2(new_n599), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(new_n341), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT95), .ZN(new_n606));
  INV_X1    g405(.A(G231gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(new_n500), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n605), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n608), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n264), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n609), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n609), .B2(new_n613), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n603), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n609), .A2(new_n613), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n615), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n609), .A2(new_n613), .A3(new_n616), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n602), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n217), .B2(new_n563), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n224), .B2(new_n563), .ZN(new_n627));
  XOR2_X1   g426(.A(G190gat), .B(G218gat), .Z(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n627), .A2(KEYINPUT98), .A3(new_n628), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT98), .B1(new_n627), .B2(new_n628), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT99), .B1(new_n630), .B2(new_n631), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  OAI221_X1 g437(.A(new_n629), .B1(KEYINPUT99), .B2(new_n638), .C1(new_n630), .C2(new_n631), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n598), .B1(new_n624), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n619), .A2(new_n623), .A3(KEYINPUT100), .A4(new_n640), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n597), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n495), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n226), .ZN(G1324gat));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n494), .ZN(new_n648));
  INV_X1    g447(.A(G8gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n230), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n230), .A2(new_n649), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n655), .B(new_n656), .C1(new_n649), .C2(new_n648), .ZN(G1325gat));
  INV_X1    g456(.A(G15gat), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n513), .A2(new_n520), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n503), .A2(new_n505), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT33), .B1(new_n660), .B2(new_n501), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n661), .A2(KEYINPUT73), .B1(KEYINPUT32), .B2(new_n510), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n510), .A2(new_n511), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n519), .B1(new_n663), .B2(new_n498), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n659), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n534), .B1(new_n665), .B2(new_n525), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n531), .A2(KEYINPUT76), .A3(new_n532), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n666), .A2(new_n528), .A3(new_n529), .A4(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT36), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n539), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n645), .A2(new_n658), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n668), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n597), .A2(new_n644), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n658), .B2(new_n674), .ZN(G1326gat));
  NOR2_X1   g474(.A1(new_n645), .A2(new_n321), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT43), .B(G22gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  NOR2_X1   g477(.A1(new_n640), .A2(KEYINPUT44), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n540), .A2(new_n547), .A3(KEYINPUT104), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT104), .B1(new_n540), .B2(new_n547), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n640), .B1(new_n540), .B2(new_n547), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n624), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n595), .B(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n687), .A2(new_n690), .A3(new_n259), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n206), .B1(new_n692), .B2(new_n543), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n687), .A2(new_n640), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n548), .A3(new_n596), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(new_n206), .A3(new_n543), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT45), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n697), .A2(KEYINPUT45), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n693), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n699), .A2(new_n698), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT105), .B1(new_n703), .B2(new_n693), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1328gat));
  INV_X1    g504(.A(new_n494), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n696), .A2(new_n207), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT46), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n207), .B1(new_n692), .B2(new_n706), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(G1329gat));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n686), .A2(new_n670), .A3(new_n691), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G43gat), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n695), .A2(G43gat), .A3(new_n668), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n715), .B1(new_n713), .B2(new_n714), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n711), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n718), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(KEYINPUT47), .A3(new_n716), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  INV_X1    g522(.A(new_n679), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n489), .A2(new_n492), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n321), .B1(new_n466), .B2(new_n472), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n497), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n670), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n538), .A2(new_n321), .A3(new_n526), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n731), .A2(KEYINPUT35), .A3(new_n495), .A4(new_n494), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n668), .A2(new_n320), .A3(new_n496), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(KEYINPUT35), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n725), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n540), .A2(new_n547), .A3(KEYINPUT104), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n724), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n683), .A2(new_n684), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n320), .B(new_n691), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT107), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n686), .A2(new_n741), .A3(new_n320), .A4(new_n691), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(G50gat), .A3(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n695), .A2(G50gat), .A3(new_n321), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n723), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  AOI211_X1 g545(.A(KEYINPUT48), .B(new_n744), .C1(new_n739), .C2(G50gat), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT108), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n747), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n311), .B1(new_n739), .B2(KEYINPUT107), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n744), .B1(new_n751), .B2(new_n742), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n749), .B(new_n750), .C1(new_n752), .C2(new_n723), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n748), .A2(new_n753), .ZN(G1331gat));
  AOI21_X1  g553(.A(new_n689), .B1(new_n735), .B2(new_n736), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n644), .A3(new_n259), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n495), .B(KEYINPUT109), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g559(.A1(new_n756), .A2(new_n494), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n756), .B2(new_n671), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n756), .A2(G71gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n668), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g568(.A1(new_n756), .A2(new_n321), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT110), .B(G78gat), .Z(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n687), .A2(new_n258), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n683), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT51), .Z(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(new_n595), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n550), .A3(new_n543), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n686), .A2(new_n595), .A3(new_n773), .ZN(new_n778));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n495), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1336gat));
  NOR3_X1   g579(.A1(new_n689), .A2(G92gat), .A3(new_n494), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G92gat), .B1(new_n778), .B2(new_n494), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n774), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n781), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(G1337gat));
  NAND3_X1  g589(.A1(new_n776), .A2(new_n516), .A3(new_n673), .ZN(new_n791));
  OAI21_X1  g590(.A(G99gat), .B1(new_n778), .B2(new_n671), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1338gat));
  AOI21_X1  g592(.A(new_n596), .B1(new_n682), .B2(new_n685), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n320), .A3(new_n773), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n794), .A2(KEYINPUT112), .A3(new_n320), .A4(new_n773), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(G106gat), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n689), .A2(G106gat), .A3(new_n321), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n775), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n795), .A2(G106gat), .B1(new_n786), .B2(new_n801), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n800), .B2(new_n804), .ZN(G1339gat));
  OAI21_X1  g604(.A(KEYINPUT54), .B1(new_n583), .B2(new_n585), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n587), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n592), .B1(new_n586), .B2(KEYINPUT54), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n587), .A2(new_n806), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n808), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n813), .A3(new_n593), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT113), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n810), .A2(new_n813), .A3(new_n816), .A4(new_n593), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n258), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n245), .A2(new_n253), .ZN(new_n819));
  INV_X1    g618(.A(new_n251), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n236), .A2(new_n237), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n240), .A2(new_n242), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n595), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n641), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n815), .A2(new_n817), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n819), .A2(new_n823), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n826), .A2(new_n640), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n624), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n642), .A2(new_n643), .A3(new_n596), .A4(new_n259), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n668), .A2(new_n320), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n706), .A2(new_n495), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n259), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n541), .B(new_n758), .C1(new_n829), .C2(new_n830), .ZN(new_n837));
  INV_X1    g636(.A(G113gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n838), .A3(new_n258), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n835), .B2(new_n689), .ZN(new_n841));
  INV_X1    g640(.A(G120gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n842), .A3(new_n595), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n835), .A2(new_n845), .A3(new_n624), .ZN(new_n846));
  AOI21_X1  g645(.A(G127gat), .B1(new_n837), .B2(new_n687), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(G1342gat));
  INV_X1    g647(.A(G134gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n837), .A2(new_n849), .A3(new_n641), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT114), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n835), .B2(new_n640), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n850), .A2(KEYINPUT114), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(KEYINPUT114), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(KEYINPUT56), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(G1343gat));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n831), .A2(new_n859), .A3(new_n320), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n671), .A2(new_n834), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT115), .B1(new_n812), .B2(new_n808), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT55), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT115), .B(new_n811), .C1(new_n812), .C2(new_n808), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n258), .A2(new_n593), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n641), .B1(new_n866), .B2(new_n824), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n624), .B1(new_n867), .B2(new_n828), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n321), .B1(new_n868), .B2(new_n830), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n860), .B(new_n862), .C1(new_n859), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G141gat), .B1(new_n870), .B2(new_n259), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n758), .B1(new_n829), .B2(new_n830), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n670), .A2(new_n321), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n873), .B2(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n258), .A2(new_n282), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT117), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n875), .A2(new_n878), .A3(new_n494), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n862), .B1(new_n869), .B2(new_n859), .ZN(new_n882));
  AOI211_X1 g681(.A(KEYINPUT57), .B(new_n321), .C1(new_n829), .C2(new_n830), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n882), .A2(new_n259), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n884), .B2(new_n282), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n872), .A2(new_n885), .A3(KEYINPUT58), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n871), .B(new_n881), .C1(KEYINPUT118), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1344gat));
  AND3_X1   g688(.A1(new_n875), .A2(new_n494), .A3(new_n878), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n890), .A2(KEYINPUT119), .A3(new_n284), .A4(new_n595), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n875), .A2(new_n878), .A3(new_n284), .A4(new_n494), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n596), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n859), .B1(new_n831), .B2(new_n320), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n320), .A2(new_n859), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n827), .A2(new_n640), .A3(new_n814), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n624), .B1(new_n867), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n899), .B2(new_n830), .ZN(new_n900));
  NOR4_X1   g699(.A1(new_n896), .A2(new_n900), .A3(new_n596), .A4(new_n861), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT59), .B1(new_n901), .B2(new_n284), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n870), .B2(new_n596), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n902), .B1(new_n284), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n895), .A2(new_n905), .ZN(G1345gat));
  NOR3_X1   g705(.A1(new_n870), .A2(new_n275), .A3(new_n624), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n687), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n275), .ZN(G1346gat));
  NOR3_X1   g708(.A1(new_n870), .A2(new_n276), .A3(new_n640), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n641), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n276), .ZN(G1347gat));
  AOI211_X1 g711(.A(new_n543), .B(new_n494), .C1(new_n829), .C2(new_n830), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n731), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n326), .A3(new_n258), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n757), .A2(new_n494), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n833), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n259), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(G1348gat));
  NOR4_X1   g718(.A1(new_n917), .A2(new_n328), .A3(new_n329), .A4(new_n689), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n914), .A2(new_n595), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n327), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(KEYINPUT120), .A3(new_n327), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n624), .A2(new_n378), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n913), .A2(new_n731), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n831), .A2(new_n687), .A3(new_n832), .A4(new_n916), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n357), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(KEYINPUT60), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1350gat));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n833), .A2(new_n641), .A3(new_n916), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(G190gat), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n941), .B2(G190gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n941), .A2(G190gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n943), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n914), .A2(new_n342), .A3(new_n641), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n949), .A3(new_n950), .ZN(G1351gat));
  XOR2_X1   g750(.A(KEYINPUT123), .B(G197gat), .Z(new_n952));
  NAND2_X1  g751(.A1(new_n913), .A2(new_n876), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n259), .ZN(new_n954));
  INV_X1    g753(.A(new_n916), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n896), .A2(new_n900), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n671), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n259), .A2(new_n952), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n954), .B(new_n961), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n831), .A2(new_n320), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n900), .B1(new_n964), .B2(KEYINPUT57), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n965), .A2(new_n671), .A3(new_n690), .A4(new_n916), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n956), .A2(KEYINPUT126), .A3(new_n671), .A4(new_n690), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(G204gat), .A3(new_n969), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n953), .A2(G204gat), .A3(new_n596), .ZN(new_n971));
  XOR2_X1   g770(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n972));
  OR2_X1    g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n970), .A2(new_n973), .A3(new_n975), .ZN(G1353gat));
  INV_X1    g775(.A(new_n953), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n264), .A3(new_n687), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n965), .A2(new_n687), .A3(new_n671), .A4(new_n916), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n957), .B2(new_n640), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n977), .A2(new_n265), .A3(new_n641), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


