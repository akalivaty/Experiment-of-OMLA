//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G58), .B2(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G77), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n203), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(G58), .A2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n206), .B(new_n227), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT67), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G222), .ZN(new_n263));
  INV_X1    g0063(.A(G223), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n261), .B(new_n263), .C1(new_n264), .C2(new_n262), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT68), .B1(new_n267), .B2(new_n228), .ZN(new_n268));
  INV_X1    g0068(.A(new_n228), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(new_n266), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n265), .B(new_n273), .C1(new_n220), .C2(new_n261), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n275), .B(G274), .C1(G41), .C2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n267), .A2(new_n228), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n278), .B1(G226), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n274), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G179), .ZN(new_n286));
  OAI21_X1  g0086(.A(G20), .B1(new_n232), .B2(G50), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n229), .A2(G33), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n287), .B1(new_n288), .B2(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n228), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n275), .A2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n213), .ZN(new_n300));
  INV_X1    g0100(.A(new_n295), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n297), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G50), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n296), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(G169), .B1(new_n274), .B2(new_n284), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n286), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n285), .A2(G200), .B1(new_n309), .B2(new_n305), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(KEYINPUT9), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n274), .A2(G190), .A3(new_n284), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n310), .A2(new_n315), .A3(new_n311), .A4(new_n312), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n308), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n303), .A2(G68), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT74), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n229), .A2(G33), .A3(G77), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n301), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n322), .A2(KEYINPUT11), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(KEYINPUT11), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT12), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT75), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n325), .A2(KEYINPUT75), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n299), .A2(new_n217), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n319), .A2(new_n323), .A3(new_n324), .A4(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n326), .B1(new_n299), .B2(new_n217), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n214), .A2(new_n262), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n237), .A2(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n261), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n272), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n276), .B(KEYINPUT66), .ZN(new_n338));
  INV_X1    g0138(.A(new_n283), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n218), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n332), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n278), .B1(G238), .B2(new_n283), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n256), .A2(new_n260), .B1(new_n237), .B2(G1698), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n333), .B1(G33), .B2(G97), .ZN(new_n344));
  OAI211_X1 g0144(.A(KEYINPUT13), .B(new_n342), .C1(new_n344), .C2(new_n272), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n341), .A2(new_n345), .A3(G200), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n332), .A2(KEYINPUT73), .ZN(new_n347));
  OR3_X1    g0147(.A1(new_n337), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n337), .B2(new_n340), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(G190), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n331), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n341), .A2(new_n345), .A3(G169), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(new_n349), .A3(G179), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n341), .A2(new_n345), .A3(new_n355), .A4(G169), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n331), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n317), .A2(new_n351), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT7), .A2(G20), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT76), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G33), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n252), .A2(KEYINPUT76), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT3), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n366), .B2(new_n257), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n252), .A2(KEYINPUT76), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(G33), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n254), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n370), .A2(KEYINPUT77), .A3(new_n253), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n361), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n370), .A2(new_n253), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT7), .B1(new_n373), .B2(G20), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(G68), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(G58), .B(G68), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(KEYINPUT16), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT76), .B(G33), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n255), .B1(new_n379), .B2(new_n254), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT7), .B1(new_n380), .B2(G20), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n256), .A2(new_n260), .A3(new_n361), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(G68), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n377), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT16), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n378), .A2(new_n295), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n299), .ZN(new_n388));
  MUX2_X1   g0188(.A(new_n302), .B(new_n388), .S(new_n291), .Z(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G223), .A2(G1698), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n262), .A2(G226), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n366), .A2(new_n257), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n252), .A2(new_n207), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n272), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n338), .B1(new_n339), .B2(new_n237), .ZN(new_n400));
  OAI21_X1  g0200(.A(G169), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR4_X1   g0201(.A1(new_n370), .A2(new_n253), .A3(new_n392), .A4(new_n394), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n273), .B1(new_n402), .B2(new_n397), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n278), .B1(G232), .B2(new_n283), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(G179), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT18), .B1(new_n391), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n404), .ZN(new_n409));
  INV_X1    g0209(.A(G200), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(G190), .B2(new_n409), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n387), .A2(new_n389), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT17), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n390), .A2(new_n415), .A3(new_n406), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n387), .A2(new_n389), .A3(new_n412), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n408), .A2(new_n414), .A3(new_n416), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n262), .A2(G232), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n261), .B(new_n421), .C1(new_n218), .C2(new_n262), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n422), .B(new_n273), .C1(G107), .C2(new_n261), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n278), .B1(G244), .B2(new_n283), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G169), .ZN(new_n426));
  INV_X1    g0226(.A(G77), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n302), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n388), .A2(new_n220), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n220), .A2(G20), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT69), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n291), .B(new_n433), .ZN(new_n434));
  XOR2_X1   g0234(.A(new_n289), .B(KEYINPUT70), .Z(new_n435));
  OAI221_X1 g0235(.A(new_n430), .B1(new_n292), .B2(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  AOI211_X1 g0236(.A(new_n428), .B(new_n429), .C1(new_n436), .C2(new_n295), .ZN(new_n437));
  OR3_X1    g0237(.A1(new_n426), .A2(KEYINPUT71), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n425), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT71), .B1(new_n426), .B2(new_n437), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n425), .A2(G190), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n437), .C1(new_n410), .C2(new_n425), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n445), .A2(KEYINPUT72), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(KEYINPUT72), .ZN(new_n447));
  AOI211_X1 g0247(.A(new_n360), .B(new_n420), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n207), .A2(G20), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n261), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT22), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT24), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n368), .A2(new_n369), .A3(new_n229), .A4(G116), .ZN(new_n454));
  OR3_X1    g0254(.A1(new_n229), .A2(KEYINPUT23), .A3(G107), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT23), .B1(new_n229), .B2(G107), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n366), .A2(KEYINPUT22), .A3(new_n257), .A4(new_n449), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n452), .A2(new_n453), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n449), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n256), .B2(new_n260), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n457), .B(new_n458), .C1(new_n461), .C2(KEYINPUT22), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT24), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n301), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n208), .A2(new_n262), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n224), .A2(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n366), .A2(new_n257), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n379), .A2(G294), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n273), .ZN(new_n471));
  INV_X1    g0271(.A(G190), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n281), .A2(G1), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n269), .A2(new_n266), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n210), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n471), .A2(new_n472), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n272), .B1(new_n468), .B2(new_n469), .ZN(new_n484));
  INV_X1    g0284(.A(new_n482), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n484), .A2(new_n479), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n483), .B1(new_n486), .B2(G200), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n295), .B1(new_n275), .B2(G33), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n388), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n209), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n299), .A2(new_n209), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT25), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n465), .A2(new_n487), .A3(new_n491), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n464), .A2(new_n490), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n486), .A2(new_n439), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n486), .B2(G169), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT79), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n219), .A2(G1698), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G238), .B2(G1698), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n366), .A3(new_n257), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n379), .A2(G116), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n272), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n473), .A2(new_n481), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n208), .B1(new_n281), .B2(G1), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n477), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n507), .A2(new_n439), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G169), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n370), .A2(new_n503), .A3(new_n253), .ZN(new_n514));
  INV_X1    g0314(.A(new_n506), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n273), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n501), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(G169), .B1(new_n507), .B2(new_n511), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(G179), .A3(new_n510), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT79), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n229), .B1(new_n336), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G97), .A2(G107), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n207), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n522), .B1(new_n292), .B2(new_n223), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n229), .B(new_n257), .C1(new_n379), .C2(new_n254), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n217), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(new_n295), .B1(new_n299), .B2(new_n432), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT80), .B1(new_n489), .B2(new_n432), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n488), .A2(new_n532), .A3(new_n388), .A4(new_n431), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n518), .A2(new_n521), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(G200), .B1(new_n507), .B2(new_n511), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n488), .A2(G87), .A3(new_n388), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT81), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n516), .A2(G190), .A3(new_n510), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n537), .A2(new_n539), .A3(new_n530), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n496), .A2(new_n500), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n368), .A2(new_n369), .A3(new_n254), .ZN(new_n544));
  AOI21_X1  g0344(.A(G20), .B1(new_n544), .B2(new_n258), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT7), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n382), .B(G107), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n550));
  XOR2_X1   g0350(.A(G97), .B(G107), .Z(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(KEYINPUT6), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n381), .A2(KEYINPUT78), .A3(G107), .A4(new_n382), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n295), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n299), .A2(new_n223), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n489), .B2(new_n223), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n561));
  OAI211_X1 g0361(.A(G244), .B(new_n257), .C1(new_n379), .C2(new_n254), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT4), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(G33), .B2(G283), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n260), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n259), .B1(new_n257), .B2(new_n258), .ZN(new_n567));
  OAI21_X1  g0367(.A(G250), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n262), .B1(new_n568), .B2(KEYINPUT4), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n273), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n482), .B1(new_n224), .B2(new_n478), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n513), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n563), .B1(new_n261), .B2(G250), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n564), .B(new_n561), .C1(new_n575), .C2(new_n262), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n571), .B1(new_n576), .B2(new_n273), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n439), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n560), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G116), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n299), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n488), .A2(G116), .A3(new_n388), .ZN(new_n582));
  AOI21_X1  g0382(.A(G20), .B1(G33), .B2(G283), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(G33), .B2(new_n223), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n584), .B(new_n295), .C1(new_n229), .C2(G116), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n581), .B(new_n582), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G169), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G257), .A2(G1698), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n210), .A2(G1698), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n373), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n256), .A2(G303), .A3(new_n260), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n272), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n478), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G270), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n596), .A2(new_n485), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT21), .B1(new_n590), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n273), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n482), .A3(new_n598), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(G169), .A4(new_n589), .ZN(new_n606));
  INV_X1    g0406(.A(new_n589), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n601), .A2(new_n606), .B1(new_n608), .B2(G179), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n558), .B1(new_n555), .B2(new_n295), .ZN(new_n610));
  AOI211_X1 g0410(.A(G190), .B(new_n571), .C1(new_n576), .C2(new_n273), .ZN(new_n611));
  AOI21_X1  g0411(.A(G200), .B1(new_n570), .B2(new_n572), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n600), .A2(G190), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(new_n607), .C1(new_n410), .C2(new_n600), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n579), .A2(new_n609), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n448), .A2(new_n543), .A3(new_n616), .ZN(G372));
  OAI21_X1  g0417(.A(new_n535), .B1(new_n517), .B2(new_n512), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n541), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n579), .A2(new_n613), .A3(new_n495), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT82), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n541), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n497), .B2(new_n487), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT82), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n579), .A4(new_n613), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n465), .A2(new_n491), .A3(new_n494), .ZN(new_n626));
  INV_X1    g0426(.A(new_n499), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n609), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT26), .B1(new_n579), .B2(new_n542), .ZN(new_n631));
  AOI21_X1  g0431(.A(G169), .B1(new_n570), .B2(new_n572), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n439), .B2(new_n577), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n633), .A2(new_n619), .A3(new_n634), .A4(new_n560), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n631), .A2(new_n618), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n448), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n442), .A2(new_n359), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n351), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n414), .A2(new_n419), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n408), .B(new_n416), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n314), .A2(new_n316), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n308), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(new_n644), .ZN(G369));
  NOR2_X1   g0445(.A1(new_n298), .A2(G20), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .A3(G1), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT27), .B1(new_n647), .B2(G1), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n607), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n609), .A2(KEYINPUT83), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT83), .B1(new_n609), .B2(new_n655), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n609), .A2(new_n615), .A3(new_n655), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G330), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT85), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT85), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n660), .A2(new_n665), .A3(G330), .A4(new_n661), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n626), .A2(new_n627), .A3(new_n652), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT86), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n628), .B(new_n495), .C1(new_n497), .C2(new_n653), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(KEYINPUT86), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n609), .A2(new_n652), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n500), .A2(new_n653), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n673), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n204), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n525), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT87), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT87), .ZN(new_n686));
  INV_X1    g0486(.A(new_n234), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n685), .B(new_n686), .C1(new_n687), .C2(new_n682), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n652), .B1(new_n630), .B2(new_n636), .ZN(new_n690));
  OR3_X1    g0490(.A1(new_n690), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n579), .A2(new_n613), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n629), .A3(new_n623), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT26), .B1(new_n579), .B2(new_n622), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n579), .A2(new_n542), .A3(KEYINPUT26), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n618), .B(KEYINPUT90), .Z(new_n696));
  NAND4_X1  g0496(.A1(new_n693), .A2(new_n694), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .A3(new_n653), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT89), .B1(new_n690), .B2(KEYINPUT29), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n691), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n616), .A2(new_n543), .A3(new_n653), .ZN(new_n701));
  NOR4_X1   g0501(.A1(new_n577), .A2(new_n600), .A3(G179), .A4(new_n486), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n507), .B2(new_n511), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n577), .A2(new_n512), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n600), .A2(new_n471), .A3(new_n480), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT88), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(KEYINPUT30), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n704), .B2(new_n705), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n703), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n652), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n711), .A2(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n700), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n689), .B1(new_n717), .B2(G1), .ZN(G364));
  AOI21_X1  g0518(.A(new_n275), .B1(new_n646), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n681), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(G330), .B1(new_n660), .B2(new_n661), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n667), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n229), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n662), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n228), .B1(G20), .B2(new_n513), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n229), .A2(new_n439), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n472), .A2(new_n410), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT92), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT92), .B1(new_n730), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n730), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n736), .A2(G190), .A3(G200), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n735), .A2(G326), .B1(G311), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G294), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n472), .A2(G179), .A3(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n229), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n738), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT95), .Z(new_n743));
  NOR2_X1   g0543(.A1(new_n229), .A2(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n472), .A3(new_n410), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G329), .ZN(new_n747));
  INV_X1    g0547(.A(G322), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n736), .A2(new_n472), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT91), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n743), .B(new_n747), .C1(new_n748), .C2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n736), .A2(new_n410), .A3(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n744), .A2(new_n472), .A3(G200), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT93), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(KEYINPUT93), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT94), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n731), .A2(new_n744), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n261), .B1(G303), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT96), .Z(new_n771));
  NOR4_X1   g0571(.A1(new_n755), .A2(new_n759), .A3(new_n767), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n765), .A2(new_n209), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n768), .A2(new_n207), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n737), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n775), .B(new_n261), .C1(new_n221), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n746), .A2(G159), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n735), .A2(G50), .B1(KEYINPUT32), .B2(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n779), .B1(KEYINPUT32), .B2(new_n778), .C1(new_n217), .C2(new_n757), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n741), .A2(new_n223), .ZN(new_n781));
  INV_X1    g0581(.A(G58), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n754), .A2(new_n782), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n777), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n729), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n366), .A2(new_n257), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT77), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n373), .A2(new_n362), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n680), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n234), .A2(new_n281), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(new_n281), .C2(new_n247), .ZN(new_n793));
  INV_X1    g0593(.A(G355), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n261), .A2(new_n204), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n793), .B1(G116), .B2(new_n204), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n727), .A2(new_n729), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g0598(.A1(new_n728), .A2(new_n785), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n724), .B1(new_n722), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT97), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  INV_X1    g0602(.A(new_n445), .ZN(new_n803));
  AND4_X1   g0603(.A1(KEYINPUT99), .A2(new_n637), .A3(new_n803), .A4(new_n653), .ZN(new_n804));
  AOI21_X1  g0604(.A(KEYINPUT99), .B1(new_n690), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n437), .A2(new_n653), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n442), .A2(new_n444), .A3(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n438), .A2(new_n440), .A3(new_n441), .A4(new_n806), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n804), .A2(new_n805), .B1(new_n690), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(new_n716), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n722), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n735), .A2(G137), .B1(G159), .B2(new_n737), .ZN(new_n814));
  INV_X1    g0614(.A(G143), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n288), .B2(new_n757), .C1(new_n754), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT34), .ZN(new_n817));
  INV_X1    g0617(.A(new_n741), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G58), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n764), .A2(G68), .B1(G50), .B2(new_n769), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n817), .A2(new_n790), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G132), .B2(new_n746), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n754), .A2(new_n739), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n781), .B(new_n823), .C1(G87), .C2(new_n764), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n776), .A2(new_n580), .B1(new_n768), .B2(new_n209), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n261), .B(new_n825), .C1(G311), .C2(new_n746), .ZN(new_n826));
  INV_X1    g0626(.A(G303), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n824), .B(new_n826), .C1(new_n827), .C2(new_n734), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G283), .B2(new_n756), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n729), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n729), .A2(new_n725), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT98), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n725), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n830), .B1(G77), .B2(new_n833), .C1(new_n834), .C2(new_n810), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n721), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n813), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n837), .A2(KEYINPUT100), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(KEYINPUT100), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  INV_X1    g0641(.A(KEYINPUT39), .ZN(new_n842));
  XNOR2_X1  g0642(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT106), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n401), .A2(new_n405), .A3(new_n650), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n387), .B2(new_n389), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n413), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT103), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT103), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n413), .A2(new_n847), .A3(new_n851), .A4(KEYINPUT37), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n845), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT37), .B1(new_n413), .B2(new_n847), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n849), .B(new_n417), .C1(new_n391), .C2(new_n846), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n851), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n848), .A2(KEYINPUT103), .A3(new_n849), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT106), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n853), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n650), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n420), .A2(new_n390), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n844), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n378), .A2(new_n295), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n375), .A2(new_n377), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(KEYINPUT16), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n389), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n407), .A2(new_n650), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n413), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n850), .A2(new_n852), .B1(new_n868), .B2(new_n849), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n420), .A2(new_n860), .A3(new_n866), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT38), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n842), .B1(new_n862), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n357), .A2(new_n358), .A3(new_n653), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT104), .Z(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n869), .A2(new_n870), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n873), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n442), .A2(new_n652), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n804), .B2(new_n805), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n358), .A2(new_n652), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n359), .A2(new_n351), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT102), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n357), .A2(new_n358), .A3(new_n652), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n879), .A2(new_n871), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n884), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n408), .A2(new_n416), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n650), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n881), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n691), .A2(new_n448), .A3(new_n698), .A4(new_n699), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n644), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n897), .B(new_n899), .Z(new_n900));
  OAI21_X1  g0700(.A(new_n810), .B1(new_n889), .B2(new_n890), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n714), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n862), .B2(new_n872), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n714), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n903), .A2(KEYINPUT40), .B1(new_n893), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n448), .A2(new_n715), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n905), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(G330), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n900), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n275), .B2(new_n646), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n580), .B1(new_n552), .B2(KEYINPUT35), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n230), .C1(KEYINPUT35), .C2(new_n552), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n217), .A2(G50), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT101), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n220), .B1(new_n782), .B2(new_n217), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(new_n687), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n298), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n913), .A3(new_n918), .ZN(G367));
  INV_X1    g0719(.A(new_n673), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n692), .B1(new_n610), .B2(new_n653), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n633), .A2(new_n560), .A3(new_n652), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT109), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n923), .ZN(new_n927));
  OR3_X1    g0727(.A1(new_n675), .A2(new_n927), .A3(KEYINPUT42), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n579), .B1(new_n921), .B2(new_n628), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n653), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT42), .B1(new_n675), .B2(new_n927), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n539), .A2(new_n530), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n652), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT107), .B1(new_n619), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n618), .A2(new_n935), .ZN(new_n937));
  MUX2_X1   g0737(.A(new_n936), .B(KEYINPUT107), .S(new_n937), .Z(new_n938));
  INV_X1    g0738(.A(KEYINPUT43), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n938), .A2(new_n939), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n933), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n933), .A2(new_n941), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n926), .B(new_n943), .C1(new_n944), .C2(new_n940), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n924), .A2(new_n925), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n681), .B(KEYINPUT41), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n675), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n672), .A2(new_n674), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n667), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n717), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT111), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n678), .A2(KEYINPUT110), .A3(new_n923), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT44), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT110), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n677), .B2(new_n927), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n677), .A2(new_n927), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT45), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n958), .B1(new_n957), .B2(new_n960), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(new_n920), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n953), .A2(KEYINPUT111), .A3(new_n717), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n920), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n956), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n949), .B1(new_n969), .B2(new_n717), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n947), .B1(new_n970), .B2(new_n720), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n797), .B1(new_n432), .B2(new_n204), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n791), .B2(new_n243), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n776), .A2(new_n213), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n261), .B1(new_n763), .B2(new_n221), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G159), .B2(new_n756), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n741), .A2(new_n217), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n815), .B2(new_n734), .C1(new_n754), .C2(new_n288), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n976), .B1(new_n979), .B2(KEYINPUT112), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n974), .B(new_n980), .C1(KEYINPUT112), .C2(new_n979), .ZN(new_n981));
  INV_X1    g0781(.A(G137), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n981), .B1(new_n782), .B2(new_n768), .C1(new_n982), .C2(new_n745), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n776), .A2(new_n766), .ZN(new_n984));
  INV_X1    g0784(.A(new_n754), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n985), .A2(G303), .B1(G107), .B2(new_n818), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n769), .A2(G116), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(new_n988), .A3(new_n789), .ZN(new_n989));
  INV_X1    g0789(.A(new_n763), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n989), .B1(G97), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n746), .A2(G317), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n735), .A2(G311), .B1(G294), .B2(new_n756), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n983), .B1(new_n984), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n973), .B1(new_n996), .B2(new_n729), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n938), .A2(new_n727), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n721), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n971), .A2(new_n999), .ZN(G387));
  NAND2_X1  g0800(.A1(new_n956), .A2(new_n967), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1001), .B(new_n681), .C1(new_n717), .C2(new_n953), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n434), .A2(G50), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(G68), .A2(G77), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1004), .A2(new_n281), .A3(new_n1005), .A4(new_n683), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n791), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n240), .B2(G45), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n795), .A2(new_n683), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(G107), .B2(new_n204), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(new_n797), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n985), .A2(G317), .B1(G311), .B2(new_n756), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n827), .B2(new_n776), .C1(new_n748), .C2(new_n734), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT48), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n766), .B2(new_n741), .C1(new_n739), .C2(new_n768), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT49), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n790), .B1(G326), .B2(new_n746), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n580), .C2(new_n763), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n789), .B1(G150), .B2(new_n746), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n291), .B2(new_n757), .C1(new_n432), .C2(new_n741), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n754), .A2(new_n213), .B1(new_n221), .B2(new_n768), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G68), .C2(new_n737), .ZN(new_n1023));
  INV_X1    g0823(.A(G159), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1023), .B1(new_n223), .B2(new_n765), .C1(new_n1024), .C2(new_n734), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n722), .B(new_n1012), .C1(new_n1026), .C2(new_n729), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n672), .A2(new_n726), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1027), .A2(new_n1028), .B1(new_n720), .B2(new_n953), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1002), .A2(new_n1029), .ZN(G393));
  NAND3_X1  g0830(.A1(new_n966), .A2(new_n720), .A3(new_n968), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n434), .A2(new_n776), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n754), .A2(new_n1024), .B1(new_n734), .B2(new_n288), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT51), .Z(new_n1034));
  OAI22_X1  g0834(.A1(new_n745), .A2(new_n815), .B1(new_n768), .B2(new_n217), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n741), .A2(new_n427), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n790), .C1(new_n207), .C2(new_n765), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1032), .B(new_n1038), .C1(G50), .C2(new_n756), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n776), .A2(new_n739), .B1(new_n757), .B2(new_n827), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G116), .B2(new_n818), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(KEYINPUT113), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n261), .B(new_n773), .C1(KEYINPUT113), .C2(new_n1041), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n985), .A2(G311), .B1(G317), .B2(new_n735), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT52), .Z(new_n1045));
  OAI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(new_n748), .C2(new_n745), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1042), .B(new_n1046), .C1(G283), .C2(new_n769), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n729), .B1(new_n1039), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n927), .A2(new_n727), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n797), .B1(new_n223), .B2(new_n204), .C1(new_n1007), .C2(new_n250), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1048), .A2(new_n721), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1031), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n966), .A2(new_n968), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n682), .B1(new_n1001), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1052), .B1(new_n1054), .B2(new_n969), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(G390));
  NAND4_X1  g0856(.A1(new_n712), .A2(new_n713), .A3(G330), .A4(new_n810), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1057), .A2(new_n891), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n884), .A2(new_n892), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1060), .A2(new_n875), .B1(new_n873), .B2(new_n880), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n697), .A2(new_n810), .A3(new_n653), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n883), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n892), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n875), .B(KEYINPUT114), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n872), .C2(new_n862), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1059), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n637), .A2(new_n803), .A3(new_n653), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT99), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n690), .A2(KEYINPUT99), .A3(new_n803), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n882), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n875), .B1(new_n1073), .B2(new_n891), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n873), .A2(new_n880), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n1066), .A3(new_n1058), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1068), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n834), .B1(new_n873), .B2(new_n880), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n832), .A2(new_n291), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT54), .B(G143), .Z(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(G125), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n776), .A2(new_n1082), .B1(new_n1083), .B2(new_n745), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n985), .A2(G132), .B1(G159), .B2(new_n818), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n768), .A2(new_n288), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT53), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n756), .A2(G137), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1087), .A3(new_n261), .A4(new_n1088), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1084), .B(new_n1089), .C1(G50), .C2(new_n990), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n735), .A2(G128), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n756), .A2(G107), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n261), .B1(new_n985), .B2(G116), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n764), .A2(G68), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n746), .A2(G294), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n774), .B(new_n1036), .C1(G97), .C2(new_n737), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G283), .B2(new_n735), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1090), .A2(new_n1091), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT116), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n729), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n721), .B(new_n1080), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1078), .A2(new_n719), .B1(new_n1079), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n448), .A2(G330), .A3(new_n715), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n898), .A2(new_n644), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1057), .A2(new_n891), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1058), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n884), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1058), .A2(new_n883), .A3(new_n1062), .A4(new_n1106), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1061), .A2(new_n1067), .A3(new_n1059), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1058), .B1(new_n1076), .B2(new_n1066), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1068), .A2(new_n1077), .A3(new_n1110), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n681), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT115), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(KEYINPUT115), .A3(new_n681), .A4(new_n1115), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1103), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(G378));
  INV_X1    g0921(.A(new_n1105), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1115), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n897), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n308), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n643), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT55), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT55), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n317), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n306), .A2(new_n650), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1128), .B1(new_n643), .B2(new_n1125), .ZN(new_n1133));
  AOI211_X1 g0933(.A(KEYINPUT55), .B(new_n308), .C1(new_n314), .C2(new_n316), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1132), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n904), .A2(new_n893), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(G330), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT119), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1137), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1136), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1131), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1133), .A2(new_n1134), .A3(new_n1130), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1132), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT119), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n905), .A2(new_n663), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1124), .B1(new_n1143), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1152), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1142), .A2(new_n1155), .A3(G330), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n905), .A2(new_n663), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n1157), .A3(new_n897), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT57), .B1(new_n1123), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1123), .A2(new_n1159), .A3(KEYINPUT57), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n681), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n720), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1155), .A2(new_n725), .ZN(new_n1165));
  INV_X1    g0965(.A(G124), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n252), .B1(new_n745), .B2(new_n1166), .ZN(new_n1167));
  OR3_X1    g0967(.A1(new_n1082), .A2(KEYINPUT117), .A3(new_n768), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT117), .B1(new_n1082), .B2(new_n768), .ZN(new_n1169));
  INV_X1    g0969(.A(G132), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1169), .C1(new_n1170), .C2(new_n757), .ZN(new_n1171));
  INV_X1    g0971(.A(G128), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n754), .A2(new_n1172), .B1(new_n288), .B2(new_n741), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G137), .C2(new_n737), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1083), .B2(new_n734), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G41), .B(new_n1167), .C1(new_n1175), .C2(KEYINPUT59), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(KEYINPUT59), .B2(new_n1175), .C1(new_n1024), .C2(new_n763), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(new_n790), .B2(G33), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1177), .B1(G50), .B2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n985), .A2(G107), .B1(G58), .B2(new_n990), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n580), .B2(new_n734), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n978), .B1(new_n766), .B2(new_n745), .C1(new_n757), .C2(new_n223), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1181), .A2(G41), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n790), .B1(new_n220), .B2(new_n769), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n432), .C2(new_n776), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT58), .Z(new_n1186));
  OAI21_X1  g0986(.A(new_n729), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n831), .A2(new_n213), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1165), .A2(new_n721), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1164), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1163), .A2(new_n1191), .ZN(G375));
  AND2_X1   g0992(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n833), .A2(G68), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n985), .A2(G283), .B1(new_n431), .B2(new_n818), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n776), .A2(new_n209), .B1(new_n768), .B2(new_n223), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n261), .B(new_n1196), .C1(G303), .C2(new_n746), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n735), .A2(G294), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n764), .A2(G77), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G116), .B2(new_n756), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n990), .A2(G58), .B1(G159), .B2(new_n769), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n213), .B2(new_n741), .C1(new_n982), .C2(new_n754), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n790), .B1(new_n1170), .B2(new_n734), .C1(new_n757), .C2(new_n1082), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n745), .A2(new_n1172), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n776), .A2(new_n288), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n729), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n721), .B(new_n1208), .C1(new_n892), .C2(new_n834), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1193), .A2(new_n719), .B1(new_n1194), .B2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT120), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1193), .A2(new_n1105), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(new_n1111), .A3(new_n948), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(G381));
  INV_X1    g1014(.A(G375), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1103), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1216), .A2(new_n1116), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(G381), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n971), .A2(new_n999), .A3(new_n1055), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(G393), .A2(G396), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n840), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT121), .Z(new_n1224));
  NAND3_X1  g1024(.A1(new_n1219), .A2(new_n1221), .A3(new_n1224), .ZN(G407));
  NAND2_X1  g1025(.A1(new_n651), .A2(G213), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT122), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(G407), .B(G213), .C1(new_n1218), .C2(new_n1228), .ZN(G409));
  NAND2_X1  g1029(.A1(new_n1212), .A2(KEYINPUT124), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n681), .B(new_n1111), .C1(new_n1230), .C2(KEYINPUT60), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1230), .A2(KEYINPUT60), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1211), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(G384), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1211), .B(new_n840), .C1(new_n1232), .C2(new_n1231), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1123), .A2(new_n1159), .A3(KEYINPUT57), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1237), .A2(new_n1160), .A3(new_n682), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1238), .A2(new_n1120), .A3(new_n1190), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT123), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1159), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1154), .A2(KEYINPUT123), .A3(new_n1158), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n720), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1123), .A2(new_n1159), .A3(new_n948), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1189), .A3(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1245), .A2(new_n1217), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1228), .B(new_n1236), .C1(new_n1239), .C2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(new_n1217), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(G375), .B2(new_n1120), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1248), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n1228), .A3(new_n1236), .A4(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1250), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1227), .A2(G2897), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1236), .B(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1252), .A2(new_n1228), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT61), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1255), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1055), .B1(new_n971), .B2(new_n999), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n801), .B1(new_n1002), .B2(new_n1029), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1222), .A2(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1265), .A2(new_n1220), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1265), .B2(new_n1220), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1255), .A2(KEYINPUT127), .A3(new_n1260), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1263), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1247), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1252), .A2(KEYINPUT63), .A3(new_n1228), .A4(new_n1236), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1278), .A2(KEYINPUT125), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(KEYINPUT125), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1275), .B(new_n1276), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1272), .A2(new_n1281), .ZN(G405));
  AOI21_X1  g1082(.A(new_n1239), .B1(G375), .B2(new_n1217), .ZN(new_n1283));
  XOR2_X1   g1083(.A(new_n1283), .B(new_n1236), .Z(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1270), .ZN(G402));
endmodule


