//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n209), .B1(new_n213), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(KEYINPUT3), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G223), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n249), .B1(new_n250), .B2(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n210), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  AND2_X1   g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n260), .A2(new_n259), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT67), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n267), .A2(new_n268), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n262), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G226), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n256), .A2(G190), .A3(new_n270), .A4(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT71), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n256), .A2(new_n270), .A3(new_n278), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n210), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT68), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT68), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n288), .A3(new_n210), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n260), .A2(G13), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n211), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT69), .B1(new_n211), .B2(G1), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT69), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(new_n260), .A3(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(G50), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT8), .B(G58), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n211), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G150), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n299), .A2(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G50), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n211), .B1(new_n201), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n290), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G13), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G1), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G20), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n298), .B(new_n307), .C1(G50), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT9), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n311), .B(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT10), .B1(new_n284), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n311), .B(KEYINPUT9), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n283), .A4(new_n281), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n282), .A2(G179), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n282), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n311), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n286), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n245), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n246), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT73), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n332), .A2(KEYINPUT73), .A3(KEYINPUT7), .A4(new_n211), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n245), .A2(new_n211), .A3(new_n246), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n329), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G68), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n216), .ZN(new_n340));
  OAI21_X1  g0140(.A(G20), .B1(new_n340), .B2(new_n201), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n302), .A2(G159), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT16), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n326), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n216), .B1(new_n336), .B2(new_n327), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n344), .B1(new_n347), .B2(new_n343), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n344), .C1(new_n347), .C2(new_n343), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n346), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n299), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n297), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT75), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT75), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n297), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n293), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n292), .A2(new_n299), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n265), .A2(new_n269), .B1(new_n271), .B2(G232), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n252), .A2(new_n248), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G1698), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(new_n366), .C1(new_n330), .C2(new_n331), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G87), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n274), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n363), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n271), .A2(G232), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n270), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n321), .B1(new_n375), .B2(new_n369), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT76), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n363), .A2(new_n370), .A3(new_n377), .A4(new_n371), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n373), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n362), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT18), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n379), .B1(new_n352), .B2(new_n361), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT18), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n375), .A2(new_n369), .ZN(new_n386));
  INV_X1    g0186(.A(G190), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n386), .B2(G200), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n352), .A3(new_n361), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n389), .A2(new_n352), .A3(KEYINPUT17), .A4(new_n361), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n382), .A2(new_n385), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n217), .B1(new_n273), .B2(new_n276), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n228), .A2(G1698), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G226), .B2(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n401), .B2(new_n332), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n255), .B1(new_n265), .B2(new_n269), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n255), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n270), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT13), .B1(new_n406), .B2(new_n396), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n407), .A3(G190), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n292), .A2(new_n216), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT12), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n302), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n250), .B2(new_n300), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n290), .A2(new_n412), .A3(KEYINPUT11), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n292), .A2(new_n286), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(G68), .A3(new_n297), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT11), .B1(new_n290), .B2(new_n412), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G200), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n404), .B2(new_n407), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n398), .B1(new_n397), .B2(new_n403), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n406), .A2(new_n396), .A3(KEYINPUT13), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT14), .ZN(new_n427));
  INV_X1    g0227(.A(new_n423), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n404), .B2(new_n407), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n404), .A2(new_n407), .A3(G179), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n418), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n422), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n332), .A2(G107), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n436), .B(new_n437), .C1(new_n251), .C2(new_n217), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n255), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n271), .A2(new_n272), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n441));
  OAI21_X1  g0241(.A(G244), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n442), .A3(new_n270), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n443), .A2(new_n321), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n299), .A2(new_n303), .B1(new_n211), .B2(new_n250), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT15), .B(G87), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n300), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n286), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n250), .B1(new_n294), .B2(new_n296), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n414), .A2(new_n449), .B1(new_n250), .B2(new_n292), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT70), .B1(new_n444), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(new_n443), .B2(new_n321), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT70), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n443), .A2(G179), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n451), .B1(new_n443), .B2(G200), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n387), .B2(new_n443), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n325), .A2(new_n395), .A3(new_n435), .A4(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(G264), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n463));
  OAI211_X1 g0263(.A(G257), .B(new_n248), .C1(new_n330), .C2(new_n331), .ZN(new_n464));
  INV_X1    g0264(.A(G303), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n463), .B(new_n464), .C1(new_n465), .C2(new_n247), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n255), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n260), .A2(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT80), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n269), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n258), .A2(G1), .ZN(new_n475));
  INV_X1    g0275(.A(new_n471), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(new_n469), .ZN(new_n477));
  OAI21_X1  g0277(.A(G274), .B1(new_n254), .B2(new_n210), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT80), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n472), .A2(new_n255), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G270), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n467), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G200), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT78), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n244), .B2(G1), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n260), .A2(KEYINPUT78), .A3(G33), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n414), .A2(G116), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n309), .A2(G20), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n285), .A2(new_n210), .B1(G20), .B2(new_n490), .ZN(new_n493));
  AOI21_X1  g0293(.A(G20), .B1(G33), .B2(G283), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(G33), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n497), .A2(new_n498), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n492), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n479), .A2(new_n474), .B1(new_n481), .B2(G270), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(G190), .A3(new_n467), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n484), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT86), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n483), .A2(KEYINPUT21), .A3(G169), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n503), .A2(G179), .A3(new_n467), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n321), .B1(new_n503), .B2(new_n467), .ZN(new_n513));
  INV_X1    g0313(.A(new_n499), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n491), .B(new_n489), .C1(new_n514), .C2(new_n500), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT21), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n508), .A2(new_n509), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT85), .B1(new_n519), .B2(new_n502), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n507), .A2(new_n512), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n522));
  OAI211_X1 g0322(.A(G250), .B(new_n248), .C1(new_n330), .C2(new_n331), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n244), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n255), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n481), .A2(G264), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n480), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n525), .A2(new_n255), .B1(new_n481), .B2(G264), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT89), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n480), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n532), .A3(G169), .ZN(new_n533));
  INV_X1    g0333(.A(new_n528), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G179), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(G20), .B1(new_n245), .B2(new_n246), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT87), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT22), .A4(G87), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n244), .A2(new_n490), .A3(G20), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n211), .A2(G107), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT23), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT23), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n211), .B2(G107), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n540), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n211), .B(G87), .C1(new_n330), .C2(new_n331), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT87), .B(KEYINPUT22), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n539), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT24), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n539), .A2(new_n545), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n326), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g0353(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n554));
  NAND2_X1  g0354(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n309), .A2(new_n541), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n291), .A2(new_n211), .A3(G107), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n287), .A2(new_n488), .A3(new_n310), .A4(new_n289), .ZN(new_n558));
  INV_X1    g0358(.A(G107), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n556), .B1(new_n555), .B2(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n536), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(G190), .B1(new_n529), .B2(new_n532), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n534), .A2(G200), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n568));
  OAI211_X1 g0368(.A(G238), .B(new_n248), .C1(new_n330), .C2(new_n331), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n244), .C2(new_n490), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n255), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n468), .B(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n255), .A2(new_n219), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n574), .B1(new_n269), .B2(new_n475), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n575), .A3(G190), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT84), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n211), .A2(G33), .A3(G97), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT19), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT83), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(KEYINPUT83), .A3(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n211), .B1(new_n399), .B2(new_n579), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G97), .A2(G107), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n218), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n537), .A2(G68), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n326), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n558), .A2(new_n218), .ZN(new_n590));
  INV_X1    g0390(.A(new_n446), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(new_n310), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n571), .A2(new_n575), .A3(new_n594), .A4(G190), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n571), .A2(new_n575), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G200), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n577), .A2(new_n593), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n558), .A2(new_n446), .ZN(new_n599));
  INV_X1    g0399(.A(new_n592), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n584), .A2(new_n588), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n326), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n596), .A2(new_n321), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n571), .A2(new_n575), .A3(new_n371), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n558), .A2(G97), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n310), .A2(new_n495), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(KEYINPUT79), .A3(new_n609), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n336), .A2(new_n327), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G107), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT6), .ZN(new_n616));
  AND2_X1   g0416(.A1(G97), .A2(G107), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(new_n586), .ZN(new_n618));
  NAND2_X1  g0418(.A1(KEYINPUT6), .A2(G97), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT77), .B1(new_n619), .B2(G107), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT77), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(new_n559), .A3(KEYINPUT6), .A4(G97), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n618), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n623), .A2(G20), .B1(G77), .B2(new_n302), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n612), .A2(new_n613), .B1(new_n286), .B2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(G250), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n627));
  INV_X1    g0427(.A(G283), .ZN(new_n628));
  OAI211_X1 g0428(.A(G244), .B(new_n248), .C1(new_n330), .C2(new_n331), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT4), .ZN(new_n630));
  OAI221_X1 g0430(.A(new_n627), .B1(new_n244), .B2(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n255), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n479), .A2(new_n474), .B1(new_n481), .B2(G257), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G190), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n627), .B1(new_n244), .B2(new_n628), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n629), .A2(new_n630), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n274), .B1(new_n639), .B2(new_n632), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n481), .A2(G257), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n480), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT81), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT81), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n626), .B(new_n636), .C1(new_n646), .C2(new_n420), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n480), .A2(new_n641), .A3(new_n644), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n480), .B2(new_n641), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n371), .B(new_n634), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n625), .A2(new_n286), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT79), .B1(new_n608), .B2(new_n609), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n608), .A2(KEYINPUT79), .A3(new_n609), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n321), .B1(new_n640), .B2(new_n642), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n650), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n607), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n462), .A2(new_n521), .A3(new_n567), .A4(new_n657), .ZN(G372));
  INV_X1    g0458(.A(KEYINPUT91), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n457), .B1(new_n454), .B2(new_n455), .ZN(new_n660));
  AOI211_X1 g0460(.A(KEYINPUT70), .B(new_n452), .C1(new_n321), .C2(new_n443), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n453), .A2(KEYINPUT91), .A3(new_n456), .A4(new_n457), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n433), .B2(new_n434), .ZN(new_n664));
  INV_X1    g0464(.A(new_n422), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n392), .A3(new_n393), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n382), .B(new_n385), .C1(new_n664), .C2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT92), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n319), .B1(new_n667), .B2(KEYINPUT92), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n324), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n593), .A2(new_n597), .A3(new_n576), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n605), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n671), .B1(new_n656), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n606), .A2(new_n656), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n605), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n561), .B1(new_n533), .B2(new_n535), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT21), .B1(new_n513), .B2(new_n515), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n679), .A2(new_n510), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n605), .A2(new_n672), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n566), .A2(new_n647), .A3(new_n682), .A4(new_n656), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n670), .B1(new_n462), .B2(new_n685), .ZN(G369));
  XOR2_X1   g0486(.A(KEYINPUT94), .B(G330), .Z(new_n687));
  OAI21_X1  g0487(.A(new_n518), .B1(new_n510), .B2(new_n511), .ZN(new_n688));
  AOI211_X1 g0488(.A(KEYINPUT85), .B(new_n502), .C1(new_n508), .C2(new_n509), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR3_X1    g0490(.A1(new_n291), .A2(KEYINPUT27), .A3(G20), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT27), .B1(new_n291), .B2(G20), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G343), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT93), .Z(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n502), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n690), .A2(new_n507), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n680), .B2(new_n510), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n687), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n695), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n562), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n563), .A2(new_n702), .A3(new_n566), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n679), .A2(new_n701), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n690), .A2(new_n701), .ZN(new_n707));
  INV_X1    g0507(.A(new_n567), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n679), .A2(new_n695), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT95), .ZN(G399));
  INV_X1    g0513(.A(new_n207), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n587), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n214), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT96), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  INV_X1    g0522(.A(new_n596), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n530), .A3(new_n634), .A4(new_n635), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n721), .B(new_n722), .C1(new_n724), .C2(new_n509), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n634), .B1(new_n648), .B2(new_n649), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(G179), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n483), .A4(new_n528), .ZN(new_n728));
  INV_X1    g0528(.A(new_n509), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n640), .A2(new_n642), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n530), .A2(new_n571), .A3(new_n575), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n721), .A2(new_n722), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n729), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n725), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT97), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT97), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n734), .A2(new_n737), .A3(KEYINPUT31), .A4(new_n701), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(new_n701), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n736), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n657), .A2(new_n567), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n690), .A3(new_n507), .A4(new_n695), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n687), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n695), .B1(new_n678), .B2(new_n684), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT98), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND4_X1   g0548(.A1(new_n566), .A2(new_n647), .A3(new_n682), .A4(new_n656), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n563), .B(new_n518), .C1(new_n502), .C2(new_n519), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n605), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n650), .A2(new_n654), .A3(new_n655), .ZN(new_n753));
  INV_X1    g0553(.A(new_n676), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n607), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n755), .B2(new_n674), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n701), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n748), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT99), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n688), .A2(new_n679), .A3(new_n689), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n683), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n520), .A2(new_n563), .A3(new_n512), .A4(new_n518), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n749), .A2(new_n764), .A3(KEYINPUT99), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n753), .A2(KEYINPUT26), .A3(new_n682), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n676), .B1(new_n606), .B2(new_n656), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n752), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n763), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT29), .A3(new_n695), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n745), .B1(new_n760), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n720), .B1(new_n771), .B2(G1), .ZN(G364));
  INV_X1    g0572(.A(new_n700), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n308), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n260), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n715), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n698), .A2(new_n687), .A3(new_n699), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n773), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n698), .A2(new_n699), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n210), .B1(G20), .B2(new_n321), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n211), .A2(new_n371), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n387), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT104), .B(G326), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n211), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(new_n387), .A3(G200), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n790), .A2(new_n791), .B1(new_n793), .B2(new_n628), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n788), .A2(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(KEYINPUT33), .A2(G317), .ZN(new_n797));
  NAND2_X1  g0597(.A1(KEYINPUT33), .A2(G317), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n387), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n371), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n794), .B(new_n799), .C1(G294), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G190), .A2(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n247), .B1(new_n806), .B2(G329), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n465), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n787), .A2(KEYINPUT102), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n787), .A2(KEYINPUT102), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n800), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n809), .B1(new_n813), .B2(G322), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n804), .B1(new_n810), .B2(new_n811), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT103), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(KEYINPUT103), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n803), .B(new_n814), .C1(new_n815), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n808), .A2(new_n218), .ZN(new_n822));
  INV_X1    g0622(.A(new_n802), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n796), .A2(new_n216), .B1(new_n823), .B2(new_n495), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(G50), .C2(new_n789), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n819), .A2(G77), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n813), .A2(G58), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n247), .B1(new_n793), .B2(new_n559), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n806), .A2(KEYINPUT32), .A3(G159), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT32), .ZN(new_n830));
  INV_X1    g0630(.A(G159), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n805), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n828), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n786), .B1(new_n821), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n783), .A2(new_n785), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n247), .A2(new_n207), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT100), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G355), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(G116), .B2(new_n207), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT101), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n714), .A2(new_n247), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(G45), .B2(new_n214), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n241), .B2(G45), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n841), .B2(new_n842), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n837), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n835), .A2(new_n848), .A3(new_n778), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n784), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n780), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G396));
  AOI22_X1  g0652(.A1(new_n795), .A2(G150), .B1(new_n789), .B2(G137), .ZN(new_n853));
  INV_X1    g0653(.A(G143), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n854), .B2(new_n812), .C1(new_n820), .C2(new_n831), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT34), .Z(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n247), .B1(new_n805), .B2(new_n857), .C1(new_n216), .C2(new_n793), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n823), .A2(new_n339), .B1(new_n808), .B2(new_n305), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n247), .B1(new_n806), .B2(G311), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n861), .B1(new_n823), .B2(new_n495), .C1(new_n812), .C2(new_n524), .ZN(new_n862));
  INV_X1    g0662(.A(new_n808), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n795), .A2(G283), .B1(new_n863), .B2(G107), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n864), .B1(new_n218), .B2(new_n793), .C1(new_n465), .C2(new_n790), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n862), .B(new_n865), .C1(G116), .C2(new_n819), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n785), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n785), .A2(new_n781), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n867), .B(new_n777), .C1(G77), .C2(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT105), .Z(new_n871));
  NOR2_X1   g0671(.A1(new_n695), .A2(new_n452), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n662), .A2(new_n663), .A3(new_n872), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n460), .B1(new_n452), .B2(new_n695), .C1(new_n660), .C2(new_n661), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n871), .B1(new_n782), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n757), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n748), .A2(new_n758), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n875), .ZN(new_n879));
  INV_X1    g0679(.A(new_n745), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n777), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n880), .B2(new_n879), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n876), .A2(new_n882), .ZN(G384));
  NOR2_X1   g0683(.A1(new_n774), .A2(new_n260), .ZN(new_n884));
  INV_X1    g0684(.A(new_n431), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n432), .B1(new_n429), .B2(new_n430), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n434), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n701), .A2(new_n434), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n665), .A3(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n434), .B(new_n701), .C1(new_n433), .C2(new_n422), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n889), .A2(new_n890), .B1(new_n873), .B2(new_n874), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NOR4_X1   g0692(.A1(new_n521), .A2(new_n657), .A3(new_n567), .A4(new_n701), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n741), .A2(new_n735), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n362), .A2(new_n693), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n381), .A2(new_n896), .A3(new_n897), .A4(new_n390), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT106), .ZN(new_n899));
  INV_X1    g0699(.A(new_n343), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n338), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n344), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n338), .A2(new_n345), .B1(new_n287), .B2(new_n289), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n360), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n693), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n338), .A2(new_n345), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n290), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT16), .B1(new_n338), .B2(new_n900), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n361), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(KEYINPUT106), .A3(new_n693), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n380), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n906), .A2(new_n911), .A3(new_n390), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n906), .A2(new_n911), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n898), .A2(new_n914), .B1(new_n394), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n898), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n394), .A2(new_n915), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n895), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n896), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n381), .A2(new_n896), .A3(new_n390), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n394), .A2(new_n923), .B1(new_n925), .B2(new_n898), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT108), .B1(new_n926), .B2(KEYINPUT38), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n394), .A2(new_n923), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n898), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT108), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n927), .A2(new_n933), .A3(new_n917), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n889), .A2(new_n890), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n875), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n741), .A2(new_n735), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n744), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n922), .B1(new_n939), .B2(KEYINPUT40), .ZN(new_n940));
  INV_X1    g0740(.A(new_n462), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n937), .A2(new_n744), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n940), .B(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n687), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n918), .A2(KEYINPUT38), .A3(new_n919), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT39), .B1(new_n947), .B2(new_n920), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT107), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT39), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n927), .A2(new_n933), .A3(new_n950), .A4(new_n917), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT107), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(KEYINPUT39), .C1(new_n947), .C2(new_n920), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n433), .A2(new_n434), .A3(new_n695), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n921), .A2(new_n917), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n458), .A2(new_n701), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n757), .B2(new_n875), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n961), .A3(new_n935), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n382), .A2(new_n385), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n905), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n957), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n760), .A2(new_n770), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n670), .B1(new_n967), .B2(new_n462), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n966), .B(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n884), .B1(new_n946), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n969), .B2(new_n946), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n623), .A2(KEYINPUT35), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n623), .A2(KEYINPUT35), .ZN(new_n973));
  NOR4_X1   g0773(.A1(new_n972), .A2(new_n973), .A3(new_n490), .A4(new_n213), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT36), .Z(new_n975));
  OR3_X1    g0775(.A1(new_n214), .A2(new_n250), .A3(new_n340), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n305), .A2(G68), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(G1), .A3(new_n308), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n971), .A2(new_n975), .A3(new_n979), .ZN(G367));
  XOR2_X1   g0780(.A(new_n715), .B(KEYINPUT41), .Z(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n647), .B(new_n656), .C1(new_n626), .C2(new_n695), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n753), .A2(new_n701), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n711), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n985), .B1(new_n709), .B2(new_n710), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n706), .ZN(new_n992));
  INV_X1    g0792(.A(new_n706), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n988), .A2(new_n993), .A3(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT114), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n709), .B1(new_n707), .B2(new_n705), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT113), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n773), .A3(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n707), .A2(new_n705), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n1000), .B(new_n709), .C1(new_n700), .C2(KEYINPUT113), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n771), .A2(new_n996), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n996), .B1(new_n771), .B2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT115), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n967), .A2(new_n1002), .A3(new_n880), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT114), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT115), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n771), .A2(new_n996), .A3(new_n1002), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n995), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n771), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n982), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n775), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n707), .A2(new_n985), .A3(new_n708), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT42), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n679), .A2(new_n647), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n701), .B1(new_n1017), .B2(new_n656), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1015), .B2(KEYINPUT42), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n695), .A2(new_n593), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(new_n605), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n682), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1016), .A2(new_n1019), .B1(KEYINPUT43), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT110), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n706), .A2(new_n985), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1031), .A2(KEYINPUT112), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT112), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1033), .A2(new_n1035), .B1(KEYINPUT111), .B2(new_n1029), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1033), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1034), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1014), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(G137), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n808), .A2(new_n339), .B1(new_n805), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n823), .A2(new_n216), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G159), .B2(new_n795), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n854), .B2(new_n790), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1044), .B(new_n1047), .C1(G150), .C2(new_n813), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n247), .B1(new_n793), .B2(new_n250), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT116), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(new_n305), .C2(new_n820), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n820), .A2(new_n628), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n790), .A2(new_n815), .B1(new_n823), .B2(new_n559), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G294), .B2(new_n795), .ZN(new_n1054));
  INV_X1    g0854(.A(G317), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n332), .B1(new_n805), .B2(new_n1055), .C1(new_n495), .C2(new_n793), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n813), .B2(G303), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n863), .A2(G116), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT46), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1051), .B1(new_n1052), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT47), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n785), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n837), .B1(new_n714), .B2(new_n591), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n234), .A2(new_n844), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n778), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n783), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1063), .B(new_n1066), .C1(new_n1067), .C2(new_n1023), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1042), .A2(new_n1068), .ZN(G387));
  NAND2_X1  g0869(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n715), .C1(new_n771), .C2(new_n1002), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n839), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1072), .A2(new_n717), .B1(G107), .B2(new_n207), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n231), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n299), .A2(G50), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n717), .B(new_n258), .C1(new_n216), .C2(new_n250), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n844), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1074), .A2(G45), .B1(KEYINPUT118), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1079), .A2(KEYINPUT118), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1073), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n777), .B1(new_n1082), .B2(new_n837), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n332), .B1(new_n806), .B2(G150), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n495), .B2(new_n793), .C1(new_n812), .C2(new_n305), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n823), .A2(new_n446), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G77), .B2(new_n863), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n831), .B2(new_n790), .C1(new_n299), .C2(new_n796), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1085), .B(new_n1088), .C1(G68), .C2(new_n819), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT119), .Z(new_n1090));
  OAI22_X1  g0890(.A1(new_n823), .A2(new_n628), .B1(new_n808), .B2(new_n524), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n795), .A2(G311), .B1(new_n789), .B2(G322), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n1055), .B2(new_n812), .C1(new_n820), .C2(new_n465), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT48), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT49), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n332), .B1(new_n805), .B2(new_n791), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n793), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(G116), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1090), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1083), .B1(new_n1103), .B2(new_n785), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n703), .A2(new_n704), .A3(new_n783), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1002), .A2(new_n776), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1071), .A2(new_n1106), .ZN(G393));
  AOI21_X1  g0907(.A(new_n716), .B1(new_n995), .B2(new_n1070), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n995), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n995), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n986), .A2(new_n783), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n836), .B1(new_n495), .B2(new_n207), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n238), .B2(new_n844), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n247), .B1(new_n806), .B2(G322), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n559), .B2(new_n793), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n796), .A2(new_n465), .B1(new_n823), .B2(new_n490), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(G283), .C2(new_n863), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n812), .A2(new_n815), .B1(new_n790), .B2(new_n1055), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT52), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(new_n524), .C2(new_n820), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n247), .B1(new_n805), .B2(new_n854), .C1(new_n218), .C2(new_n793), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n796), .A2(new_n305), .B1(new_n823), .B2(new_n250), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(G68), .C2(new_n863), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n299), .B2(new_n820), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n813), .A2(G159), .B1(G150), .B2(new_n789), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT51), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1121), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n778), .B(new_n1114), .C1(new_n1128), .C2(new_n785), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1111), .A2(new_n776), .B1(new_n1112), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1110), .A2(new_n1130), .ZN(G390));
  INV_X1    g0931(.A(new_n935), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n955), .B1(new_n960), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n949), .A2(new_n951), .A3(new_n953), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n769), .A2(new_n695), .A3(new_n875), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n959), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n935), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n955), .A3(new_n934), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G330), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n937), .B2(new_n744), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(new_n936), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n745), .A2(new_n875), .A3(new_n935), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1134), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1143), .A2(new_n462), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n670), .C1(new_n462), .C2(new_n967), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n935), .B1(new_n745), .B2(new_n875), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n961), .B1(new_n1154), .B2(new_n1144), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n935), .B1(new_n1142), .B2(new_n875), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(new_n1137), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1146), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT120), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n716), .B1(new_n1149), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1148), .A2(new_n1161), .A3(new_n1160), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1149), .A2(new_n776), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n777), .B1(new_n353), .B2(new_n869), .ZN(new_n1167));
  INV_X1    g0967(.A(G125), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n247), .B1(new_n805), .B2(new_n1168), .C1(new_n796), .C2(new_n1043), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n813), .B2(G132), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n823), .A2(new_n831), .B1(new_n793), .B2(new_n305), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G128), .B2(new_n789), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n808), .A2(new_n301), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT53), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n820), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n820), .A2(new_n495), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n247), .B(new_n822), .C1(G294), .C2(new_n806), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n813), .A2(G116), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G68), .A2(new_n1100), .B1(new_n802), .B2(G77), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n795), .A2(G107), .B1(new_n789), .B2(G283), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1175), .A2(new_n1177), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1167), .B1(new_n1184), .B2(new_n785), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n954), .B2(new_n782), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1165), .A2(new_n1166), .A3(new_n1186), .ZN(G378));
  AOI21_X1  g0987(.A(KEYINPUT121), .B1(new_n318), .B2(new_n323), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n311), .A2(new_n693), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT55), .Z(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n318), .A2(KEYINPUT121), .A3(new_n323), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1189), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n318), .A2(KEYINPUT121), .A3(new_n323), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1191), .B1(new_n1195), .B2(new_n1188), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1197), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n940), .A2(new_n1141), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1200), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1198), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n958), .A2(new_n892), .A3(new_n938), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n942), .A2(new_n891), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT38), .B1(new_n928), .B2(new_n929), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1207), .A2(new_n931), .B1(new_n916), .B2(KEYINPUT38), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1206), .B1(new_n1208), .B2(new_n927), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1205), .B1(new_n1209), .B2(new_n892), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1204), .B1(new_n1210), .B2(G330), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n966), .B1(new_n1202), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1201), .B1(new_n940), .B2(new_n1141), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(G330), .A3(new_n1204), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n957), .A4(new_n965), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1145), .A2(new_n1147), .A3(new_n1159), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1153), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT57), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT123), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1215), .A2(new_n1212), .B1(new_n1217), .B2(new_n1153), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT123), .B1(new_n1222), .B2(KEYINPUT57), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n716), .B1(new_n1222), .B2(KEYINPUT57), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1216), .A2(new_n776), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n869), .A2(G50), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n257), .B(new_n332), .C1(new_n805), .C2(new_n628), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1228), .B(new_n1045), .C1(G107), .C2(new_n813), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n796), .A2(new_n495), .B1(new_n250), .B2(new_n808), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n790), .A2(new_n490), .B1(new_n793), .B2(new_n339), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1229), .B(new_n1232), .C1(new_n820), .C2(new_n446), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT58), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n332), .A2(new_n257), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G50), .B1(new_n244), .B2(new_n257), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1233), .A2(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n790), .A2(new_n1168), .B1(new_n808), .B2(new_n1176), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n796), .A2(new_n857), .B1(new_n823), .B2(new_n301), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(G128), .C2(new_n813), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1043), .B2(new_n820), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1100), .A2(G159), .ZN(new_n1243));
  AOI211_X1 g1043(.A(G33), .B(G41), .C1(new_n806), .C2(G124), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1237), .B1(new_n1234), .B2(new_n1233), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n778), .B(new_n1227), .C1(new_n1247), .C2(new_n785), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1204), .B2(new_n782), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1226), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1225), .A2(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n1132), .A2(new_n781), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n819), .A2(G150), .B1(G50), .B2(new_n802), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT124), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n789), .A2(G132), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1256), .B1(new_n831), .B2(new_n808), .C1(new_n796), .C2(new_n1176), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n332), .B1(new_n806), .B2(G128), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1258), .B1(new_n339), .B2(new_n793), .C1(new_n812), .C2(new_n1043), .ZN(new_n1259));
  OR3_X1    g1059(.A1(new_n1255), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n796), .A2(new_n490), .B1(new_n495), .B2(new_n808), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1086), .B(new_n1261), .C1(G294), .C2(new_n789), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n332), .B1(new_n805), .B2(new_n465), .C1(new_n250), .C2(new_n793), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n813), .B2(G283), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1262), .B(new_n1264), .C1(new_n559), .C2(new_n820), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n786), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n778), .B(new_n1266), .C1(new_n216), .C2(new_n868), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1159), .A2(new_n776), .B1(new_n1253), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n981), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1152), .A2(new_n1155), .A3(new_n1158), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(G381));
  NOR2_X1   g1073(.A1(G375), .A2(G378), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1040), .B1(new_n1013), .B2(new_n775), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1068), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1275), .A2(G390), .A3(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1071), .A2(new_n851), .A3(new_n1106), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(G381), .A2(G384), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1274), .A2(new_n1277), .A3(new_n1279), .ZN(G407));
  INV_X1    g1080(.A(G343), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(G213), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1274), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(G407), .A2(G213), .A3(new_n1284), .ZN(G409));
  INV_X1    g1085(.A(G2897), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G384), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n1155), .A4(new_n1158), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n715), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1160), .A2(KEYINPUT60), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n1271), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1293), .B2(new_n1269), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1271), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(KEYINPUT60), .B2(new_n1160), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G384), .B(new_n1268), .C1(new_n1296), .C2(new_n1291), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT125), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1288), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  AOI211_X1 g1100(.A(KEYINPUT125), .B(new_n1287), .C1(new_n1294), .C2(new_n1297), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n1300), .A2(new_n1301), .B1(new_n1299), .B2(new_n1298), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1216), .A2(new_n1218), .A3(KEYINPUT57), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n715), .B(new_n1304), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1222), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G378), .B(new_n1251), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1166), .A2(new_n1186), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1222), .A2(new_n982), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n1250), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1307), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1282), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT61), .B1(new_n1303), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1313), .B2(new_n1298), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1278), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n851), .B1(new_n1071), .B2(new_n1106), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AND2_X1   g1119(.A1(new_n1110), .A2(new_n1130), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1320), .B1(new_n1042), .B2(new_n1068), .ZN(new_n1321));
  OAI211_X1 g1121(.A(KEYINPUT126), .B(new_n1319), .C1(new_n1321), .C2(new_n1277), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1042), .A2(new_n1068), .A3(new_n1320), .ZN(new_n1323));
  OR2_X1    g1123(.A1(new_n1319), .A2(KEYINPUT126), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1319), .A2(KEYINPUT126), .ZN(new_n1325));
  OAI21_X1  g1125(.A(G390), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1322), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1283), .B1(new_n1307), .B2(new_n1311), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1298), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1314), .A2(new_n1316), .A3(new_n1329), .A4(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1330), .A2(new_n1334), .A3(new_n1331), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT61), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1330), .B2(new_n1302), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1334), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1335), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1333), .B1(new_n1339), .B2(new_n1329), .ZN(G405));
  INV_X1    g1140(.A(new_n1307), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G378), .B1(new_n1225), .B2(new_n1251), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1331), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(G375), .A2(new_n1309), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1344), .A2(new_n1298), .A3(new_n1307), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1343), .A2(new_n1328), .A3(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1328), .B1(new_n1343), .B2(new_n1345), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT127), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1346), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  AOI211_X1 g1149(.A(KEYINPUT127), .B(new_n1328), .C1(new_n1343), .C2(new_n1345), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(G402));
endmodule


