//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n205), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n217), .A2(new_n218), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n212), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT65), .Z(new_n225));
  INV_X1    g0025(.A(KEYINPUT1), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n212), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n210), .ZN(new_n233));
  INV_X1    g0033(.A(new_n201), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n231), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  AND3_X1   g0037(.A1(new_n227), .A2(new_n228), .A3(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  INV_X1    g0044(.A(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT2), .B(G226), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n252), .B(new_n255), .Z(G351));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G58), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT8), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n258), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n232), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n266), .A2(new_n268), .B1(new_n202), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT71), .B1(new_n210), .B2(G1), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT71), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(new_n209), .A3(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  XOR2_X1   g0076(.A(new_n276), .B(KEYINPUT72), .Z(new_n277));
  INV_X1    g0077(.A(KEYINPUT70), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n270), .B2(new_n268), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n269), .A2(KEYINPUT70), .A3(new_n232), .A4(new_n267), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n271), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT9), .ZN(new_n283));
  INV_X1    g0083(.A(G200), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G222), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n288), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n295), .A2(G223), .B1(G77), .B2(new_n294), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n286), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  AOI21_X1  g0099(.A(G1), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(new_n286), .A3(G274), .ZN(new_n301));
  INV_X1    g0101(.A(G226), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n286), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n301), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n283), .B1(new_n284), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n306), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT75), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OR3_X1    g0110(.A1(new_n307), .A2(KEYINPUT10), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT10), .B1(new_n307), .B2(new_n310), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G68), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n270), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT12), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n270), .A2(new_n268), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(G68), .A3(new_n275), .ZN(new_n318));
  INV_X1    g0118(.A(G77), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n265), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n257), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n321), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n268), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT11), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n316), .B(new_n318), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n245), .A2(G1698), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(G226), .B2(G1698), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n331), .B2(new_n294), .ZN(new_n332));
  INV_X1    g0132(.A(new_n286), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n286), .A2(G238), .A3(new_n303), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT76), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n301), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n301), .B2(new_n335), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT13), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n334), .B(new_n341), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(G169), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(G179), .A3(new_n342), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n344), .B1(new_n343), .B2(G169), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n328), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n327), .B1(new_n343), .B2(new_n309), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n284), .B1(new_n340), .B2(new_n342), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G169), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n308), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n306), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n282), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G244), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n301), .B1(new_n360), .B2(new_n304), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n287), .A2(G238), .A3(G1698), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n363), .C1(new_n206), .C2(new_n287), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n361), .B1(new_n364), .B2(new_n333), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n284), .ZN(new_n366));
  AOI211_X1 g0166(.A(new_n309), .B(new_n361), .C1(new_n364), .C2(new_n333), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n275), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n319), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n317), .B1(new_n319), .B2(new_n270), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT8), .B(G58), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n372), .A2(new_n321), .B1(new_n210), .B2(new_n319), .ZN(new_n373));
  XOR2_X1   g0173(.A(KEYINPUT15), .B(G87), .Z(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(KEYINPUT73), .B1(new_n264), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n376), .B1(new_n210), .B2(new_n319), .C1(new_n372), .C2(new_n321), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT74), .B1(new_n378), .B2(new_n268), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  INV_X1    g0180(.A(new_n268), .ZN(new_n381));
  AOI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n375), .C2(new_n377), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n368), .B(new_n371), .C1(new_n379), .C2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n365), .A2(G169), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n357), .B2(new_n365), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n371), .B1(new_n379), .B2(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n313), .A2(new_n354), .A3(new_n359), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT77), .B1(new_n263), .B2(KEYINPUT3), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(new_n292), .A3(G33), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n390), .A2(new_n392), .A3(new_n291), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT7), .B1(new_n393), .B2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n392), .A3(new_n291), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n210), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(G68), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n201), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT78), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n257), .A2(G159), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT78), .B(G20), .C1(new_n400), .C2(new_n201), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n396), .B1(new_n287), .B2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n294), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n314), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n409), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(new_n413), .A3(new_n268), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n262), .A2(new_n269), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n369), .B1(new_n279), .B2(new_n280), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(new_n262), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT79), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT79), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n415), .C1(new_n416), .C2(new_n262), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n302), .A2(G1698), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G223), .B2(G1698), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n395), .A2(new_n423), .B1(new_n263), .B2(new_n214), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n333), .ZN(new_n425));
  INV_X1    g0225(.A(new_n304), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n286), .A2(G274), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n426), .A2(G232), .B1(new_n427), .B2(new_n300), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n425), .A2(G190), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n284), .B1(new_n425), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n414), .A2(new_n421), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(KEYINPUT80), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT80), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n414), .A2(new_n421), .A3(new_n431), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n438), .B2(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n414), .A2(new_n421), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n425), .A2(new_n428), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n357), .B2(new_n441), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT18), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n389), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT84), .ZN(new_n450));
  AND2_X1   g0250(.A1(KEYINPUT4), .A2(G244), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n291), .A2(new_n293), .A3(new_n451), .A4(new_n288), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n291), .A2(new_n293), .A3(G250), .A4(G1698), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n360), .A2(G1698), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n390), .A2(new_n392), .A3(new_n291), .A4(new_n456), .ZN(new_n457));
  XOR2_X1   g0257(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n286), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n298), .A2(KEYINPUT5), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n209), .B(G45), .C1(new_n298), .C2(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(KEYINPUT83), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n299), .A2(G1), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G41), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n464), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G257), .B(new_n286), .C1(new_n463), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n462), .A2(KEYINPUT83), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n464), .A3(new_n467), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n427), .A2(new_n470), .A3(new_n461), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n450), .B1(new_n460), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n457), .A2(new_n458), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n333), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n477), .A2(KEYINPUT84), .A3(new_n472), .A4(new_n469), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n355), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n460), .A2(new_n473), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n205), .A2(KEYINPUT81), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT81), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G97), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G97), .A2(G107), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT6), .B1(new_n207), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(G20), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n319), .B2(new_n321), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n206), .B1(new_n410), .B2(new_n411), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n268), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n269), .A2(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n209), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n269), .A2(new_n494), .A3(new_n232), .A4(new_n267), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n496), .B2(G97), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n357), .A2(new_n481), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n473), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n284), .B1(new_n499), .B2(new_n477), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n492), .A2(new_n497), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n474), .A2(new_n478), .A3(G190), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n480), .A2(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n393), .A2(KEYINPUT88), .A3(new_n210), .A4(G87), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT88), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n390), .A2(new_n392), .A3(new_n210), .A4(new_n291), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n214), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(KEYINPUT22), .A3(new_n509), .ZN(new_n510));
  OR4_X1    g0310(.A1(KEYINPUT22), .A2(new_n294), .A3(G20), .A4(new_n214), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT23), .B1(new_n206), .B2(G20), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n513), .A2(new_n514), .B1(G20), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n505), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(KEYINPUT24), .B(new_n516), .C1(new_n510), .C2(new_n511), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n268), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT25), .B1(new_n270), .B2(new_n206), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n523), .B1(G107), .B2(new_n496), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n216), .A2(G1698), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(G250), .B2(G1698), .ZN(new_n526));
  INV_X1    g0326(.A(G294), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n395), .A2(new_n526), .B1(new_n263), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n333), .ZN(new_n529));
  OAI211_X1 g0329(.A(G264), .B(new_n286), .C1(new_n463), .C2(new_n468), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n472), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n309), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(G200), .B2(new_n531), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n520), .A2(new_n524), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n374), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n270), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n496), .A2(G87), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  XNOR2_X1  g0338(.A(KEYINPUT81), .B(G97), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(new_n265), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n210), .B1(new_n329), .B2(new_n538), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n483), .A2(new_n485), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n214), .A2(new_n206), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  OR3_X1    g0345(.A1(new_n508), .A2(KEYINPUT85), .A3(new_n314), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT85), .B1(new_n508), .B2(new_n314), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n536), .B(new_n537), .C1(new_n548), .C2(new_n381), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n215), .B1(new_n299), .B2(G1), .ZN(new_n551));
  INV_X1    g0351(.A(G274), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n209), .A2(new_n552), .A3(G45), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n286), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n360), .A2(G1698), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G238), .B2(G1698), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n515), .B1(new_n395), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n555), .B1(new_n558), .B2(new_n333), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(new_n284), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(G190), .B2(new_n559), .ZN(new_n561));
  OAI221_X1 g0361(.A(new_n536), .B1(new_n535), .B2(new_n495), .C1(new_n548), .C2(new_n381), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n559), .A2(G169), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n357), .B2(new_n559), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n550), .A2(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n504), .A2(new_n534), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n454), .A2(new_n210), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n542), .B2(new_n263), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT20), .ZN(new_n570));
  INV_X1    g0370(.A(G116), .ZN(new_n571));
  AOI22_X1  g0371(.A1(KEYINPUT86), .A2(new_n570), .B1(new_n571), .B2(G20), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n268), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n567), .B(KEYINPUT20), .C1(new_n569), .C2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n210), .B(new_n454), .C1(new_n539), .C2(G33), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n567), .A2(KEYINPUT20), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n575), .A2(new_n268), .A3(new_n572), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n269), .A2(new_n571), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n496), .B2(new_n571), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n574), .A2(new_n577), .A3(new_n579), .A4(KEYINPUT87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n463), .A2(new_n468), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n292), .A2(G33), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n587));
  OAI21_X1  g0387(.A(G303), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n216), .A2(new_n288), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G264), .B2(new_n288), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n395), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n427), .A2(new_n585), .B1(new_n591), .B2(new_n333), .ZN(new_n592));
  OAI211_X1 g0392(.A(G270), .B(new_n286), .C1(new_n463), .C2(new_n468), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n355), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n584), .A2(KEYINPUT21), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n333), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(G179), .A3(new_n593), .A4(new_n472), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n584), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT21), .B1(new_n584), .B2(new_n594), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n531), .A2(new_n355), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G179), .B2(new_n531), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n512), .A2(new_n517), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT24), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n512), .A2(new_n505), .A3(new_n517), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n381), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n524), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n596), .A2(new_n472), .A3(new_n593), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n584), .B1(G200), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n309), .B2(new_n612), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n602), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n449), .A2(new_n566), .A3(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n359), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n349), .B1(new_n352), .B2(new_n387), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n439), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT90), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n440), .A2(new_n443), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n620), .B1(new_n440), .B2(new_n443), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n445), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n623), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(KEYINPUT18), .A3(new_n621), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n617), .B1(new_n628), .B2(new_n313), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n504), .A2(new_n534), .A3(new_n565), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT89), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n602), .A2(new_n611), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n584), .A2(new_n594), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n599), .A3(new_n595), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n604), .B1(new_n520), .B2(new_n524), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT89), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n630), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n550), .A2(new_n561), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n562), .A2(new_n564), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n480), .A2(new_n498), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n565), .A2(KEYINPUT26), .A3(new_n480), .A4(new_n498), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n645), .A2(new_n646), .B1(new_n562), .B2(new_n564), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n639), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n629), .B1(new_n449), .B2(new_n649), .ZN(G369));
  NAND3_X1  g0450(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n584), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n602), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(G330), .A3(new_n614), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n609), .B2(new_n610), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n534), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n611), .ZN(new_n662));
  INV_X1    g0462(.A(new_n656), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n637), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n637), .B1(new_n660), .B2(new_n534), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n636), .A2(new_n663), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(G399));
  NOR3_X1   g0472(.A1(new_n542), .A2(G116), .A3(new_n543), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT91), .ZN(new_n674));
  INV_X1    g0474(.A(new_n229), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n235), .B2(new_n677), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT94), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT93), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT92), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n592), .A2(new_n683), .A3(G179), .A4(new_n593), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n597), .A2(KEYINPUT92), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n559), .A2(new_n530), .A3(new_n529), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n479), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT30), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n474), .A2(new_n478), .A3(KEYINPUT30), .ZN(new_n691));
  INV_X1    g0491(.A(new_n559), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n612), .A2(new_n692), .A3(new_n357), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n531), .B1(new_n460), .B2(new_n473), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n690), .A2(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n656), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n694), .A2(new_n693), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n474), .A2(new_n478), .A3(KEYINPUT30), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n699), .B1(new_n687), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n690), .B2(new_n479), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n682), .B1(new_n698), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT31), .B1(new_n704), .B2(new_n656), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT93), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n681), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AOI211_X1 g0509(.A(new_n697), .B(new_n663), .C1(new_n701), .C2(new_n703), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT93), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n698), .A2(new_n682), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(KEYINPUT94), .A3(new_n712), .ZN(new_n713));
  OR3_X1    g0513(.A1(new_n615), .A2(new_n566), .A3(new_n656), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT95), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(KEYINPUT95), .A3(G330), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n636), .A2(new_n637), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n647), .B1(new_n566), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .A3(new_n663), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n656), .B1(new_n639), .B2(new_n647), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(KEYINPUT29), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n718), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n680), .B1(new_n726), .B2(G1), .ZN(G364));
  INV_X1    g0527(.A(G13), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n209), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n676), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n659), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n658), .A2(new_n614), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(G330), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n229), .A2(G355), .A3(new_n287), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G116), .B2(new_n229), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n393), .B(new_n675), .C1(new_n299), .C2(new_n236), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n252), .A2(new_n299), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n232), .B1(G20), .B2(new_n355), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n732), .B1(new_n742), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n210), .A2(G179), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G190), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G159), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n753), .A2(KEYINPUT32), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT32), .ZN(new_n756));
  INV_X1    g0556(.A(new_n753), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(G159), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n751), .A2(new_n309), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n755), .B(new_n758), .C1(G107), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n210), .A2(new_n357), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G190), .A3(new_n284), .ZN(new_n763));
  INV_X1    g0563(.A(G58), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n287), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n751), .A2(G190), .A3(G200), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n766), .A2(new_n202), .B1(new_n767), .B2(new_n214), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n762), .A2(new_n309), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n765), .B(new_n768), .C1(G68), .C2(new_n770), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n762), .A2(KEYINPUT96), .A3(new_n752), .ZN(new_n772));
  AOI21_X1  g0572(.A(KEYINPUT96), .B1(new_n762), .B2(new_n752), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G77), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n309), .A2(G200), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n210), .B1(new_n777), .B2(new_n357), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT97), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G97), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n761), .A2(new_n771), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  INV_X1    g0582(.A(new_n763), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n770), .A2(new_n782), .B1(new_n783), .B2(G322), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT98), .ZN(new_n785));
  INV_X1    g0585(.A(G303), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n767), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G283), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n778), .A2(new_n527), .B1(new_n759), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n766), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n787), .B(new_n789), .C1(G326), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n762), .A2(new_n752), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n287), .B(new_n794), .C1(G329), .C2(new_n757), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n781), .B1(new_n785), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n750), .B1(new_n797), .B2(new_n747), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n736), .B2(new_n746), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n737), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  AND3_X1   g0601(.A1(new_n715), .A2(KEYINPUT95), .A3(G330), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT95), .B1(new_n715), .B2(G330), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n386), .A2(new_n656), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n383), .A2(new_n387), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT100), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT100), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n383), .A2(new_n387), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n723), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n385), .A2(new_n386), .A3(new_n656), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n807), .A2(new_n813), .A3(new_n809), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n723), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n733), .B1(new_n804), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT101), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n816), .A2(KEYINPUT101), .B1(new_n804), .B2(new_n815), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n814), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n743), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n747), .A2(new_n743), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n732), .B1(G77), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n775), .A2(G116), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n769), .A2(new_n788), .B1(new_n767), .B2(new_n206), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n766), .A2(new_n786), .B1(new_n759), .B2(new_n214), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n294), .B1(new_n753), .B2(new_n793), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G294), .B2(new_n783), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n780), .A2(new_n825), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n783), .A2(G143), .B1(new_n790), .B2(G137), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n832), .B1(new_n833), .B2(new_n769), .C1(new_n774), .C2(new_n754), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n395), .B1(new_n757), .B2(G132), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n778), .A2(new_n764), .B1(new_n767), .B2(new_n202), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n759), .A2(new_n314), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n837), .B(new_n840), .C1(new_n834), .C2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n831), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT99), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n748), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n824), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n821), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n819), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n729), .A2(new_n209), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n347), .A2(new_n348), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n328), .B(new_n656), .C1(new_n853), .C2(new_n352), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n328), .A2(new_n656), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n349), .A2(new_n353), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n615), .A2(new_n566), .A3(new_n656), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n698), .A2(new_n705), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n814), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  INV_X1    g0661(.A(new_n654), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n440), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n627), .B2(new_n439), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n444), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n438), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n432), .B(new_n863), .C1(new_n622), .C2(new_n623), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n861), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n435), .A2(new_n437), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n408), .A2(new_n268), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n398), .B2(new_n407), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n421), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT102), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT102), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n421), .B(new_n876), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n862), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n443), .A3(new_n877), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n871), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  INV_X1    g0681(.A(new_n867), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n878), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n447), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n852), .B(new_n860), .C1(new_n870), .C2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT104), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n867), .B1(new_n880), .B2(KEYINPUT37), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n878), .B1(new_n439), .B2(new_n446), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n861), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n860), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n888), .B1(new_n892), .B2(KEYINPUT40), .ZN(new_n893));
  INV_X1    g0693(.A(new_n856), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n855), .B1(new_n349), .B2(new_n353), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n814), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n859), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n714), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n883), .B2(new_n885), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n889), .A2(new_n890), .A3(new_n861), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n852), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n887), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n714), .A2(new_n897), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n448), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(G330), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n448), .B2(new_n904), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT105), .Z(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n624), .A2(new_n626), .A3(new_n654), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n656), .B(new_n810), .C1(new_n639), .C2(new_n647), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n387), .A2(new_n656), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n857), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n886), .A2(new_n891), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n911), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT103), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n870), .A2(new_n886), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n853), .A2(new_n328), .A3(new_n663), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n891), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT103), .B(new_n911), .C1(new_n914), .C2(new_n916), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n919), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n629), .B1(new_n449), .B2(new_n724), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n928), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n851), .B1(new_n910), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n910), .B2(new_n930), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n486), .A2(new_n488), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(KEYINPUT35), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(KEYINPUT35), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n934), .A2(G116), .A3(new_n233), .A4(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n236), .A2(G77), .A3(new_n399), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(G50), .B2(new_n314), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(G1), .A3(new_n728), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n932), .A2(new_n937), .A3(new_n940), .ZN(G367));
  NOR2_X1   g0741(.A1(new_n675), .A2(new_n393), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n242), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n749), .B1(new_n675), .B2(new_n374), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n733), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT108), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n549), .A2(new_n656), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n565), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n642), .A2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(G317), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n395), .B1(new_n753), .B2(new_n951), .C1(new_n763), .C2(new_n786), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n775), .B2(G283), .ZN(new_n953));
  INV_X1    g0753(.A(new_n767), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(G116), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT46), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n778), .A2(new_n206), .B1(new_n769), .B2(new_n527), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n766), .A2(new_n793), .B1(new_n759), .B2(new_n539), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n953), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT109), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n779), .A2(G68), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n759), .A2(new_n319), .ZN(new_n963));
  INV_X1    g0763(.A(G143), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n964), .A2(new_n766), .B1(new_n769), .B2(new_n754), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(G58), .C2(new_n954), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n775), .A2(G50), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT110), .B(G137), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n287), .B1(new_n753), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G150), .B2(new_n783), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n966), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n961), .B1(new_n962), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(KEYINPUT47), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n747), .B1(new_n972), .B2(KEYINPUT47), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n946), .B1(new_n950), .B2(new_n746), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n501), .A2(new_n656), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n504), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n644), .A2(new_n663), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n670), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n979), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n671), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n670), .B2(new_n979), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(KEYINPUT106), .A3(new_n666), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n982), .A2(new_n990), .A3(new_n987), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT107), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n665), .B2(new_n669), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n659), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n994), .A2(new_n659), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n996), .A2(new_n997), .B1(new_n665), .B2(new_n669), .ZN(new_n998));
  INV_X1    g0798(.A(new_n997), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n665), .A2(new_n669), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n995), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n726), .B1(new_n992), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n676), .B(KEYINPUT41), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n731), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n950), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1000), .A2(new_n983), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT42), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n502), .A2(new_n503), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n637), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n656), .B1(new_n1014), .B2(new_n644), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1011), .B2(KEYINPUT42), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1007), .B(new_n1010), .C1(new_n1012), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n667), .A2(new_n979), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1012), .A2(new_n1016), .A3(new_n1009), .A4(new_n1008), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1020), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1022), .A2(new_n1017), .B1(new_n667), .B2(new_n979), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n975), .B1(new_n1006), .B2(new_n1024), .ZN(G387));
  NOR3_X1   g0825(.A1(new_n674), .A2(new_n675), .A3(new_n294), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n206), .B2(new_n675), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT111), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n674), .B(new_n299), .C1(new_n314), .C2(new_n319), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT112), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n372), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n942), .B1(new_n299), .B2(new_n248), .C1(new_n1031), .C2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n732), .B1(new_n1036), .B2(new_n749), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT113), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n779), .A2(new_n374), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n319), .A2(new_n767), .B1(new_n759), .B2(new_n205), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G159), .B2(new_n790), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n763), .A2(new_n202), .B1(new_n792), .B2(new_n314), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(KEYINPUT114), .B(G150), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1044), .B1(new_n757), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n262), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n395), .B1(new_n1047), .B2(new_n770), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1041), .A2(new_n1043), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n393), .B1(G326), .B2(new_n757), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n778), .A2(new_n788), .B1(new_n767), .B2(new_n527), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n793), .A2(new_n769), .B1(new_n763), .B2(new_n951), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G322), .B2(new_n790), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n786), .B2(new_n774), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1050), .B1(new_n571), .B2(new_n759), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n747), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1040), .A2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1039), .B(new_n1063), .C1(new_n665), .C2(new_n745), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n998), .A2(new_n1001), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n731), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n804), .A2(new_n1065), .A3(new_n724), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n676), .B(KEYINPUT115), .Z(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n726), .A2(new_n1065), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(G393));
  XNOR2_X1  g0871(.A(new_n988), .B(new_n667), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n731), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n779), .A2(G77), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n774), .A2(new_n372), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n769), .A2(new_n202), .B1(new_n759), .B2(new_n214), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G68), .B2(new_n954), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n395), .B1(new_n757), .B2(G143), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n763), .A2(new_n754), .B1(new_n766), .B2(new_n833), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  OAI22_X1  g0881(.A1(new_n763), .A2(new_n793), .B1(new_n766), .B2(new_n951), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  OAI22_X1  g0883(.A1(new_n769), .A2(new_n786), .B1(new_n759), .B2(new_n206), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n778), .A2(new_n571), .B1(new_n767), .B2(new_n788), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n287), .B1(new_n757), .B2(G322), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n527), .C2(new_n792), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1079), .A2(new_n1081), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n747), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n942), .A2(new_n255), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n749), .B1(new_n675), .B2(new_n542), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n733), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1090), .B(new_n1093), .C1(new_n983), .C2(new_n746), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1072), .B1(new_n726), .B2(new_n1065), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1068), .B1(new_n1067), .B2(new_n992), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1073), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(G390));
  NAND2_X1  g0897(.A1(new_n904), .A2(G330), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(new_n896), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n925), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT39), .B1(new_n870), .B2(new_n886), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n857), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n913), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n812), .B2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1101), .A2(new_n1102), .B1(new_n1105), .B2(new_n924), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n721), .A2(new_n663), .A3(new_n811), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1104), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n857), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n924), .B1(new_n870), .B2(new_n886), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1100), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n922), .A2(new_n925), .B1(new_n914), .B2(new_n923), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1111), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n814), .B(new_n857), .C1(new_n802), .C2(new_n803), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n731), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n743), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n206), .A2(new_n769), .B1(new_n766), .B2(new_n788), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n839), .B(new_n1120), .C1(G87), .C2(new_n954), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n775), .A2(new_n542), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n294), .B1(new_n763), .B2(new_n571), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G294), .B2(new_n757), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1074), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n954), .A2(new_n1045), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT53), .Z(new_n1127));
  INV_X1    g0927(.A(G125), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n753), .A2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n294), .B(new_n1129), .C1(G132), .C2(new_n783), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT116), .Z(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1127), .B(new_n1130), .C1(new_n774), .C2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G128), .A2(new_n790), .B1(new_n760), .B2(G50), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n779), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1135), .B1(new_n769), .B2(new_n968), .C1(new_n1136), .C2(new_n754), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1125), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n747), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n733), .B1(new_n262), .B2(new_n822), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1119), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n904), .A2(G330), .A3(new_n814), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1108), .B1(new_n1142), .B2(new_n1103), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1116), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n814), .B1(new_n802), .B2(new_n803), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1099), .B1(new_n1145), .B2(new_n1103), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n912), .A2(new_n913), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n449), .A2(new_n1098), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n929), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1117), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1068), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1117), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1118), .B(new_n1141), .C1(new_n1152), .C2(new_n1153), .ZN(G378));
  OAI21_X1  g0954(.A(new_n732), .B1(G50), .B2(new_n823), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n282), .A2(new_n862), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n313), .A2(new_n359), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n313), .B2(new_n359), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  OR3_X1    g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1163), .A2(new_n744), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n395), .A2(new_n298), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n535), .A2(new_n792), .B1(new_n788), .B2(new_n753), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(G107), .C2(new_n783), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n954), .A2(G77), .B1(new_n760), .B2(G58), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n770), .A2(G97), .B1(new_n790), .B2(G116), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n962), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT117), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1166), .B1(new_n1172), .B2(KEYINPUT58), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT118), .Z(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(KEYINPUT58), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n766), .A2(new_n1128), .ZN(new_n1176));
  INV_X1    g0976(.A(G128), .ZN(new_n1177));
  INV_X1    g0977(.A(G137), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n763), .A2(new_n1177), .B1(new_n792), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(G132), .C2(new_n770), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n833), .B2(new_n1136), .C1(new_n767), .C2(new_n1133), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n760), .A2(G159), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n757), .C2(G124), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1174), .B(new_n1175), .C1(new_n1182), .C2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1155), .B(new_n1164), .C1(new_n747), .C2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT119), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n927), .A2(new_n926), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1105), .A2(new_n915), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT103), .B1(new_n1191), .B2(new_n911), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n893), .A2(new_n902), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n920), .A2(KEYINPUT40), .A3(new_n898), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1194), .A2(new_n1163), .A3(G330), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1163), .B1(new_n903), .B2(G330), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1193), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n892), .A2(new_n888), .A3(KEYINPUT40), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT104), .B1(new_n901), .B2(new_n852), .ZN(new_n1201));
  OAI211_X1 g1001(.A(G330), .B(new_n1195), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1163), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1204), .A2(new_n1189), .A3(new_n928), .A4(new_n1196), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1199), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1188), .B1(new_n1206), .B2(new_n731), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1204), .A2(new_n1208), .A3(new_n1196), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1208), .B1(new_n1204), .B2(new_n1196), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT57), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1150), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1148), .B2(new_n1117), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1068), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n820), .B1(new_n718), .B2(new_n719), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1100), .B1(new_n1216), .B2(new_n857), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1147), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1217), .A2(new_n1218), .B1(new_n1116), .B2(new_n1143), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1115), .B2(new_n1100), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1150), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1207), .B1(new_n1215), .B2(new_n1223), .ZN(G375));
  NAND2_X1  g1024(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1213), .B(new_n1144), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1005), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1103), .A2(new_n743), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n732), .B1(G68), .B2(new_n823), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n766), .A2(new_n527), .B1(new_n767), .B2(new_n205), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n963), .B(new_n1230), .C1(G116), .C2(new_n770), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n775), .A2(G107), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n294), .B1(new_n753), .B2(new_n786), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G283), .B2(new_n783), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1231), .A2(new_n1041), .A3(new_n1232), .A4(new_n1234), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1136), .A2(new_n202), .B1(new_n833), .B2(new_n792), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT120), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n764), .A2(new_n759), .B1(new_n767), .B2(new_n754), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G132), .B2(new_n790), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n763), .A2(new_n968), .B1(new_n753), .B2(new_n1177), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(new_n395), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1239), .B(new_n1241), .C1(new_n1133), .C2(new_n769), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1229), .B1(new_n1243), .B2(new_n747), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1148), .A2(new_n731), .B1(new_n1228), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1227), .A2(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT121), .Z(G381));
  XNOR2_X1  g1047(.A(G375), .B(KEYINPUT122), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(G384), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n975), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1006), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1024), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1250), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1118), .A2(new_n1141), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1152), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1153), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1249), .A2(new_n1253), .A3(new_n1257), .ZN(new_n1258));
  OR3_X1    g1058(.A1(new_n1248), .A2(G381), .A3(new_n1258), .ZN(G407));
  NAND2_X1  g1059(.A1(new_n655), .A2(G213), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G407), .B(G213), .C1(new_n1248), .C2(new_n1262), .ZN(G409));
  NAND3_X1  g1063(.A1(new_n1199), .A2(new_n1205), .A3(new_n1005), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT123), .B1(new_n1264), .B2(new_n1214), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n928), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1209), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1188), .B1(new_n1267), .B2(new_n731), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1264), .A2(new_n1214), .A3(KEYINPUT123), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1257), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G378), .B(new_n1207), .C1(new_n1215), .C2(new_n1223), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1068), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1226), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1278), .A2(KEYINPUT60), .A3(new_n1213), .A4(new_n1144), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1245), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n849), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G384), .A2(new_n1245), .A3(new_n1280), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1273), .A2(new_n1260), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT62), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1260), .A2(KEYINPUT125), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1282), .A2(new_n1283), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1261), .A2(G2897), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1289), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1282), .A2(new_n1283), .A3(new_n1291), .A4(new_n1287), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1273), .A2(new_n1260), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1273), .A2(new_n1297), .A3(new_n1260), .A4(new_n1284), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1286), .A2(new_n1295), .A3(new_n1296), .A4(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G390), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(G387), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G390), .B(new_n975), .C1(new_n1006), .C2(new_n1024), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1253), .B2(G390), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(G393), .B(new_n800), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1303), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1301), .A2(new_n1306), .A3(new_n1302), .A4(new_n1304), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1299), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT124), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1285), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT63), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1308), .A2(new_n1296), .A3(new_n1309), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT127), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1308), .A2(new_n1317), .A3(new_n1296), .A4(new_n1309), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1316), .A2(new_n1318), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1285), .A2(new_n1312), .A3(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1314), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1311), .A2(new_n1322), .ZN(G405));
  XNOR2_X1  g1123(.A(G375), .B(G378), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(new_n1310), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1284), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OR2_X1    g1127(.A1(new_n1324), .A2(new_n1310), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1324), .A2(new_n1310), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n1284), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1327), .A2(new_n1330), .ZN(G402));
endmodule


