//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960;
  AND2_X1   g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT7), .ZN(new_n204));
  NOR2_X1   g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206));
  AOI211_X1 g005(.A(KEYINPUT94), .B(new_n205), .C1(KEYINPUT8), .C2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G85gat), .ZN(new_n208));
  INV_X1    g007(.A(G92gat), .ZN(new_n209));
  AOI22_X1  g008(.A1(KEYINPUT8), .A2(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT94), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n204), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G99gat), .B(G106gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(new_n204), .C1(new_n207), .C2(new_n212), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT95), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT95), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n213), .A2(new_n219), .A3(new_n215), .ZN(new_n220));
  NAND2_X1  g019(.A1(G71gat), .A2(G78gat), .ZN(new_n221));
  OR2_X1    g020(.A1(G71gat), .A2(G78gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G64gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G57gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT92), .ZN(new_n227));
  INV_X1    g026(.A(G57gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G64gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT91), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n224), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n226), .A2(new_n229), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n221), .B(new_n222), .C1(new_n232), .C2(new_n223), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n220), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n234), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(new_n216), .A3(new_n217), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n220), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT10), .A3(new_n236), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n202), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n235), .A2(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n202), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G120gat), .B(G148gat), .ZN(new_n248));
  INV_X1    g047(.A(G176gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G204gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n244), .A2(new_n246), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259));
  INV_X1    g058(.A(G141gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(G148gat), .ZN(new_n261));
  INV_X1    g060(.A(G148gat), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT75), .B1(new_n262), .B2(G141gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n260), .A2(G148gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT76), .ZN(new_n266));
  XNOR2_X1  g065(.A(G155gat), .B(G162gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT2), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT76), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n270), .B(new_n261), .C1(new_n263), .C2(new_n264), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n266), .A2(new_n267), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G141gat), .B(G148gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(KEYINPUT2), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n274), .A2(new_n267), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  INV_X1    g076(.A(G127gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G134gat), .ZN(new_n279));
  INV_X1    g078(.A(G134gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G127gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n278), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n283), .B(new_n284), .C1(KEYINPUT1), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  INV_X1    g086(.A(G120gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G113gat), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G120gat), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT1), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n284), .A4(new_n283), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n291), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n292), .A2(KEYINPUT68), .A3(new_n298), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n272), .A2(new_n306), .A3(new_n275), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n277), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n305), .A2(KEYINPUT4), .A3(new_n276), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n302), .A2(new_n303), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n287), .B2(new_n295), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n272), .A2(new_n275), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n258), .B(new_n308), .C1(new_n309), .C2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n313), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n305), .A2(new_n276), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n258), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT4), .B1(new_n305), .B2(new_n276), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(new_n313), .A3(new_n310), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n276), .A2(KEYINPUT3), .B1(new_n296), .B2(new_n304), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n321), .A2(new_n322), .B1(new_n323), .B2(new_n307), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n320), .B1(new_n324), .B2(new_n258), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n317), .B1(new_n325), .B2(new_n316), .ZN(new_n326));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT0), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G57gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(new_n208), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n257), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(new_n317), .C1(new_n325), .C2(new_n316), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n257), .ZN(new_n335));
  OR3_X1    g134(.A1(new_n326), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G226gat), .ZN(new_n338));
  INV_X1    g137(.A(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT24), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(new_n342), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  OR2_X1    g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(KEYINPUT24), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G169gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n249), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n343), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT64), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT25), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT25), .B1(new_n352), .B2(KEYINPUT23), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n343), .A2(new_n346), .A3(new_n350), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT26), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT65), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n348), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT65), .B1(new_n365), .B2(new_n352), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT26), .B1(new_n354), .B2(new_n355), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n345), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT27), .B(G183gat), .ZN(new_n370));
  INV_X1    g169(.A(G190gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT28), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n357), .B(new_n359), .C1(new_n369), .C2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n340), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT73), .B(KEYINPUT22), .Z(new_n381));
  INV_X1    g180(.A(G211gat), .ZN(new_n382));
  INV_X1    g181(.A(G218gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G197gat), .B(G204gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G211gat), .B(G218gat), .Z(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n377), .A2(new_n340), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n380), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n377), .A2(KEYINPUT74), .A3(new_n340), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n379), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n391), .B1(new_n395), .B2(new_n389), .ZN(new_n396));
  XNOR2_X1  g195(.A(G8gat), .B(G36gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(new_n225), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(new_n209), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n391), .B(new_n399), .C1(new_n395), .C2(new_n389), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT30), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(KEYINPUT30), .ZN(new_n404));
  INV_X1    g203(.A(new_n394), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT74), .B1(new_n377), .B2(new_n340), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n380), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n388), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n399), .B1(new_n408), .B2(new_n391), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  INV_X1    g211(.A(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT79), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n415), .B(KEYINPUT31), .Z(new_n416));
  AND2_X1   g215(.A1(new_n416), .A2(KEYINPUT81), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(KEYINPUT81), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n386), .A2(new_n387), .ZN(new_n420));
  INV_X1    g219(.A(new_n387), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n384), .B2(new_n385), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n378), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n313), .B1(new_n423), .B2(new_n306), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G22gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n307), .A2(new_n378), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n389), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n388), .B1(new_n378), .B2(new_n307), .ZN(new_n430));
  OAI21_X1  g229(.A(G22gat), .B1(new_n430), .B2(new_n424), .ZN(new_n431));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n430), .B2(KEYINPUT80), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n429), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n429), .B2(new_n431), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n419), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n429), .A2(new_n431), .ZN(new_n437));
  INV_X1    g236(.A(new_n433), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n429), .A2(new_n431), .A3(new_n433), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n418), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n436), .A2(new_n441), .A3(KEYINPUT82), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n337), .A2(new_n411), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n318), .A2(new_n319), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(G225gat), .A3(G233gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n316), .B1(new_n315), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT5), .B1(new_n324), .B2(new_n258), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT84), .B(new_n317), .C1(new_n325), .C2(new_n316), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n332), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n331), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n333), .A2(new_n335), .ZN(new_n456));
  INV_X1    g255(.A(new_n390), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n388), .B1(new_n457), .B2(new_n379), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT37), .B(new_n458), .C1(new_n407), .C2(new_n388), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT38), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n400), .B1(new_n396), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n409), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n455), .A2(new_n456), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT85), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n462), .B2(new_n396), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT38), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n455), .A2(new_n464), .A3(new_n469), .A4(new_n456), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n404), .A2(new_n409), .ZN(new_n473));
  INV_X1    g272(.A(new_n396), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n474), .A2(KEYINPUT30), .A3(new_n399), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n403), .A2(new_n410), .A3(KEYINPUT83), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OR3_X1    g277(.A1(new_n324), .A2(KEYINPUT39), .A3(new_n258), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n318), .A2(new_n319), .A3(new_n258), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT39), .B(new_n480), .C1(new_n324), .C2(new_n258), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n330), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT40), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n479), .A2(new_n484), .A3(new_n330), .A4(new_n481), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n486), .A2(new_n454), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n442), .B1(new_n478), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n446), .B1(new_n471), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n369), .A2(new_n376), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n357), .A2(new_n359), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n305), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n312), .A2(new_n377), .ZN(new_n493));
  INV_X1    g292(.A(G227gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(new_n339), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT32), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT33), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G43gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT69), .ZN(new_n501));
  XOR2_X1   g300(.A(G71gat), .B(G99gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n496), .B(KEYINPUT32), .C1(new_n498), .C2(new_n503), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n495), .B1(new_n492), .B2(new_n493), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n510), .B2(KEYINPUT70), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n508), .A2(new_n509), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n516), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT36), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT72), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n520), .A3(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n517), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT36), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n489), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n334), .A2(new_n336), .B1(new_n410), .B2(new_n403), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n442), .B1(new_n526), .B2(new_n525), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n476), .A2(new_n477), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n533), .A2(new_n535), .A3(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n455), .A2(new_n456), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n256), .B1(new_n530), .B2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G43gat), .B(G50gat), .Z(new_n541));
  INV_X1    g340(.A(KEYINPUT15), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(G29gat), .A2(G36gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT14), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT14), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n548), .A2(KEYINPUT86), .ZN(new_n549));
  NAND2_X1  g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n548), .B2(KEYINPUT86), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n543), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n541), .A2(new_n542), .ZN(new_n553));
  INV_X1    g352(.A(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n541), .A2(new_n542), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n550), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(new_n220), .A3(new_n218), .ZN(new_n559));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT96), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n241), .A2(new_n557), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n559), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT97), .ZN(new_n566));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n559), .A2(new_n563), .A3(new_n564), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n561), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n565), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n573), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT20), .Z(new_n579));
  XNOR2_X1  g378(.A(G15gat), .B(G22gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT16), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(G1gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(G1gat), .B2(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT87), .ZN(new_n584));
  INV_X1    g383(.A(G8gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT87), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT88), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(G8gat), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n236), .A2(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT93), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT93), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(new_n595), .A3(new_n592), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(KEYINPUT19), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT19), .B1(new_n594), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n579), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n596), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT19), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n579), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n597), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n236), .A2(KEYINPUT21), .ZN(new_n606));
  XOR2_X1   g405(.A(G183gat), .B(G211gat), .Z(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n606), .B(new_n609), .Z(new_n610));
  NAND3_X1  g409(.A1(new_n600), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n600), .B2(new_n605), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n577), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT98), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n605), .ZN(new_n616));
  INV_X1    g415(.A(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n611), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n577), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n591), .A2(new_n558), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT90), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n589), .A2(new_n590), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n557), .ZN(new_n627));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n623), .A2(new_n625), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT89), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT90), .B1(new_n630), .B2(new_n624), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n589), .A2(new_n552), .A3(new_n556), .A4(new_n590), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n628), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n623), .A2(new_n631), .A3(new_n627), .A4(new_n628), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n633), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G197gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT11), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n347), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n633), .A2(new_n645), .A3(new_n638), .A4(new_n639), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n540), .A2(new_n622), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n337), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(G1gat), .Z(G1324gat));
  NAND4_X1  g451(.A1(new_n540), .A2(new_n622), .A3(new_n649), .A4(new_n478), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT16), .B(G8gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n656), .B(KEYINPUT100), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n654), .B1(new_n653), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n653), .A2(G8gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT103), .ZN(G1325gat));
  INV_X1    g465(.A(G15gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n518), .A2(new_n521), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(new_n650), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT104), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n525), .A2(new_n527), .A3(new_n526), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n527), .B1(new_n525), .B2(new_n526), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n522), .A2(KEYINPUT105), .A3(new_n528), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n650), .A2(new_n667), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n670), .A2(new_n677), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n444), .A2(new_n445), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n650), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n530), .A2(new_n539), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n684), .B1(new_n685), .B2(new_n576), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n538), .B1(new_n489), .B2(new_n676), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n576), .B(KEYINPUT108), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n649), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n256), .B(KEYINPUT106), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR4_X1   g493(.A1(new_n691), .A2(new_n619), .A3(new_n692), .A4(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G29gat), .B1(new_n696), .B2(new_n337), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n612), .A2(new_n613), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n540), .A2(new_n576), .A3(new_n698), .A4(new_n649), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n699), .A2(G29gat), .A3(new_n337), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT45), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(G1328gat));
  OAI21_X1  g501(.A(G36gat), .B1(new_n696), .B2(new_n535), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n699), .A2(G36gat), .A3(new_n535), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  OAI21_X1  g506(.A(G43gat), .B1(new_n696), .B2(new_n676), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n699), .A2(G43gat), .A3(new_n668), .ZN(new_n709));
  AOI211_X1 g508(.A(KEYINPUT109), .B(new_n707), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n707), .A2(KEYINPUT109), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(KEYINPUT109), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n711), .A2(new_n708), .A3(new_n712), .A4(new_n709), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n710), .A2(new_n713), .ZN(G1330gat));
  INV_X1    g513(.A(new_n442), .ZN(new_n715));
  OAI21_X1  g514(.A(G50gat), .B1(new_n696), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n699), .A2(G50gat), .A3(new_n680), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(KEYINPUT48), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n695), .A2(new_n679), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(G50gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n721), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g521(.A(new_n687), .ZN(new_n723));
  AND4_X1   g522(.A1(new_n622), .A2(new_n723), .A3(new_n692), .A4(new_n694), .ZN(new_n724));
  INV_X1    g523(.A(new_n337), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g526(.A(new_n535), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT110), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n730), .B(new_n731), .Z(G1333gat));
  INV_X1    g531(.A(new_n676), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n724), .A2(G71gat), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n668), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n724), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n736), .B2(G71gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n724), .A2(new_n679), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g539(.A1(new_n686), .A2(new_n690), .ZN(new_n741));
  INV_X1    g540(.A(new_n256), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n619), .A2(new_n649), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G85gat), .B1(new_n744), .B2(new_n337), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n698), .A2(new_n576), .A3(new_n692), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n471), .A2(new_n488), .ZN(new_n748));
  INV_X1    g547(.A(new_n446), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n749), .A3(new_n676), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n747), .B1(new_n750), .B2(new_n539), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT111), .B1(new_n751), .B2(KEYINPUT51), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NOR4_X1   g553(.A1(new_n687), .A2(new_n753), .A3(new_n754), .A4(new_n747), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n746), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n687), .B2(new_n747), .ZN(new_n757));
  INV_X1    g556(.A(new_n747), .ZN(new_n758));
  AOI221_X4 g557(.A(new_n446), .B1(new_n674), .B2(new_n675), .C1(new_n471), .C2(new_n488), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT51), .B(new_n758), .C1(new_n759), .C2(new_n538), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n753), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n751), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(KEYINPUT112), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n756), .A2(new_n757), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n208), .A3(new_n725), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n745), .B1(new_n765), .B2(new_n742), .ZN(G1336gat));
  NOR3_X1   g565(.A1(new_n693), .A2(G92gat), .A3(new_n535), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT113), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n478), .B(new_n743), .C1(new_n686), .C2(new_n690), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n209), .B1(new_n770), .B2(KEYINPUT114), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n741), .A2(new_n772), .A3(new_n478), .A4(new_n743), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n764), .A2(new_n775), .A3(new_n767), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n769), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n770), .A2(G92gat), .ZN(new_n778));
  INV_X1    g577(.A(new_n757), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n761), .B2(new_n762), .ZN(new_n780));
  INV_X1    g579(.A(new_n767), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT52), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT115), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n777), .A2(new_n786), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n744), .B2(new_n676), .ZN(new_n789));
  INV_X1    g588(.A(G99gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n764), .A2(new_n790), .A3(new_n256), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n791), .B2(new_n668), .ZN(G1338gat));
  NAND3_X1  g591(.A1(new_n741), .A2(new_n679), .A3(new_n743), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n693), .A2(G106gat), .A3(new_n715), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT53), .B1(new_n764), .B2(new_n795), .ZN(new_n799));
  OAI21_X1  g598(.A(G106gat), .B1(new_n744), .B2(new_n715), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1339gat));
  INV_X1    g601(.A(KEYINPUT108), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n576), .B(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n254), .B1(new_n243), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n240), .A2(new_n202), .A3(new_n242), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n243), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT116), .B1(new_n808), .B2(KEYINPUT54), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  NOR4_X1   g609(.A1(new_n807), .A2(new_n243), .A3(new_n810), .A4(new_n805), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT55), .B(new_n806), .C1(new_n809), .C2(new_n811), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n649), .A3(new_n255), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n635), .A2(new_n637), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n628), .B1(new_n623), .B2(new_n627), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n644), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT117), .B(new_n644), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n822), .A2(new_n648), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n256), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n804), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n816), .A2(new_n255), .A3(new_n824), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n689), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n698), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n615), .A2(new_n621), .A3(new_n692), .A4(new_n742), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n829), .B2(new_n830), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n832), .A2(new_n833), .A3(new_n478), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n725), .ZN(new_n835));
  INV_X1    g634(.A(new_n533), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n838), .A2(new_n290), .A3(new_n649), .A4(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n835), .A2(new_n679), .A3(new_n668), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n692), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(G1340gat));
  NAND4_X1  g643(.A1(new_n838), .A2(new_n288), .A3(new_n256), .A4(new_n839), .ZN(new_n845));
  OAI21_X1  g644(.A(G120gat), .B1(new_n842), .B2(new_n693), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1341gat));
  AOI21_X1  g646(.A(G127gat), .B1(new_n837), .B2(new_n619), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n698), .A2(new_n278), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n841), .B2(new_n849), .ZN(G1342gat));
  NAND3_X1  g649(.A1(new_n837), .A2(new_n280), .A3(new_n576), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n852));
  OAI21_X1  g651(.A(G134gat), .B1(new_n842), .B2(new_n577), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(G1343gat));
  NOR3_X1   g654(.A1(new_n832), .A2(new_n833), .A3(new_n715), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n733), .A2(new_n337), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n692), .A2(G141gat), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n535), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n856), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n814), .A2(new_n255), .A3(new_n815), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n814), .A2(new_n255), .A3(new_n868), .A4(new_n815), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n649), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n576), .B1(new_n870), .B2(new_n825), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n698), .B1(new_n871), .B2(new_n828), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n830), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT57), .B1(new_n873), .B2(new_n680), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n535), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n865), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G141gat), .B1(new_n877), .B2(new_n692), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n856), .A2(new_n876), .A3(new_n861), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n881), .B2(new_n863), .ZN(G1344gat));
  NAND4_X1  g681(.A1(new_n860), .A2(new_n262), .A3(new_n535), .A4(new_n256), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n865), .A2(new_n256), .A3(new_n874), .A4(new_n876), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(G148gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n884), .A2(KEYINPUT122), .A3(new_n885), .A4(G148gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n827), .A2(new_n577), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n871), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n871), .B2(new_n892), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n698), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n830), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT124), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n895), .A2(new_n898), .A3(new_n830), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n897), .A2(new_n899), .A3(new_n864), .A4(new_n679), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n856), .A2(new_n864), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n256), .A4(new_n876), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n885), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n883), .B1(new_n890), .B2(new_n903), .ZN(G1345gat));
  NAND3_X1  g703(.A1(new_n860), .A2(new_n619), .A3(new_n535), .ZN(new_n905));
  INV_X1    g704(.A(G155gat), .ZN(new_n906));
  INV_X1    g705(.A(new_n877), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n698), .A2(new_n906), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT125), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n905), .A2(new_n906), .B1(new_n907), .B2(new_n909), .ZN(G1346gat));
  XOR2_X1   g709(.A(KEYINPUT77), .B(G162gat), .Z(new_n911));
  NAND4_X1  g710(.A1(new_n860), .A2(new_n576), .A3(new_n535), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n907), .A2(KEYINPUT126), .A3(new_n804), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n877), .B2(new_n689), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n912), .B1(new_n916), .B2(new_n911), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n832), .A2(new_n833), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n725), .A2(new_n535), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n918), .A2(new_n680), .A3(new_n735), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G169gat), .B1(new_n920), .B2(new_n692), .ZN(new_n921));
  INV_X1    g720(.A(new_n919), .ZN(new_n922));
  NOR4_X1   g721(.A1(new_n832), .A2(new_n833), .A3(new_n836), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n347), .A3(new_n649), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(G1348gat));
  OAI21_X1  g724(.A(G176gat), .B1(new_n920), .B2(new_n693), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n249), .A3(new_n256), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT127), .ZN(G1349gat));
  OAI21_X1  g728(.A(G183gat), .B1(new_n920), .B2(new_n698), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n923), .A2(new_n619), .A3(new_n370), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n923), .A2(new_n371), .A3(new_n804), .ZN(new_n934));
  OAI21_X1  g733(.A(G190gat), .B1(new_n920), .B2(new_n577), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(G1351gat));
  AND2_X1   g738(.A1(new_n900), .A2(new_n901), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n733), .A2(new_n922), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n649), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G197gat), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n856), .A2(new_n941), .ZN(new_n944));
  INV_X1    g743(.A(G197gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n945), .A3(new_n649), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n946), .ZN(G1352gat));
  NAND3_X1  g746(.A1(new_n940), .A2(new_n694), .A3(new_n941), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G204gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n944), .A2(new_n251), .A3(new_n256), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n944), .A2(new_n382), .A3(new_n619), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n900), .A2(new_n901), .A3(new_n619), .A4(new_n941), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  AOI21_X1  g756(.A(G218gat), .B1(new_n944), .B2(new_n804), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n940), .A2(new_n941), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n577), .A2(new_n383), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(G1355gat));
endmodule


