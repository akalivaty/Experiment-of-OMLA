//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n190), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n188), .B2(G143), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n194), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n193), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT11), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n205), .A2(G134), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n202), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n205), .B2(G134), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(KEYINPUT65), .A3(G134), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n202), .A2(KEYINPUT66), .A3(G137), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n213), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n201), .A2(new_n211), .A3(new_n219), .ZN(new_n220));
  AOI211_X1 g034(.A(G131), .B(new_n209), .C1(new_n203), .C2(new_n206), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n208), .B1(new_n207), .B2(new_n210), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n189), .A2(new_n191), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n198), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n220), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G116), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT67), .A3(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(G116), .ZN(new_n236));
  INV_X1    g050(.A(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT2), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G113), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n235), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT68), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n232), .A2(new_n234), .B1(G116), .B2(new_n231), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n241), .ZN(new_n246));
  OAI22_X1  g060(.A1(new_n243), .A2(new_n246), .B1(new_n245), .B2(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n229), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT71), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n228), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT69), .B(new_n225), .C1(new_n198), .C2(new_n227), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n223), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n245), .A2(new_n241), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n242), .A2(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n245), .A2(new_n244), .A3(new_n241), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n259), .A3(new_n220), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n229), .A2(new_n261), .A3(new_n247), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n249), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT28), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT70), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(G210), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n229), .A2(new_n261), .A3(new_n247), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n261), .B1(new_n229), .B2(new_n247), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n277), .B1(new_n280), .B2(new_n260), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n260), .A2(new_n277), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT72), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n265), .B(new_n276), .C1(new_n281), .C2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n255), .A2(KEYINPUT30), .A3(new_n220), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n229), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n247), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n275), .A3(new_n260), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n275), .A4(new_n260), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G472), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT73), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n298), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n281), .A2(new_n283), .ZN(new_n304));
  INV_X1    g118(.A(new_n265), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n275), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n288), .A2(new_n260), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n276), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n220), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n253), .B2(new_n254), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(new_n247), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n282), .B1(new_n313), .B2(new_n277), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n276), .A2(new_n307), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n295), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n187), .B1(new_n303), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n263), .A2(KEYINPUT28), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT72), .A3(new_n282), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n276), .B1(new_n321), .B2(new_n265), .ZN(new_n322));
  INV_X1    g136(.A(new_n309), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n322), .A2(KEYINPUT29), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n317), .ZN(new_n325));
  OAI21_X1  g139(.A(G472), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n326), .A2(KEYINPUT74), .A3(new_n301), .A4(new_n302), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n270), .A2(G227), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G140), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n333));
  INV_X1    g147(.A(G104), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n333), .A2(KEYINPUT3), .B1(new_n334), .B2(G107), .ZN(new_n335));
  OAI22_X1  g149(.A1(new_n333), .A2(KEYINPUT3), .B1(new_n334), .B2(G107), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n337));
  INV_X1    g151(.A(G107), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT80), .A4(G104), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G101), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n335), .A2(new_n336), .A3(new_n342), .A4(new_n339), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(KEYINPUT4), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n345), .A3(G101), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n338), .A3(G104), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT81), .B1(new_n338), .B2(G104), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n334), .A2(G107), .ZN(new_n351));
  OAI211_X1 g165(.A(G101), .B(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n193), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n199), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n189), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n357), .A2(new_n358), .B1(new_n189), .B2(new_n191), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n353), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n347), .A2(new_n253), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n353), .A2(KEYINPUT10), .A3(new_n201), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(KEYINPUT84), .A3(new_n223), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n253), .A2(new_n346), .A3(new_n344), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n361), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n223), .A4(new_n363), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n332), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n362), .A2(new_n363), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n254), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n360), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n353), .A2(new_n201), .ZN(new_n375));
  OAI211_X1 g189(.A(KEYINPUT12), .B(new_n254), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n254), .B1(new_n374), .B2(new_n375), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n364), .A2(new_n369), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n332), .B1(new_n380), .B2(KEYINPUT85), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n364), .A2(new_n369), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n376), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n382), .A2(KEYINPUT85), .A3(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(G469), .B(new_n373), .C1(new_n381), .C2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G469), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n370), .A2(new_n383), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n331), .B1(new_n382), .B2(new_n372), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n386), .B(new_n296), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(G469), .A2(G902), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT9), .B(G234), .Z(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G221), .B1(new_n393), .B2(G902), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n397));
  INV_X1    g211(.A(G125), .ZN(new_n398));
  OR3_X1    g212(.A1(new_n398), .A2(KEYINPUT16), .A3(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT76), .B1(new_n400), .B2(new_n188), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(G146), .A3(new_n399), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT24), .B(G110), .Z(new_n404));
  XNOR2_X1  g218(.A(G119), .B(G128), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT23), .B1(new_n199), .B2(G119), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n199), .A2(G119), .ZN(new_n408));
  MUX2_X1   g222(.A(KEYINPUT23), .B(new_n407), .S(new_n408), .Z(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G110), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n397), .A2(KEYINPUT76), .A3(G146), .A4(new_n399), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n403), .A2(new_n406), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  OAI22_X1  g226(.A1(new_n409), .A2(G110), .B1(new_n405), .B2(new_n404), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n396), .A2(new_n188), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n402), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT22), .B(G137), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n417), .A2(KEYINPUT77), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n417), .A2(KEYINPUT77), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n418), .B2(new_n420), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n421), .A2(KEYINPUT78), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT78), .B1(new_n421), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n422), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n412), .A2(new_n427), .A3(new_n415), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n296), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT25), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT75), .B(G217), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(G234), .B2(new_n296), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G902), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT79), .Z(new_n436));
  AND2_X1   g250(.A1(new_n426), .A2(new_n428), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n431), .A2(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n395), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n235), .A2(KEYINPUT5), .A3(new_n236), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n236), .A2(KEYINPUT5), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(G113), .A3(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n353), .B(new_n444), .C1(new_n243), .C2(new_n246), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n344), .A2(new_n346), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n445), .B(new_n446), .C1(new_n447), .C2(new_n259), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n228), .A2(G125), .ZN(new_n449));
  INV_X1    g263(.A(G224), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(G953), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n398), .B(new_n193), .C1(new_n198), .C2(new_n200), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n449), .A2(KEYINPUT7), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  AOI211_X1 g271(.A(KEYINPUT87), .B(new_n457), .C1(new_n449), .C2(new_n453), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n189), .A2(new_n191), .A3(new_n224), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT64), .B1(new_n190), .B2(G146), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n189), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n224), .A2(new_n226), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n453), .B1(new_n465), .B2(new_n398), .ZN(new_n466));
  INV_X1    g280(.A(new_n457), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n446), .B(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n444), .B1(new_n243), .B2(new_n246), .ZN(new_n472));
  INV_X1    g286(.A(new_n353), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n474), .B2(new_n445), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n455), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n441), .B1(new_n476), .B2(G902), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n445), .B1(new_n447), .B2(new_n259), .ZN(new_n478));
  INV_X1    g292(.A(new_n446), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n448), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n466), .B(new_n451), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n483), .A3(new_n479), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n458), .A2(new_n468), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n474), .A2(new_n445), .ZN(new_n487));
  INV_X1    g301(.A(new_n471), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(KEYINPUT88), .B(new_n296), .C1(new_n490), .C2(new_n455), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n477), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G210), .B1(G237), .B2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n477), .A2(new_n491), .A3(new_n493), .A4(new_n485), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(KEYINPUT89), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G214), .B1(G237), .B2(G902), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n499), .A3(new_n494), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT90), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n497), .A2(new_n503), .A3(new_n498), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n403), .A2(new_n411), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n270), .A2(G214), .A3(new_n271), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n190), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n270), .A2(G143), .A3(G214), .A4(new_n271), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT17), .A3(G131), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(G131), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n208), .A3(new_n509), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n506), .B(new_n511), .C1(new_n514), .C2(KEYINPUT17), .ZN(new_n515));
  XNOR2_X1  g329(.A(G113), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n334), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n508), .B(new_n509), .C1(new_n518), .C2(new_n208), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n396), .B(new_n188), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(new_n520), .C1(new_n512), .C2(new_n518), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n517), .ZN(new_n523));
  INV_X1    g337(.A(new_n521), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n396), .B(KEYINPUT19), .Z(new_n525));
  OAI21_X1  g339(.A(new_n402), .B1(new_n525), .B2(G146), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n512), .B2(new_n513), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n523), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G475), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n296), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT20), .ZN(new_n532));
  AOI21_X1  g346(.A(G475), .B1(new_n522), .B2(new_n528), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT20), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n296), .ZN(new_n535));
  INV_X1    g349(.A(new_n522), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n517), .B1(new_n515), .B2(new_n521), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n296), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n532), .A2(new_n535), .B1(G475), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n544));
  XNOR2_X1  g358(.A(G116), .B(G122), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n545), .A2(new_n546), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(G107), .ZN(new_n550));
  XOR2_X1   g364(.A(G116), .B(G122), .Z(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT91), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n338), .B1(new_n552), .B2(new_n547), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n544), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G128), .B(G143), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n202), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(KEYINPUT13), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n190), .A2(G128), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n557), .B(G134), .C1(KEYINPUT13), .C2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G107), .B1(new_n548), .B2(new_n549), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(new_n547), .A3(new_n338), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(KEYINPUT92), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n554), .A2(new_n556), .A3(new_n559), .A4(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n555), .B(new_n202), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n233), .A2(KEYINPUT14), .A3(G122), .ZN(new_n565));
  OAI211_X1 g379(.A(G107), .B(new_n565), .C1(new_n551), .C2(KEYINPUT14), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n393), .A2(new_n433), .A3(G953), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n563), .B2(new_n567), .ZN(new_n571));
  OAI221_X1 g385(.A(new_n296), .B1(new_n542), .B2(new_n543), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n570), .A2(new_n571), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(G902), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n574), .B2(new_n542), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n539), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(G234), .A2(G237), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n578), .A2(G952), .A3(new_n266), .ZN(new_n579));
  INV_X1    g393(.A(new_n270), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n580), .A2(G902), .A3(new_n578), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT21), .B(G898), .Z(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n328), .A2(new_n440), .A3(new_n505), .A4(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  AOI21_X1  g401(.A(G902), .B1(new_n284), .B2(new_n293), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n588), .A2(new_n295), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n299), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n440), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT94), .ZN(new_n593));
  INV_X1    g407(.A(new_n498), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n492), .A2(new_n494), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n495), .A2(KEYINPUT95), .A3(new_n496), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n540), .A2(new_n296), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n573), .A2(KEYINPUT33), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n570), .B2(new_n571), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n601), .B1(new_n605), .B2(G478), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n574), .A2(new_n540), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n538), .A2(G475), .ZN(new_n609));
  INV_X1    g423(.A(new_n535), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n534), .B1(new_n533), .B2(new_n296), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n584), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n600), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  NAND2_X1  g431(.A1(new_n539), .A2(new_n575), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n584), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n600), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G107), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NAND2_X1  g436(.A1(new_n431), .A2(new_n434), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n425), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n416), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n436), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n395), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n505), .A2(new_n585), .A3(new_n629), .A4(new_n591), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  INV_X1    g446(.A(new_n599), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n579), .B1(new_n581), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n618), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n328), .A2(new_n633), .A3(new_n629), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  XNOR2_X1  g452(.A(new_n635), .B(KEYINPUT39), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n391), .A2(new_n394), .A3(new_n640), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n641), .A2(KEYINPUT40), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n497), .A2(new_n500), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT38), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n644), .A2(new_n594), .A3(new_n627), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n612), .A2(new_n575), .ZN(new_n646));
  INV_X1    g460(.A(new_n303), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n313), .A2(new_n276), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n296), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n276), .B1(new_n288), .B2(new_n260), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n646), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n641), .A2(KEYINPUT40), .ZN(new_n653));
  AND4_X1   g467(.A1(new_n642), .A2(new_n645), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n190), .ZN(G45));
  NOR2_X1   g469(.A1(new_n613), .A2(new_n635), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n328), .A2(new_n633), .A3(new_n629), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G146), .ZN(G48));
  NAND2_X1  g472(.A1(new_n382), .A2(new_n372), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n659), .A2(new_n332), .B1(new_n370), .B2(new_n383), .ZN(new_n660));
  OAI21_X1  g474(.A(G469), .B1(new_n660), .B2(G902), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n661), .A2(new_n389), .A3(new_n394), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n662), .A2(new_n597), .A3(new_n598), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n328), .A2(new_n438), .A3(new_n614), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT41), .B(G113), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G15));
  NAND4_X1  g480(.A1(new_n328), .A2(new_n438), .A3(new_n619), .A4(new_n663), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G116), .ZN(G18));
  NAND4_X1  g482(.A1(new_n328), .A2(new_n585), .A3(new_n627), .A4(new_n663), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G119), .ZN(G21));
  NOR2_X1   g484(.A1(new_n539), .A2(new_n576), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n662), .A2(new_n597), .A3(new_n671), .A4(new_n598), .ZN(new_n672));
  INV_X1    g486(.A(new_n584), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n293), .B1(new_n315), .B2(new_n275), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n298), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n589), .A2(new_n438), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT96), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n598), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n498), .B1(new_n495), .B2(KEYINPUT95), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n678), .A2(new_n646), .A3(new_n679), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n675), .B(new_n438), .C1(new_n295), .C2(new_n588), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n584), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT96), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n680), .A2(new_n682), .A3(new_n683), .A4(new_n662), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT97), .B(G122), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G24));
  NAND3_X1  g501(.A1(new_n589), .A2(new_n627), .A3(new_n675), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT98), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n589), .A2(new_n627), .A3(KEYINPUT98), .A4(new_n675), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n656), .A3(new_n663), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  AOI21_X1  g508(.A(new_n439), .B1(new_n319), .B2(new_n327), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n643), .B2(new_n498), .ZN(new_n698));
  AOI211_X1 g512(.A(KEYINPUT100), .B(new_n594), .C1(new_n497), .C2(new_n500), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n390), .B(KEYINPUT99), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n385), .A2(new_n389), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n394), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n696), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT101), .A4(new_n703), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n656), .B(new_n695), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n656), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n643), .A2(new_n498), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n643), .A2(new_n697), .A3(new_n498), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n704), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT101), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n700), .A2(new_n696), .A3(new_n704), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n710), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n439), .B1(new_n647), .B2(new_n326), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n707), .A2(new_n709), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n208), .ZN(G33));
  NAND2_X1  g535(.A1(new_n715), .A2(new_n716), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n636), .A3(new_n695), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G134), .ZN(G36));
  NAND2_X1  g538(.A1(new_n608), .A2(new_n539), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT43), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n590), .A3(new_n627), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n700), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n381), .A2(new_n384), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n373), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(KEYINPUT45), .A3(new_n373), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(G469), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(KEYINPUT46), .A3(new_n701), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n389), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT46), .B1(new_n737), .B2(new_n701), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n394), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n730), .A2(new_n731), .A3(new_n639), .A4(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT103), .B(G137), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G39));
  INV_X1    g558(.A(new_n741), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT47), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n741), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n328), .ZN(new_n750));
  INV_X1    g564(.A(new_n700), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n710), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n749), .A2(new_n750), .A3(new_n439), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n328), .B1(new_n746), .B2(new_n748), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n756), .A3(new_n439), .A4(new_n752), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  OAI211_X1 g573(.A(new_n656), .B(new_n692), .C1(new_n705), .C2(new_n706), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n722), .A2(KEYINPUT108), .A3(new_n656), .A4(new_n692), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n762), .A2(new_n723), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n720), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n664), .A2(new_n667), .A3(new_n669), .A4(new_n685), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n590), .A2(new_n395), .A3(new_n439), .ZN(new_n767));
  INV_X1    g581(.A(new_n619), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n502), .B2(new_n504), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n769), .B2(KEYINPUT107), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n771), .B(new_n768), .C1(new_n502), .C2(new_n504), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n630), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n613), .B(KEYINPUT106), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n673), .A3(new_n505), .A4(new_n767), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n586), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n577), .A2(new_n635), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n700), .A2(new_n328), .A3(new_n629), .A4(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n766), .A2(new_n773), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n635), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n704), .A2(KEYINPUT109), .A3(new_n628), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n628), .A2(new_n702), .A3(new_n394), .A4(new_n781), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n782), .A2(new_n652), .A3(new_n633), .A4(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n637), .A2(new_n657), .A3(new_n786), .A4(new_n693), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n764), .A2(new_n765), .A3(new_n780), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n762), .A2(new_n723), .A3(new_n763), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n664), .A2(new_n667), .A3(new_n669), .A4(new_n685), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n585), .A2(new_n505), .A3(new_n591), .A4(new_n629), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n505), .A2(new_n619), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n592), .B1(new_n796), .B2(new_n771), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n769), .A2(KEYINPUT107), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n775), .A2(new_n586), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n794), .A2(new_n799), .A3(new_n800), .A4(new_n778), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n793), .A2(new_n801), .A3(new_n720), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n637), .A2(new_n657), .A3(new_n693), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT110), .A3(KEYINPUT52), .A4(new_n786), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n787), .B2(new_n788), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n787), .A2(new_n788), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n802), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n792), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n764), .A2(new_n808), .A3(new_n765), .A4(new_n780), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n791), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n802), .A2(KEYINPUT53), .A3(new_n789), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT112), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n816), .A2(new_n817), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n820), .B(new_n812), .C1(new_n821), .C2(new_n814), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n644), .A2(new_n394), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n661), .A2(new_n389), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n579), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n681), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n727), .A2(new_n594), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT50), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n726), .A2(new_n828), .A3(new_n498), .A4(new_n681), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n826), .A4(new_n825), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n751), .A2(new_n828), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n662), .A3(new_n692), .A4(new_n727), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n647), .A2(new_n438), .A3(new_n651), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n608), .A2(new_n612), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n835), .A2(new_n662), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n831), .A2(new_n834), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n726), .A2(new_n828), .A3(new_n681), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n826), .B(KEYINPUT105), .Z(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n394), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n700), .B(new_n843), .C1(new_n749), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n842), .A2(KEYINPUT51), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  INV_X1    g664(.A(new_n846), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n850), .B1(new_n851), .B2(new_n840), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n842), .A2(KEYINPUT114), .A3(KEYINPUT51), .A4(new_n846), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n849), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n835), .A2(new_n662), .A3(new_n718), .A4(new_n727), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT48), .ZN(new_n856));
  INV_X1    g670(.A(G952), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n857), .B(G953), .C1(new_n843), .C2(new_n663), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n835), .A2(new_n662), .A3(new_n837), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n856), .B(new_n858), .C1(new_n613), .C2(new_n859), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT115), .Z(new_n861));
  NAND4_X1  g675(.A1(new_n823), .A2(new_n824), .A3(new_n854), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(new_n266), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n854), .A2(new_n819), .A3(new_n822), .A4(new_n861), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT116), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n594), .B(new_n725), .C1(new_n844), .C2(KEYINPUT49), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n844), .A2(KEYINPUT49), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n837), .A3(new_n825), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n866), .A2(new_n869), .ZN(G75));
  AOI21_X1  g684(.A(new_n296), .B1(new_n792), .B2(new_n809), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n871), .B2(G210), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n481), .A2(new_n484), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(new_n482), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n872), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n270), .A2(G952), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT117), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(G51));
  NOR2_X1   g693(.A1(new_n815), .A2(new_n791), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT53), .B1(new_n802), .B2(new_n789), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n810), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT119), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n792), .A2(new_n809), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n810), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n812), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n792), .A2(new_n809), .A3(KEYINPUT118), .A4(new_n811), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n883), .A2(new_n886), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n701), .B(KEYINPUT57), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n660), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n890), .A2(KEYINPUT120), .A3(new_n891), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n737), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n871), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n877), .B1(new_n897), .B2(new_n899), .ZN(G54));
  NAND3_X1  g714(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(new_n529), .Z(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n877), .ZN(G60));
  XNOR2_X1  g717(.A(new_n601), .B(KEYINPUT59), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n605), .B1(new_n823), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n878), .ZN(new_n906));
  INV_X1    g720(.A(new_n904), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n890), .A2(new_n604), .A3(new_n602), .A4(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT60), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n792), .B2(new_n809), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n437), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n878), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n625), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n914), .B(new_n915), .C1(KEYINPUT121), .C2(KEYINPUT61), .ZN(new_n916));
  NAND2_X1  g730(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G66));
  OAI21_X1  g732(.A(G953), .B1(new_n583), .B2(new_n450), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n766), .A2(new_n773), .A3(new_n776), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n580), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n873), .B1(G898), .B2(new_n270), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT122), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n921), .B(new_n923), .ZN(G69));
  NAND4_X1  g738(.A1(new_n745), .A2(new_n640), .A3(new_n680), .A4(new_n718), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n803), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n742), .A2(new_n926), .A3(new_n720), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n758), .A2(new_n723), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT127), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n758), .A2(new_n927), .A3(new_n930), .A4(new_n723), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n270), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n285), .A2(new_n287), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(new_n525), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n580), .A2(G900), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n654), .B1(new_n938), .B2(KEYINPUT62), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n803), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT124), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n742), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n940), .A2(new_n942), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n774), .B1(new_n539), .B2(new_n575), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n641), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n695), .A3(new_n700), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n758), .A2(new_n943), .A3(new_n944), .A4(new_n947), .ZN(new_n948));
  AOI22_X1  g762(.A1(new_n948), .A2(new_n270), .B1(KEYINPUT123), .B2(new_n934), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n934), .A2(KEYINPUT123), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n949), .A2(KEYINPUT125), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT125), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n937), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n270), .B1(G227), .B2(G900), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n937), .B2(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OAI221_X1 g770(.A(new_n937), .B1(KEYINPUT126), .B2(new_n954), .C1(new_n951), .C2(new_n952), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  INV_X1    g774(.A(new_n920), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n948), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n650), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(G952), .B2(new_n270), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n929), .A2(new_n920), .A3(new_n931), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n275), .B(new_n308), .C1(new_n965), .C2(new_n960), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n821), .B1(new_n289), .B2(new_n309), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n964), .B(new_n966), .C1(new_n960), .C2(new_n967), .ZN(G57));
endmodule


