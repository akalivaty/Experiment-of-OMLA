

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792;

  BUF_X1 U379 ( .A(n712), .Z(n357) );
  NAND2_X1 U380 ( .A1(n369), .A2(n412), .ZN(n588) );
  AND2_X1 U381 ( .A1(n627), .A2(n575), .ZN(n582) );
  XNOR2_X1 U382 ( .A(n778), .B(G146), .ZN(n568) );
  XNOR2_X1 U383 ( .A(G902), .B(KEYINPUT15), .ZN(n662) );
  BUF_X1 U384 ( .A(G116), .Z(n360) );
  XOR2_X2 U385 ( .A(n684), .B(n683), .Z(n377) );
  XOR2_X2 U386 ( .A(n673), .B(n672), .Z(n379) );
  XOR2_X2 U387 ( .A(n678), .B(n677), .Z(n380) );
  INV_X2 U388 ( .A(G116), .ZN(n438) );
  OR2_X2 U389 ( .A1(n684), .A2(G902), .ZN(n570) );
  XNOR2_X1 U390 ( .A(n622), .B(KEYINPUT39), .ZN(n657) );
  XOR2_X1 U391 ( .A(G119), .B(G128), .Z(n358) );
  AND2_X1 U392 ( .A1(n461), .A2(n670), .ZN(n359) );
  AND2_X2 U393 ( .A1(n420), .A2(n600), .ZN(n419) );
  AND2_X2 U394 ( .A1(n435), .A2(n474), .ZN(n473) );
  NAND2_X2 U395 ( .A1(n594), .A2(n574), .ZN(n721) );
  XNOR2_X2 U396 ( .A(n502), .B(n501), .ZN(n594) );
  NAND2_X2 U397 ( .A1(n462), .A2(n478), .ZN(n461) );
  NAND2_X2 U398 ( .A1(n463), .A2(n461), .ZN(n407) );
  AND2_X2 U399 ( .A1(n464), .A2(n479), .ZN(n463) );
  BUF_X2 U400 ( .A(n752), .Z(n759) );
  XNOR2_X2 U401 ( .A(n520), .B(n511), .ZN(n778) );
  XNOR2_X2 U402 ( .A(n554), .B(KEYINPUT4), .ZN(n520) );
  NOR2_X1 U403 ( .A1(n368), .A2(n398), .ZN(n397) );
  OR2_X1 U404 ( .A1(n644), .A2(n643), .ZN(n368) );
  AND2_X1 U405 ( .A1(n392), .A2(n593), .ZN(n692) );
  AND2_X1 U406 ( .A1(n415), .A2(n410), .ZN(n369) );
  INV_X2 U407 ( .A(n642), .ZN(n695) );
  NOR2_X1 U408 ( .A1(n721), .A2(n616), .ZN(n618) );
  XNOR2_X1 U409 ( .A(n386), .B(G478), .ZN(n572) );
  XNOR2_X1 U410 ( .A(n467), .B(n558), .ZN(n757) );
  INV_X1 U411 ( .A(n567), .ZN(n441) );
  XNOR2_X1 U412 ( .A(n443), .B(n442), .ZN(n567) );
  INV_X2 U413 ( .A(G953), .ZN(n516) );
  INV_X1 U414 ( .A(n401), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n624), .B(n623), .ZN(n682) );
  XNOR2_X2 U416 ( .A(n452), .B(KEYINPUT19), .ZN(n634) );
  NAND2_X2 U417 ( .A1(n608), .A2(n714), .ZN(n452) );
  NAND2_X1 U418 ( .A1(n392), .A2(n593), .ZN(n362) );
  NAND2_X1 U419 ( .A1(n661), .A2(n709), .ZN(n428) );
  BUF_X1 U420 ( .A(n608), .Z(n652) );
  XNOR2_X1 U421 ( .A(n363), .B(KEYINPUT106), .ZN(n392) );
  NOR2_X1 U422 ( .A1(n592), .A2(n650), .ZN(n363) );
  XNOR2_X2 U423 ( .A(n364), .B(n365), .ZN(n712) );
  NAND2_X1 U424 ( .A1(n582), .A2(n650), .ZN(n364) );
  XNOR2_X1 U425 ( .A(KEYINPUT107), .B(KEYINPUT33), .ZN(n365) );
  XNOR2_X2 U426 ( .A(n428), .B(n481), .ZN(n477) );
  XNOR2_X2 U427 ( .A(n765), .B(n469), .ZN(n676) );
  XNOR2_X1 U428 ( .A(n764), .B(KEYINPUT69), .ZN(n521) );
  XNOR2_X1 U429 ( .A(n652), .B(KEYINPUT38), .ZN(n406) );
  INV_X1 U430 ( .A(n598), .ZN(n389) );
  NAND2_X1 U431 ( .A1(n432), .A2(n367), .ZN(n669) );
  INV_X1 U432 ( .A(KEYINPUT72), .ZN(n480) );
  INV_X1 U433 ( .A(KEYINPUT79), .ZN(n481) );
  XNOR2_X1 U434 ( .A(n457), .B(n456), .ZN(n535) );
  XNOR2_X1 U435 ( .A(KEYINPUT20), .B(KEYINPUT94), .ZN(n456) );
  NAND2_X1 U436 ( .A1(n662), .A2(G234), .ZN(n457) );
  XNOR2_X1 U437 ( .A(n471), .B(KEYINPUT17), .ZN(n470) );
  INV_X1 U438 ( .A(KEYINPUT18), .ZN(n471) );
  XNOR2_X1 U439 ( .A(n385), .B(n562), .ZN(n592) );
  XNOR2_X1 U440 ( .A(KEYINPUT22), .B(KEYINPUT66), .ZN(n562) );
  XNOR2_X1 U441 ( .A(n460), .B(n459), .ZN(n458) );
  XNOR2_X1 U442 ( .A(n567), .B(n565), .ZN(n460) );
  INV_X1 U443 ( .A(KEYINPUT28), .ZN(n436) );
  XNOR2_X1 U444 ( .A(n396), .B(n609), .ZN(n735) );
  NOR2_X1 U445 ( .A1(n713), .A2(n406), .ZN(n396) );
  XNOR2_X1 U446 ( .A(n557), .B(n560), .ZN(n467) );
  XNOR2_X1 U447 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n482) );
  XNOR2_X1 U448 ( .A(n387), .B(n512), .ZN(n753) );
  AND2_X1 U449 ( .A1(n637), .A2(KEYINPUT47), .ZN(n644) );
  NAND2_X1 U450 ( .A1(n704), .A2(n405), .ZN(n398) );
  INV_X1 U451 ( .A(n789), .ZN(n405) );
  INV_X1 U452 ( .A(G146), .ZN(n486) );
  AND2_X1 U453 ( .A1(n418), .A2(n417), .ZN(n416) );
  NOR2_X1 U454 ( .A1(n668), .A2(n480), .ZN(n478) );
  INV_X1 U455 ( .A(G237), .ZN(n523) );
  INV_X1 U456 ( .A(G902), .ZN(n524) );
  XNOR2_X1 U457 ( .A(KEYINPUT5), .B(G137), .ZN(n566) );
  XNOR2_X1 U458 ( .A(n360), .B(G113), .ZN(n564) );
  INV_X1 U459 ( .A(KEYINPUT10), .ZN(n489) );
  XOR2_X1 U460 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n546) );
  XNOR2_X1 U461 ( .A(KEYINPUT97), .B(KEYINPUT99), .ZN(n545) );
  XNOR2_X1 U462 ( .A(G143), .B(G131), .ZN(n539) );
  XOR2_X1 U463 ( .A(KEYINPUT101), .B(G140), .Z(n540) );
  XOR2_X1 U464 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n544) );
  XNOR2_X1 U465 ( .A(G134), .B(G131), .ZN(n511) );
  INV_X1 U466 ( .A(G101), .ZN(n507) );
  NAND2_X1 U467 ( .A1(n668), .A2(n480), .ZN(n479) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n528) );
  XNOR2_X1 U469 ( .A(n660), .B(KEYINPUT81), .ZN(n709) );
  NAND2_X1 U470 ( .A1(n724), .A2(n613), .ZN(n625) );
  INV_X1 U471 ( .A(KEYINPUT6), .ZN(n409) );
  XNOR2_X1 U472 ( .A(KEYINPUT3), .B(G119), .ZN(n442) );
  XNOR2_X1 U473 ( .A(n522), .B(G101), .ZN(n443) );
  INV_X1 U474 ( .A(KEYINPUT89), .ZN(n522) );
  XOR2_X1 U475 ( .A(G137), .B(G140), .Z(n508) );
  XOR2_X1 U476 ( .A(G107), .B(G104), .Z(n484) );
  XNOR2_X1 U477 ( .A(n384), .B(n472), .ZN(n469) );
  XNOR2_X1 U478 ( .A(n521), .B(n519), .ZN(n472) );
  XNOR2_X1 U479 ( .A(n520), .B(n470), .ZN(n384) );
  BUF_X1 U480 ( .A(n709), .Z(n776) );
  NAND2_X1 U481 ( .A1(n450), .A2(n439), .ZN(n622) );
  NOR2_X1 U482 ( .A1(n621), .A2(n406), .ZN(n439) );
  NOR2_X1 U483 ( .A1(n583), .A2(KEYINPUT34), .ZN(n413) );
  INV_X1 U484 ( .A(KEYINPUT0), .ZN(n468) );
  XNOR2_X1 U485 ( .A(n454), .B(n453), .ZN(n733) );
  INV_X1 U486 ( .A(KEYINPUT96), .ZN(n453) );
  NAND2_X1 U487 ( .A1(n455), .A2(n650), .ZN(n454) );
  AND2_X1 U488 ( .A1(n575), .A2(n440), .ZN(n455) );
  NOR2_X1 U489 ( .A1(G902), .A2(n760), .ZN(n502) );
  NOR2_X1 U490 ( .A1(n757), .A2(G902), .ZN(n386) );
  BUF_X1 U491 ( .A(n728), .Z(n440) );
  INV_X1 U492 ( .A(n594), .ZN(n724) );
  INV_X1 U493 ( .A(KEYINPUT42), .ZN(n394) );
  XNOR2_X1 U494 ( .A(n762), .B(n761), .ZN(n422) );
  XNOR2_X1 U495 ( .A(n758), .B(n757), .ZN(n383) );
  XNOR2_X1 U496 ( .A(n756), .B(n755), .ZN(n423) );
  INV_X1 U497 ( .A(KEYINPUT56), .ZN(n425) );
  XOR2_X1 U498 ( .A(n569), .B(G472), .Z(n366) );
  XNOR2_X1 U499 ( .A(KEYINPUT76), .B(n666), .ZN(n367) );
  XOR2_X1 U500 ( .A(KEYINPUT68), .B(KEYINPUT24), .Z(n370) );
  AND2_X1 U501 ( .A1(n404), .A2(n403), .ZN(n371) );
  AND2_X1 U502 ( .A1(n359), .A2(n463), .ZN(n372) );
  AND2_X1 U503 ( .A1(n506), .A2(n505), .ZN(n373) );
  NAND2_X1 U504 ( .A1(n527), .A2(G214), .ZN(n714) );
  XOR2_X1 U505 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n374) );
  XOR2_X1 U506 ( .A(KEYINPUT84), .B(KEYINPUT46), .Z(n375) );
  OR2_X1 U507 ( .A1(n662), .A2(n705), .ZN(n376) );
  AND2_X1 U508 ( .A1(n376), .A2(KEYINPUT65), .ZN(n378) );
  XNOR2_X1 U509 ( .A(KEYINPUT60), .B(KEYINPUT123), .ZN(n381) );
  XNOR2_X1 U510 ( .A(KEYINPUT114), .B(KEYINPUT63), .ZN(n382) );
  AND2_X1 U511 ( .A1(n675), .A2(G953), .ZN(n763) );
  INV_X1 U512 ( .A(n763), .ZN(n429) );
  XNOR2_X1 U513 ( .A(n449), .B(n507), .ZN(n448) );
  XNOR2_X1 U514 ( .A(n437), .B(n436), .ZN(n615) );
  XNOR2_X1 U515 ( .A(n431), .B(KEYINPUT83), .ZN(n667) );
  NAND2_X1 U516 ( .A1(n421), .A2(n362), .ZN(n420) );
  XNOR2_X1 U517 ( .A(n664), .B(n603), .ZN(n605) );
  NAND2_X1 U518 ( .A1(n601), .A2(n602), .ZN(n664) );
  NOR2_X1 U519 ( .A1(n383), .A2(n763), .ZN(G63) );
  NAND2_X1 U520 ( .A1(n561), .A2(n577), .ZN(n385) );
  INV_X1 U521 ( .A(n568), .ZN(n387) );
  XNOR2_X1 U522 ( .A(n388), .B(n648), .ZN(n656) );
  NAND2_X1 U523 ( .A1(n397), .A2(n399), .ZN(n388) );
  AND2_X2 U524 ( .A1(n572), .A2(n584), .ZN(n698) );
  AND2_X2 U525 ( .A1(n391), .A2(n389), .ZN(n421) );
  NAND2_X1 U526 ( .A1(n390), .A2(n598), .ZN(n417) );
  INV_X1 U527 ( .A(n391), .ZN(n390) );
  XNOR2_X1 U528 ( .A(n391), .B(G119), .ZN(G21) );
  XNOR2_X2 U529 ( .A(n597), .B(n374), .ZN(n391) );
  NAND2_X1 U530 ( .A1(n393), .A2(n574), .ZN(n465) );
  NAND2_X1 U531 ( .A1(n393), .A2(n714), .ZN(n713) );
  NOR2_X1 U532 ( .A1(n716), .A2(n393), .ZN(n717) );
  XNOR2_X2 U533 ( .A(n466), .B(KEYINPUT104), .ZN(n393) );
  XNOR2_X2 U534 ( .A(n395), .B(n394), .ZN(n792) );
  NAND2_X1 U535 ( .A1(n635), .A2(n735), .ZN(n395) );
  NAND2_X1 U536 ( .A1(n371), .A2(n400), .ZN(n399) );
  NAND2_X1 U537 ( .A1(n402), .A2(n401), .ZN(n400) );
  INV_X1 U538 ( .A(n682), .ZN(n401) );
  NOR2_X1 U539 ( .A1(n792), .A2(n375), .ZN(n402) );
  NAND2_X1 U540 ( .A1(n792), .A2(n375), .ZN(n403) );
  NAND2_X1 U541 ( .A1(n682), .A2(n375), .ZN(n404) );
  NOR2_X1 U542 ( .A1(n717), .A2(n406), .ZN(n718) );
  INV_X1 U543 ( .A(n407), .ZN(n708) );
  NAND2_X1 U544 ( .A1(n407), .A2(KEYINPUT65), .ZN(n474) );
  NAND2_X1 U545 ( .A1(n728), .A2(n714), .ZN(n619) );
  NOR2_X1 U546 ( .A1(n625), .A2(n408), .ZN(n437) );
  INV_X1 U547 ( .A(n728), .ZN(n408) );
  XNOR2_X2 U548 ( .A(n728), .B(n409), .ZN(n627) );
  XNOR2_X2 U549 ( .A(n570), .B(n366), .ZN(n728) );
  AND2_X1 U550 ( .A1(n411), .A2(n645), .ZN(n410) );
  NAND2_X1 U551 ( .A1(n583), .A2(KEYINPUT34), .ZN(n411) );
  NAND2_X1 U552 ( .A1(n414), .A2(n413), .ZN(n412) );
  INV_X1 U553 ( .A(n712), .ZN(n414) );
  NAND2_X1 U554 ( .A1(n712), .A2(KEYINPUT34), .ZN(n415) );
  NAND2_X1 U555 ( .A1(n419), .A2(n416), .ZN(n601) );
  NAND2_X1 U556 ( .A1(n692), .A2(n598), .ZN(n418) );
  NOR2_X1 U557 ( .A1(n422), .A2(n763), .ZN(G66) );
  NAND2_X1 U558 ( .A1(n589), .A2(n590), .ZN(n591) );
  NOR2_X1 U559 ( .A1(n423), .A2(n763), .ZN(G54) );
  XNOR2_X1 U560 ( .A(n424), .B(n381), .ZN(G60) );
  NAND2_X1 U561 ( .A1(n430), .A2(n429), .ZN(n424) );
  XNOR2_X1 U562 ( .A(n426), .B(n425), .ZN(G51) );
  NAND2_X1 U563 ( .A1(n427), .A2(n429), .ZN(n426) );
  XNOR2_X1 U564 ( .A(n679), .B(n380), .ZN(n427) );
  NAND2_X1 U565 ( .A1(n656), .A2(n655), .ZN(n431) );
  XNOR2_X1 U566 ( .A(n674), .B(n379), .ZN(n430) );
  INV_X1 U567 ( .A(n771), .ZN(n432) );
  XNOR2_X1 U568 ( .A(n433), .B(n382), .ZN(G57) );
  NAND2_X1 U569 ( .A1(n434), .A2(n429), .ZN(n433) );
  XNOR2_X1 U570 ( .A(n685), .B(n377), .ZN(n434) );
  NAND2_X1 U571 ( .A1(n477), .A2(n378), .ZN(n435) );
  XNOR2_X1 U572 ( .A(n447), .B(n521), .ZN(n510) );
  XNOR2_X2 U573 ( .A(n559), .B(KEYINPUT16), .ZN(n446) );
  XNOR2_X2 U574 ( .A(n438), .B(G107), .ZN(n559) );
  NAND2_X1 U575 ( .A1(n681), .A2(n667), .ZN(n660) );
  NOR2_X1 U576 ( .A1(G902), .A2(n671), .ZN(n552) );
  XNOR2_X1 U577 ( .A(n465), .B(KEYINPUT105), .ZN(n561) );
  NOR2_X2 U578 ( .A1(n585), .A2(n584), .ZN(n466) );
  XNOR2_X1 U579 ( .A(n498), .B(n777), .ZN(n760) );
  NAND2_X1 U580 ( .A1(n618), .A2(n617), .ZN(n621) );
  XNOR2_X2 U581 ( .A(n444), .B(n441), .ZN(n765) );
  XNOR2_X2 U582 ( .A(n446), .B(n537), .ZN(n444) );
  XNOR2_X2 U583 ( .A(n445), .B(G122), .ZN(n537) );
  XNOR2_X2 U584 ( .A(G113), .B(G104), .ZN(n445) );
  XNOR2_X2 U585 ( .A(G110), .B(KEYINPUT88), .ZN(n764) );
  XNOR2_X1 U586 ( .A(n448), .B(n373), .ZN(n447) );
  NAND2_X1 U587 ( .A1(n516), .A2(G227), .ZN(n449) );
  INV_X1 U588 ( .A(n620), .ZN(n450) );
  NOR2_X1 U589 ( .A1(n620), .A2(n621), .ZN(n451) );
  NAND2_X1 U590 ( .A1(n451), .A2(n646), .ZN(n647) );
  NAND2_X1 U591 ( .A1(n634), .A2(n533), .ZN(n534) );
  XNOR2_X2 U592 ( .A(n526), .B(n525), .ZN(n608) );
  NAND2_X1 U593 ( .A1(n733), .A2(n577), .ZN(n576) );
  XNOR2_X1 U594 ( .A(n568), .B(n458), .ZN(n684) );
  XNOR2_X1 U595 ( .A(n564), .B(n566), .ZN(n459) );
  INV_X1 U596 ( .A(n669), .ZN(n462) );
  NAND2_X1 U597 ( .A1(n669), .A2(n480), .ZN(n464) );
  XNOR2_X2 U598 ( .A(n534), .B(n468), .ZN(n577) );
  NAND2_X2 U599 ( .A1(n473), .A2(n475), .ZN(n752) );
  NAND2_X1 U600 ( .A1(n372), .A2(n476), .ZN(n475) );
  NAND2_X1 U601 ( .A1(n477), .A2(n376), .ZN(n476) );
  OR2_X1 U602 ( .A1(n742), .A2(G953), .ZN(n483) );
  INV_X1 U603 ( .A(n663), .ZN(n603) );
  INV_X1 U604 ( .A(KEYINPUT48), .ZN(n648) );
  INV_X1 U605 ( .A(KEYINPUT80), .ZN(n606) );
  XNOR2_X1 U606 ( .A(n599), .B(KEYINPUT86), .ZN(n598) );
  BUF_X1 U607 ( .A(n735), .Z(n743) );
  XNOR2_X1 U608 ( .A(n538), .B(n537), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n490), .B(n358), .ZN(n493) );
  XNOR2_X1 U610 ( .A(n493), .B(n492), .ZN(n497) );
  INV_X1 U611 ( .A(n776), .ZN(n779) );
  BUF_X1 U612 ( .A(n671), .Z(n673) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n512) );
  INV_X1 U614 ( .A(G125), .ZN(n485) );
  NAND2_X1 U615 ( .A1(G146), .A2(n485), .ZN(n488) );
  NAND2_X1 U616 ( .A1(n486), .A2(G125), .ZN(n487) );
  NAND2_X2 U617 ( .A1(n488), .A2(n487), .ZN(n518) );
  XNOR2_X2 U618 ( .A(n518), .B(n489), .ZN(n538) );
  XOR2_X1 U619 ( .A(n508), .B(n538), .Z(n777) );
  XOR2_X1 U620 ( .A(KEYINPUT93), .B(G110), .Z(n490) );
  XNOR2_X1 U621 ( .A(KEYINPUT92), .B(KEYINPUT23), .ZN(n491) );
  XNOR2_X1 U622 ( .A(n370), .B(n491), .ZN(n492) );
  NAND2_X1 U623 ( .A1(n516), .A2(G234), .ZN(n495) );
  XNOR2_X1 U624 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n494) );
  XNOR2_X1 U625 ( .A(n495), .B(n494), .ZN(n556) );
  NAND2_X1 U626 ( .A1(G221), .A2(n556), .ZN(n496) );
  XNOR2_X1 U627 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U628 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n500) );
  NAND2_X1 U629 ( .A1(G217), .A2(n535), .ZN(n499) );
  XNOR2_X1 U630 ( .A(n500), .B(n499), .ZN(n501) );
  INV_X1 U631 ( .A(KEYINPUT73), .ZN(n503) );
  NAND2_X1 U632 ( .A1(KEYINPUT74), .A2(n503), .ZN(n506) );
  INV_X1 U633 ( .A(KEYINPUT74), .ZN(n504) );
  NAND2_X1 U634 ( .A1(n504), .A2(KEYINPUT73), .ZN(n505) );
  XNOR2_X1 U635 ( .A(n508), .B(n484), .ZN(n509) );
  XNOR2_X2 U636 ( .A(G143), .B(G128), .ZN(n554) );
  NAND2_X1 U637 ( .A1(n753), .A2(n524), .ZN(n514) );
  INV_X1 U638 ( .A(G469), .ZN(n513) );
  XNOR2_X2 U639 ( .A(n514), .B(n513), .ZN(n614) );
  INV_X1 U640 ( .A(KEYINPUT1), .ZN(n515) );
  XNOR2_X2 U641 ( .A(n614), .B(n515), .ZN(n650) );
  INV_X1 U642 ( .A(n650), .ZN(n722) );
  NAND2_X1 U643 ( .A1(n516), .A2(G224), .ZN(n517) );
  XNOR2_X1 U644 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U645 ( .A1(n676), .A2(n662), .ZN(n526) );
  NAND2_X1 U646 ( .A1(n524), .A2(n523), .ZN(n527) );
  AND2_X1 U647 ( .A1(n527), .A2(G210), .ZN(n525) );
  XNOR2_X1 U648 ( .A(n528), .B(KEYINPUT90), .ZN(n529) );
  XNOR2_X1 U649 ( .A(KEYINPUT14), .B(n529), .ZN(n530) );
  NAND2_X1 U650 ( .A1(G952), .A2(n530), .ZN(n742) );
  NAND2_X1 U651 ( .A1(n530), .A2(G902), .ZN(n531) );
  XNOR2_X1 U652 ( .A(n531), .B(KEYINPUT91), .ZN(n610) );
  NOR2_X1 U653 ( .A1(G898), .A2(n516), .ZN(n767) );
  NAND2_X1 U654 ( .A1(n610), .A2(n767), .ZN(n532) );
  NAND2_X1 U655 ( .A1(n483), .A2(n532), .ZN(n533) );
  NAND2_X1 U656 ( .A1(n535), .A2(G221), .ZN(n536) );
  XNOR2_X1 U657 ( .A(n536), .B(KEYINPUT21), .ZN(n725) );
  INV_X1 U658 ( .A(n725), .ZN(n574) );
  XNOR2_X1 U659 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U660 ( .A(n542), .B(n541), .ZN(n550) );
  NOR2_X1 U661 ( .A1(G953), .A2(G237), .ZN(n563) );
  NAND2_X1 U662 ( .A1(G214), .A2(n563), .ZN(n543) );
  XNOR2_X1 U663 ( .A(n544), .B(n543), .ZN(n548) );
  XNOR2_X1 U664 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U665 ( .A(n548), .B(n547), .Z(n549) );
  XNOR2_X1 U666 ( .A(n550), .B(n549), .ZN(n671) );
  XNOR2_X1 U667 ( .A(KEYINPUT13), .B(G475), .ZN(n551) );
  XNOR2_X2 U668 ( .A(n552), .B(n551), .ZN(n584) );
  XOR2_X1 U669 ( .A(G122), .B(KEYINPUT102), .Z(n553) );
  XNOR2_X1 U670 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U671 ( .A(n555), .B(n482), .ZN(n558) );
  NAND2_X1 U672 ( .A1(G217), .A2(n556), .ZN(n557) );
  XNOR2_X1 U673 ( .A(G134), .B(n559), .ZN(n560) );
  INV_X1 U674 ( .A(n572), .ZN(n585) );
  NAND2_X1 U675 ( .A1(n563), .A2(G210), .ZN(n565) );
  INV_X1 U676 ( .A(KEYINPUT70), .ZN(n569) );
  NOR2_X2 U677 ( .A1(n592), .A2(n627), .ZN(n596) );
  NAND2_X1 U678 ( .A1(n722), .A2(n596), .ZN(n571) );
  NOR2_X1 U679 ( .A1(n724), .A2(n571), .ZN(n686) );
  OR2_X1 U680 ( .A1(n584), .A2(n572), .ZN(n658) );
  INV_X1 U681 ( .A(n658), .ZN(n700) );
  NOR2_X1 U682 ( .A1(n700), .A2(n698), .ZN(n573) );
  XNOR2_X1 U683 ( .A(KEYINPUT103), .B(n573), .ZN(n715) );
  INV_X1 U684 ( .A(n715), .ZN(n638) );
  INV_X1 U685 ( .A(n721), .ZN(n575) );
  XNOR2_X1 U686 ( .A(n576), .B(KEYINPUT31), .ZN(n701) );
  INV_X1 U687 ( .A(n577), .ZN(n583) );
  NOR2_X1 U688 ( .A1(n721), .A2(n440), .ZN(n578) );
  INV_X1 U689 ( .A(n614), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n578), .A2(n617), .ZN(n579) );
  NOR2_X1 U691 ( .A1(n583), .A2(n579), .ZN(n688) );
  NOR2_X1 U692 ( .A1(n701), .A2(n688), .ZN(n580) );
  NOR2_X1 U693 ( .A1(n638), .A2(n580), .ZN(n581) );
  NOR2_X1 U694 ( .A1(n686), .A2(n581), .ZN(n590) );
  NAND2_X1 U695 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U696 ( .A(n586), .B(KEYINPUT108), .Z(n645) );
  XNOR2_X1 U697 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n587) );
  XNOR2_X2 U698 ( .A(n588), .B(n587), .ZN(n791) );
  NAND2_X1 U699 ( .A1(n791), .A2(KEYINPUT44), .ZN(n589) );
  XNOR2_X1 U700 ( .A(n591), .B(KEYINPUT85), .ZN(n602) );
  NOR2_X1 U701 ( .A1(n594), .A2(n440), .ZN(n593) );
  NOR2_X1 U702 ( .A1(n722), .A2(n594), .ZN(n595) );
  NAND2_X1 U703 ( .A1(n596), .A2(n595), .ZN(n597) );
  INV_X1 U704 ( .A(KEYINPUT44), .ZN(n599) );
  NAND2_X1 U705 ( .A1(n599), .A2(n791), .ZN(n600) );
  XOR2_X1 U706 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n663) );
  INV_X1 U707 ( .A(n662), .ZN(n604) );
  NAND2_X1 U708 ( .A1(n605), .A2(n604), .ZN(n607) );
  XNOR2_X1 U709 ( .A(n607), .B(n606), .ZN(n661) );
  XNOR2_X1 U710 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n609) );
  NAND2_X1 U711 ( .A1(G953), .A2(n610), .ZN(n611) );
  OR2_X1 U712 ( .A1(n611), .A2(G900), .ZN(n612) );
  AND2_X1 U713 ( .A1(n483), .A2(n612), .ZN(n616) );
  NOR2_X1 U714 ( .A1(n616), .A2(n725), .ZN(n613) );
  NOR2_X1 U715 ( .A1(n615), .A2(n614), .ZN(n635) );
  XNOR2_X1 U716 ( .A(n619), .B(KEYINPUT30), .ZN(n620) );
  NAND2_X1 U717 ( .A1(n657), .A2(n698), .ZN(n624) );
  XOR2_X1 U718 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n623) );
  INV_X1 U719 ( .A(n698), .ZN(n626) );
  NOR2_X1 U720 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U721 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U722 ( .A(n629), .B(KEYINPUT109), .ZN(n630) );
  NAND2_X1 U723 ( .A1(n630), .A2(n714), .ZN(n649) );
  INV_X1 U724 ( .A(n652), .ZN(n631) );
  NOR2_X1 U725 ( .A1(n649), .A2(n631), .ZN(n632) );
  XNOR2_X1 U726 ( .A(n632), .B(KEYINPUT36), .ZN(n633) );
  NAND2_X1 U727 ( .A1(n633), .A2(n650), .ZN(n704) );
  NAND2_X1 U728 ( .A1(n635), .A2(n634), .ZN(n642) );
  NOR2_X1 U729 ( .A1(KEYINPUT71), .A2(n638), .ZN(n636) );
  NAND2_X1 U730 ( .A1(n695), .A2(n636), .ZN(n637) );
  XNOR2_X1 U731 ( .A(n638), .B(KEYINPUT71), .ZN(n640) );
  INV_X1 U732 ( .A(KEYINPUT47), .ZN(n639) );
  NAND2_X1 U733 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U734 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U735 ( .A1(n652), .A2(n645), .ZN(n646) );
  XNOR2_X1 U736 ( .A(n647), .B(KEYINPUT111), .ZN(n789) );
  NOR2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U738 ( .A(n651), .B(KEYINPUT43), .ZN(n653) );
  NOR2_X1 U739 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U740 ( .A(n654), .B(KEYINPUT110), .ZN(n788) );
  INV_X1 U741 ( .A(n788), .ZN(n655) );
  INV_X1 U742 ( .A(n657), .ZN(n659) );
  OR2_X1 U743 ( .A1(n659), .A2(n658), .ZN(n681) );
  INV_X1 U744 ( .A(KEYINPUT2), .ZN(n705) );
  XNOR2_X1 U745 ( .A(n664), .B(n663), .ZN(n771) );
  INV_X1 U746 ( .A(n681), .ZN(n665) );
  NOR2_X1 U747 ( .A1(n665), .A2(n705), .ZN(n666) );
  INV_X1 U748 ( .A(n667), .ZN(n668) );
  INV_X1 U749 ( .A(KEYINPUT65), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n752), .A2(G475), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n672) );
  INV_X1 U752 ( .A(G952), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n752), .A2(G210), .ZN(n679) );
  XOR2_X1 U754 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n678) );
  XNOR2_X1 U755 ( .A(n676), .B(KEYINPUT77), .ZN(n677) );
  XOR2_X1 U756 ( .A(G134), .B(KEYINPUT117), .Z(n680) );
  XNOR2_X1 U757 ( .A(n681), .B(n680), .ZN(G36) );
  XOR2_X1 U758 ( .A(n361), .B(G131), .Z(G33) );
  NAND2_X1 U759 ( .A1(n752), .A2(G472), .ZN(n685) );
  XOR2_X1 U760 ( .A(KEYINPUT87), .B(KEYINPUT62), .Z(n683) );
  XOR2_X1 U761 ( .A(G101), .B(n686), .Z(G3) );
  NAND2_X1 U762 ( .A1(n688), .A2(n698), .ZN(n687) );
  XNOR2_X1 U763 ( .A(n687), .B(G104), .ZN(G6) );
  XOR2_X1 U764 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n690) );
  NAND2_X1 U765 ( .A1(n688), .A2(n700), .ZN(n689) );
  XNOR2_X1 U766 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U767 ( .A(G107), .B(n691), .ZN(G9) );
  XOR2_X1 U768 ( .A(n692), .B(G110), .Z(G12) );
  XOR2_X1 U769 ( .A(G128), .B(KEYINPUT29), .Z(n694) );
  NAND2_X1 U770 ( .A1(n695), .A2(n700), .ZN(n693) );
  XNOR2_X1 U771 ( .A(n694), .B(n693), .ZN(G30) );
  NAND2_X1 U772 ( .A1(n695), .A2(n698), .ZN(n696) );
  XNOR2_X1 U773 ( .A(n696), .B(KEYINPUT116), .ZN(n697) );
  XNOR2_X1 U774 ( .A(G146), .B(n697), .ZN(G48) );
  NAND2_X1 U775 ( .A1(n701), .A2(n698), .ZN(n699) );
  XNOR2_X1 U776 ( .A(n699), .B(G113), .ZN(G15) );
  NAND2_X1 U777 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U778 ( .A(n702), .B(n360), .ZN(G18) );
  XOR2_X1 U779 ( .A(G125), .B(KEYINPUT37), .Z(n703) );
  XNOR2_X1 U780 ( .A(n704), .B(n703), .ZN(G27) );
  NAND2_X1 U781 ( .A1(n771), .A2(n705), .ZN(n706) );
  XNOR2_X1 U782 ( .A(KEYINPUT78), .B(n706), .ZN(n707) );
  NAND2_X1 U783 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U784 ( .A1(n776), .A2(KEYINPUT2), .ZN(n710) );
  NOR2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n749) );
  INV_X1 U786 ( .A(n713), .ZN(n719) );
  AND2_X1 U787 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U788 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U789 ( .A1(n357), .A2(n720), .ZN(n739) );
  NAND2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U791 ( .A(KEYINPUT50), .B(n723), .ZN(n731) );
  XOR2_X1 U792 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n727) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U794 ( .A(n727), .B(n726), .ZN(n729) );
  NOR2_X1 U795 ( .A1(n729), .A2(n440), .ZN(n730) );
  AND2_X1 U796 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U797 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U798 ( .A(KEYINPUT51), .B(n734), .ZN(n736) );
  NAND2_X1 U799 ( .A1(n736), .A2(n743), .ZN(n737) );
  XOR2_X1 U800 ( .A(KEYINPUT120), .B(n737), .Z(n738) );
  NOR2_X1 U801 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U802 ( .A(n740), .B(KEYINPUT52), .ZN(n741) );
  NOR2_X1 U803 ( .A1(n742), .A2(n741), .ZN(n746) );
  INV_X1 U804 ( .A(n743), .ZN(n744) );
  NOR2_X1 U805 ( .A1(n357), .A2(n744), .ZN(n745) );
  NOR2_X1 U806 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U807 ( .A(n747), .B(KEYINPUT121), .ZN(n748) );
  NOR2_X1 U808 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U809 ( .A1(n516), .A2(n750), .ZN(n751) );
  XOR2_X1 U810 ( .A(KEYINPUT53), .B(n751), .Z(G75) );
  NAND2_X1 U811 ( .A1(n759), .A2(G469), .ZN(n756) );
  XOR2_X1 U812 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n754) );
  XOR2_X1 U813 ( .A(n754), .B(n753), .Z(n755) );
  NAND2_X1 U814 ( .A1(n759), .A2(G478), .ZN(n758) );
  NAND2_X1 U815 ( .A1(n759), .A2(G217), .ZN(n762) );
  XNOR2_X1 U816 ( .A(n760), .B(KEYINPUT124), .ZN(n761) );
  XNOR2_X1 U817 ( .A(n765), .B(n764), .ZN(n766) );
  NOR2_X1 U818 ( .A1(n767), .A2(n766), .ZN(n775) );
  XOR2_X1 U819 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n769) );
  NAND2_X1 U820 ( .A1(G224), .A2(G953), .ZN(n768) );
  XNOR2_X1 U821 ( .A(n769), .B(n768), .ZN(n770) );
  NAND2_X1 U822 ( .A1(n770), .A2(G898), .ZN(n773) );
  OR2_X1 U823 ( .A1(n771), .A2(G953), .ZN(n772) );
  NAND2_X1 U824 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U825 ( .A(n775), .B(n774), .ZN(G69) );
  XOR2_X1 U826 ( .A(n778), .B(n777), .Z(n781) );
  XNOR2_X1 U827 ( .A(n779), .B(n781), .ZN(n780) );
  NAND2_X1 U828 ( .A1(n780), .A2(n516), .ZN(n785) );
  XNOR2_X1 U829 ( .A(n781), .B(G227), .ZN(n782) );
  NAND2_X1 U830 ( .A1(n782), .A2(G900), .ZN(n783) );
  NAND2_X1 U831 ( .A1(n783), .A2(G953), .ZN(n784) );
  NAND2_X1 U832 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U833 ( .A(KEYINPUT126), .B(n786), .ZN(G72) );
  XOR2_X1 U834 ( .A(G140), .B(KEYINPUT118), .Z(n787) );
  XNOR2_X1 U835 ( .A(n788), .B(n787), .ZN(G42) );
  XNOR2_X1 U836 ( .A(G143), .B(n789), .ZN(n790) );
  XNOR2_X1 U837 ( .A(n790), .B(KEYINPUT115), .ZN(G45) );
  XOR2_X1 U838 ( .A(n791), .B(G122), .Z(G24) );
  XOR2_X1 U839 ( .A(n792), .B(G137), .Z(G39) );
endmodule

