//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(G101), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT4), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT4), .ZN(new_n199));
  AOI21_X1  g013(.A(G101), .B1(new_n190), .B2(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(new_n200), .A3(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n191), .A2(new_n200), .A3(new_n194), .A4(KEYINPUT80), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n199), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n198), .B1(new_n205), .B2(new_n197), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G116), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT2), .B(G113), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT68), .ZN(new_n215));
  INV_X1    g029(.A(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT2), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G116), .B(G119), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n207), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n215), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n222), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n224), .B1(new_n223), .B2(new_n207), .ZN(new_n228));
  AOI211_X1 g042(.A(KEYINPUT67), .B(KEYINPUT68), .C1(new_n220), .C2(new_n221), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n206), .A2(new_n226), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G101), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n193), .A2(G104), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n195), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n203), .B2(new_n204), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n209), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n216), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n221), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n240), .A2(new_n242), .B1(new_n221), .B2(new_n220), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n235), .A2(new_n243), .A3(KEYINPUT85), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT85), .B1(new_n235), .B2(new_n243), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n187), .B(new_n189), .C1(new_n231), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT6), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n203), .A2(new_n204), .ZN(new_n250));
  INV_X1    g064(.A(new_n234), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n242), .ZN(new_n253));
  OAI21_X1  g067(.A(G113), .B1(new_n241), .B2(new_n209), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n223), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n249), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n235), .A2(new_n243), .A3(KEYINPUT85), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n206), .A2(new_n226), .A3(new_n230), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n188), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n187), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n248), .A2(new_n261), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n228), .A2(new_n229), .A3(new_n227), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n222), .B1(new_n215), .B2(new_n225), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n265), .A2(new_n206), .B1(new_n256), .B2(new_n257), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT87), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n188), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n258), .A2(new_n188), .A3(new_n259), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT87), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n260), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT88), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n260), .A2(KEYINPUT88), .A3(new_n272), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n262), .A2(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G128), .ZN(new_n278));
  INV_X1    g092(.A(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT64), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G146), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n282), .A3(G143), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n278), .B1(new_n283), .B2(KEYINPUT1), .ZN(new_n284));
  INV_X1    g098(.A(G143), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(G146), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n282), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n285), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT65), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n290));
  INV_X1    g104(.A(new_n286), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT64), .B(G146), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(G143), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n292), .B2(G143), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n290), .B(new_n293), .C1(new_n295), .C2(new_n278), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G125), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n279), .A2(G143), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n283), .A2(new_n294), .A3(G128), .A4(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT89), .ZN(new_n303));
  AND2_X1   g117(.A1(KEYINPUT0), .A2(G128), .ZN(new_n304));
  NOR2_X1   g118(.A1(KEYINPUT0), .A2(G128), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n299), .B1(new_n292), .B2(G143), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n293), .A2(new_n306), .B1(new_n307), .B2(new_n304), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n303), .B1(new_n308), .B2(new_n298), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n293), .A2(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n304), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n298), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT89), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G224), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(G953), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n314), .B(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT7), .B1(new_n315), .B2(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n301), .ZN(new_n319));
  AOI211_X1 g133(.A(G125), .B(new_n319), .C1(new_n289), .C2(new_n296), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n320), .B2(new_n312), .ZN(new_n321));
  INV_X1    g135(.A(new_n318), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n302), .A2(new_n309), .A3(new_n313), .A4(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n221), .A2(KEYINPUT5), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n223), .B1(new_n324), .B2(new_n254), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n235), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n188), .B(KEYINPUT8), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(new_n235), .C2(new_n255), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n321), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n268), .B2(new_n270), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT90), .B1(new_n330), .B2(G902), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n319), .B1(new_n289), .B2(new_n296), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n312), .B1(new_n332), .B2(new_n298), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n328), .B1(new_n333), .B2(new_n322), .ZN(new_n334));
  AND4_X1   g148(.A1(new_n302), .A2(new_n309), .A3(new_n313), .A4(new_n322), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n267), .B1(new_n266), .B2(new_n188), .ZN(new_n337));
  AND4_X1   g151(.A1(new_n267), .A2(new_n258), .A3(new_n188), .A4(new_n259), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT90), .ZN(new_n340));
  INV_X1    g154(.A(G902), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n277), .A2(new_n317), .B1(new_n331), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G210), .B1(G237), .B2(G902), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT91), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n331), .A2(new_n342), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT86), .B1(new_n266), .B2(new_n188), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n271), .A2(KEYINPUT6), .A3(new_n348), .A4(new_n247), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n275), .A2(new_n276), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n317), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT91), .ZN(new_n353));
  INV_X1    g167(.A(new_n344), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n345), .A2(new_n346), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G237), .A2(G953), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n357), .A2(G143), .A3(G214), .ZN(new_n358));
  AOI21_X1  g172(.A(G143), .B1(new_n357), .B2(G214), .ZN(new_n359));
  OAI211_X1 g173(.A(KEYINPUT17), .B(G131), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT92), .ZN(new_n361));
  INV_X1    g175(.A(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G125), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n298), .A2(G140), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT16), .ZN(new_n365));
  OR3_X1    g179(.A1(new_n298), .A2(KEYINPUT16), .A3(G140), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(G146), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT73), .A4(G146), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n366), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n279), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT93), .B1(new_n361), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n358), .A2(new_n359), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G131), .ZN(new_n377));
  INV_X1    g191(.A(G131), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n380), .A2(KEYINPUT17), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n360), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n373), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT93), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n374), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(new_n190), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n376), .A2(KEYINPUT18), .A3(G131), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n363), .A2(new_n364), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n292), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n279), .B2(new_n391), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT18), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n375), .B1(new_n394), .B2(new_n378), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n391), .B(KEYINPUT19), .Z(new_n398));
  OAI211_X1 g212(.A(new_n380), .B(new_n367), .C1(new_n398), .C2(new_n287), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n396), .ZN(new_n400));
  INV_X1    g214(.A(new_n389), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(G475), .A2(G902), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT20), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  INV_X1    g222(.A(new_n397), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n389), .B1(new_n387), .B2(new_n396), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n341), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n406), .A2(new_n408), .B1(G475), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(G116), .B(G122), .Z(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(G107), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n285), .A2(G128), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT96), .ZN(new_n416));
  INV_X1    g230(.A(G134), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n285), .A2(G128), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT94), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n422));
  OR2_X1    g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n422), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n416), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n421), .B1(new_n425), .B2(G134), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n210), .A2(G122), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n193), .B1(new_n427), .B2(KEYINPUT14), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(new_n413), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n416), .A2(new_n419), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G134), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n429), .B1(new_n431), .B2(new_n420), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT9), .B(G234), .ZN(new_n434));
  INV_X1    g248(.A(G217), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(G953), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n436), .B1(new_n426), .B2(new_n432), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G902), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n412), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G952), .ZN(new_n446));
  AOI211_X1 g260(.A(G953), .B(new_n446), .C1(G234), .C2(G237), .ZN(new_n447));
  INV_X1    g261(.A(G953), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n341), .B(new_n448), .C1(G234), .C2(G237), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(G898), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G214), .B1(G237), .B2(G902), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n356), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n435), .B1(G234), .B2(new_n341), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT23), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n208), .B2(G128), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n208), .A2(G128), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n278), .A2(KEYINPUT23), .A3(G119), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT24), .B(G110), .Z(new_n462));
  XNOR2_X1  g276(.A(G119), .B(G128), .ZN(new_n463));
  OAI22_X1  g277(.A1(new_n461), .A2(G110), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n392), .A3(new_n367), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT22), .B(G137), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n448), .A2(G221), .A3(G234), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n466), .B(new_n467), .Z(new_n468));
  AND2_X1   g282(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n461), .A2(G110), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT72), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n461), .A2(new_n472), .A3(G110), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n474), .A2(new_n373), .A3(KEYINPUT74), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT74), .B1(new_n474), .B2(new_n373), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n465), .B(new_n468), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT76), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n474), .A2(new_n373), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT74), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n474), .A2(KEYINPUT74), .A3(new_n373), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n484), .A2(KEYINPUT76), .A3(new_n465), .A4(new_n468), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT75), .B(new_n465), .C1(new_n475), .C2(new_n476), .ZN(new_n490));
  INV_X1    g304(.A(new_n468), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n493), .B2(KEYINPUT77), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n486), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n493), .A2(KEYINPUT77), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n456), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n496), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n486), .A2(new_n492), .A3(new_n498), .A4(new_n494), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n486), .A2(new_n492), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n455), .A2(G902), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n497), .A2(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G221), .B1(new_n434), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT11), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n417), .B2(G137), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n417), .A2(G137), .ZN(new_n508));
  INV_X1    g322(.A(G137), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT11), .A3(G134), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G131), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n507), .A2(new_n510), .A3(new_n378), .A4(new_n508), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(KEYINPUT69), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n278), .B1(new_n291), .B2(KEYINPUT1), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n301), .B1(new_n307), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n235), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT10), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n206), .A2(new_n308), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT81), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n297), .A2(new_n301), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n235), .A2(KEYINPUT10), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n332), .A2(KEYINPUT81), .A3(new_n526), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n518), .B(new_n523), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n332), .A2(KEYINPUT82), .A3(new_n252), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT82), .B1(new_n332), .B2(new_n252), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n521), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n518), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT12), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n514), .A2(KEYINPUT12), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT82), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n525), .B2(new_n235), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n332), .A2(KEYINPUT82), .A3(new_n252), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n540), .B2(new_n521), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n530), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n448), .A2(G227), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT78), .ZN(new_n544));
  XOR2_X1   g358(.A(G110), .B(G140), .Z(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n546), .B(KEYINPUT79), .Z(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT83), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT83), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n551), .B(new_n523), .C1(new_n528), .C2(new_n529), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n534), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n530), .A2(new_n546), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n542), .A2(new_n548), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G469), .B1(new_n556), .B2(G902), .ZN(new_n557));
  INV_X1    g371(.A(G469), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n546), .B1(new_n553), .B2(new_n530), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n538), .A2(new_n539), .B1(new_n235), .B2(new_n520), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(new_n518), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n533), .A2(KEYINPUT12), .A3(new_n514), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n554), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n558), .B(new_n341), .C1(new_n559), .C2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n505), .B1(new_n557), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n357), .A2(G210), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n567), .B(KEYINPUT27), .Z(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT26), .B(G101), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n568), .B(new_n569), .Z(new_n570));
  NAND2_X1  g384(.A1(new_n230), .A2(new_n226), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n516), .A2(new_n308), .A3(new_n517), .ZN(new_n572));
  INV_X1    g386(.A(new_n508), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n417), .A2(G137), .ZN(new_n574));
  OAI21_X1  g388(.A(G131), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n513), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n571), .B(new_n572), .C1(new_n332), .C2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT28), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n577), .A2(KEYINPUT71), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT71), .B1(new_n577), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n310), .A2(new_n311), .ZN(new_n582));
  INV_X1    g396(.A(new_n514), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n576), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n525), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n577), .B1(new_n586), .B2(new_n571), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT28), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n570), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n525), .A2(new_n585), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT70), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT30), .A4(new_n572), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n572), .B(KEYINPUT30), .C1(new_n332), .C2(new_n576), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT70), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT66), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n586), .A2(new_n597), .A3(KEYINPUT30), .ZN(new_n598));
  OAI22_X1  g412(.A1(new_n332), .A2(new_n576), .B1(new_n582), .B2(new_n583), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT30), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT66), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n596), .B(new_n265), .C1(new_n598), .C2(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n577), .A2(new_n570), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n602), .A2(KEYINPUT31), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT31), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n590), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(G472), .A2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT32), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n572), .B1(new_n332), .B2(new_n576), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n265), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n578), .B1(new_n613), .B2(new_n577), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n614), .A2(new_n579), .A3(new_n580), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n570), .A2(KEYINPUT29), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n570), .B1(new_n602), .B2(new_n577), .ZN(new_n618));
  INV_X1    g432(.A(new_n580), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n577), .A2(KEYINPUT71), .A3(new_n578), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n588), .A2(new_n619), .A3(new_n620), .A4(new_n570), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT29), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n617), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(G472), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n611), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT32), .B1(new_n606), .B2(new_n607), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n503), .B(new_n566), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n454), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n232), .ZN(G3));
  AND3_X1   g444(.A1(new_n347), .A2(new_n344), .A3(new_n351), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n344), .B1(new_n347), .B2(new_n351), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n453), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT97), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n635), .B(new_n453), .C1(new_n631), .C2(new_n632), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n637));
  INV_X1    g451(.A(new_n404), .ZN(new_n638));
  AOI211_X1 g452(.A(KEYINPUT20), .B(new_n638), .C1(new_n397), .C2(new_n402), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n387), .A2(new_n396), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n401), .ZN(new_n641));
  AOI21_X1  g455(.A(G902), .B1(new_n641), .B2(new_n397), .ZN(new_n642));
  INV_X1    g456(.A(G475), .ZN(new_n643));
  OAI22_X1  g457(.A1(new_n637), .A2(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n438), .A2(new_n645), .A3(new_n439), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT98), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n438), .A2(new_n439), .A3(new_n648), .A4(new_n645), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n433), .B1(new_n650), .B2(new_n436), .ZN(new_n651));
  OAI211_X1 g465(.A(KEYINPUT99), .B(new_n437), .C1(new_n426), .C2(new_n432), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(KEYINPUT33), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n442), .A2(G902), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n647), .A2(new_n649), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n442), .B1(new_n440), .B2(G902), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n644), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n451), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n634), .A2(new_n636), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n606), .A2(new_n607), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n602), .A2(new_n603), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT31), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n602), .A2(KEYINPUT31), .A3(new_n603), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n589), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n666), .B2(G902), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n566), .A2(new_n661), .A3(new_n667), .A4(new_n503), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT34), .B(G104), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  INV_X1    g485(.A(new_n444), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n412), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n451), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n634), .A2(new_n636), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n668), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT35), .B(G107), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n491), .A2(KEYINPUT36), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT75), .B1(new_n484), .B2(new_n465), .ZN(new_n681));
  INV_X1    g495(.A(new_n490), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n489), .B(new_n490), .C1(KEYINPUT36), .C2(new_n491), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n683), .A2(new_n684), .A3(new_n502), .ZN(new_n685));
  AOI211_X1 g499(.A(new_n679), .B(new_n685), .C1(new_n497), .C2(new_n499), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n495), .A2(new_n496), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n499), .A3(new_n455), .ZN(new_n688));
  INV_X1    g502(.A(new_n685), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT100), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n661), .A3(new_n566), .A4(new_n667), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n454), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT37), .B(G110), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G12));
  AND2_X1   g509(.A1(new_n634), .A2(new_n636), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n606), .A2(new_n610), .B1(new_n624), .B2(G472), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n609), .B1(new_n666), .B2(new_n608), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n686), .A2(new_n690), .ZN(new_n700));
  INV_X1    g514(.A(new_n566), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n449), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n447), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n673), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n696), .A2(new_n699), .A3(new_n702), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  XOR2_X1   g524(.A(new_n356), .B(KEYINPUT38), .Z(new_n711));
  INV_X1    g525(.A(new_n662), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n570), .B1(new_n613), .B2(new_n577), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT101), .Z(new_n714));
  OAI21_X1  g528(.A(new_n341), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G472), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n698), .A2(new_n611), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n688), .A2(new_n689), .ZN(new_n718));
  INV_X1    g532(.A(new_n453), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n718), .A2(new_n444), .A3(new_n412), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n711), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n706), .B(KEYINPUT39), .Z(new_n725));
  NOR2_X1   g539(.A1(new_n701), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT40), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  NOR2_X1   g543(.A1(new_n626), .A2(new_n627), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n644), .A2(new_n657), .A3(new_n706), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n696), .A2(new_n702), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  INV_X1    g548(.A(new_n503), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n697), .B2(new_n698), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n341), .B1(new_n559), .B2(new_n564), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(new_n504), .A3(new_n565), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n660), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT41), .B(G113), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  OR2_X1    g557(.A1(new_n675), .A2(new_n740), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  NOR2_X1   g559(.A1(new_n730), .A2(new_n700), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n452), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n634), .A2(new_n636), .A3(new_n739), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT103), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n634), .A2(new_n750), .A3(new_n636), .A4(new_n739), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n208), .ZN(G21));
  NOR2_X1   g567(.A1(new_n412), .A2(new_n444), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n634), .A2(new_n636), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(G472), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n606), .B2(new_n341), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n664), .A2(new_n665), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n615), .A2(new_n570), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n608), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n451), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n739), .A3(new_n762), .A4(new_n503), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n755), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NAND2_X1  g579(.A1(new_n749), .A2(new_n751), .ZN(new_n766));
  INV_X1    g580(.A(new_n760), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n667), .A3(new_n718), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n731), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n644), .A2(new_n657), .A3(KEYINPUT104), .A4(new_n706), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  NAND2_X1  g589(.A1(new_n699), .A2(new_n503), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT107), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n770), .A2(new_n771), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(KEYINPUT42), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n719), .B1(new_n343), .B2(new_n344), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n566), .A2(new_n780), .A3(new_n345), .A4(new_n355), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n736), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n777), .A2(new_n779), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n345), .A2(new_n780), .A3(new_n355), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n736), .A3(new_n566), .A4(new_n778), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n787), .A2(KEYINPUT106), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT106), .B1(new_n787), .B2(new_n789), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  NAND4_X1  g607(.A1(new_n786), .A2(new_n736), .A3(new_n566), .A4(new_n708), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  NAND2_X1  g609(.A1(new_n412), .A2(new_n657), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT43), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT109), .Z(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n797), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT108), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n667), .A2(new_n661), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n718), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OR3_X1    g619(.A1(new_n805), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n556), .A2(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n556), .A2(KEYINPUT45), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(G469), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(G469), .A2(G902), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT46), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n565), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n809), .A2(KEYINPUT46), .A3(new_n810), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n505), .B(new_n725), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT110), .B1(new_n805), .B2(KEYINPUT44), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n345), .A2(new_n780), .A3(new_n355), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n805), .B2(KEYINPUT44), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n806), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  AOI21_X1  g634(.A(new_n505), .B1(new_n813), .B2(new_n814), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n658), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n730), .A2(new_n735), .A3(new_n824), .A4(new_n706), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n823), .A2(new_n817), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  NOR2_X1   g641(.A1(new_n802), .A2(new_n705), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n503), .A3(new_n761), .ZN(new_n829));
  INV_X1    g643(.A(new_n766), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n786), .A2(new_n739), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT117), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n717), .A2(new_n735), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n835), .A2(new_n447), .A3(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n446), .B(G953), .C1(new_n837), .C2(new_n824), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n833), .A2(KEYINPUT120), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n777), .A2(new_n784), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n828), .A2(new_n840), .A3(new_n835), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT48), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT120), .B1(new_n833), .B2(new_n838), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n711), .A2(new_n719), .A3(new_n739), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n829), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n848), .B2(KEYINPUT50), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(KEYINPUT50), .B2(new_n848), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n738), .A2(new_n565), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n823), .B1(new_n504), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n829), .A2(new_n817), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n848), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n718), .A2(new_n828), .A3(new_n761), .A4(new_n835), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n644), .A2(new_n657), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n858), .B1(new_n837), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT51), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT51), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n845), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n566), .A2(new_n688), .A3(new_n689), .A4(new_n706), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT115), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n755), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n717), .A3(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n774), .A2(new_n872), .A3(new_n709), .A4(new_n733), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n873), .B(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n660), .A2(new_n740), .B1(new_n454), .B2(new_n692), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n356), .A2(new_n453), .ZN(new_n879));
  INV_X1    g693(.A(new_n674), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n668), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n878), .A2(new_n744), .A3(new_n764), .A4(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n659), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n879), .A2(new_n668), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT112), .B1(new_n885), .B2(new_n629), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n356), .A2(new_n452), .A3(new_n453), .ZN(new_n887));
  INV_X1    g701(.A(new_n628), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT112), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n553), .A2(new_n555), .ZN(new_n891));
  INV_X1    g705(.A(new_n530), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n562), .B2(new_n563), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n891), .B(G469), .C1(new_n893), .C2(new_n547), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n810), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n503), .B(new_n504), .C1(new_n812), .C2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n803), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n453), .A3(new_n356), .A4(new_n659), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n889), .A2(new_n890), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n886), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n883), .A2(new_n900), .A3(new_n752), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n445), .A2(new_n707), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n746), .A2(new_n782), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT113), .B1(new_n773), .B2(new_n782), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n905));
  NOR4_X1   g719(.A1(new_n781), .A2(new_n768), .A3(new_n772), .A4(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n903), .B(new_n794), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n787), .A2(new_n789), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT106), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n787), .A2(KEYINPUT106), .A3(new_n789), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n907), .B1(new_n912), .B2(new_n785), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n876), .B1(new_n901), .B2(new_n913), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n675), .A2(new_n740), .B1(new_n755), .B2(new_n763), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n915), .A2(new_n877), .A3(new_n881), .ZN(new_n916));
  INV_X1    g730(.A(new_n752), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n886), .A4(new_n899), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n699), .A2(new_n691), .A3(new_n902), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n794), .B1(new_n781), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n904), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n773), .A2(new_n782), .A3(KEYINPUT113), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n792), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n918), .A2(new_n924), .A3(KEYINPUT114), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n875), .B1(new_n914), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT53), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n873), .B(KEYINPUT52), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n774), .A2(new_n709), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT52), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n901), .A2(KEYINPUT53), .A3(new_n913), .A4(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT54), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n928), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n926), .B1(new_n927), .B2(new_n931), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT114), .B1(new_n918), .B2(new_n924), .ZN(new_n938));
  NOR4_X1   g752(.A1(new_n752), .A2(new_n915), .A3(new_n877), .A4(new_n881), .ZN(new_n939));
  INV_X1    g753(.A(new_n900), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n913), .A2(new_n939), .A3(new_n876), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT53), .B1(new_n942), .B2(new_n875), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n936), .B1(new_n944), .B2(new_n935), .ZN(new_n945));
  OAI22_X1  g759(.A1(new_n867), .A2(new_n945), .B1(G952), .B2(G953), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n851), .B(KEYINPUT49), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n796), .A2(new_n719), .A3(new_n505), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n711), .A2(new_n836), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n946), .A2(new_n949), .ZN(G75));
  NAND2_X1  g764(.A1(new_n928), .A2(new_n934), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(G210), .A3(G902), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT56), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n277), .B(KEYINPUT121), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT55), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(new_n317), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n952), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n952), .B2(new_n953), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n448), .A2(G952), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G51));
  XNOR2_X1  g774(.A(new_n951), .B(new_n935), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n810), .B(KEYINPUT57), .ZN(new_n962));
  OAI22_X1  g776(.A1(new_n961), .A2(new_n962), .B1(new_n559), .B2(new_n564), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n951), .A2(G902), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(new_n809), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n959), .B1(new_n963), .B2(new_n965), .ZN(G54));
  INV_X1    g780(.A(new_n959), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT58), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n964), .A2(new_n968), .A3(new_n643), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n969), .B2(new_n403), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n403), .B2(new_n969), .ZN(G60));
  AND3_X1   g785(.A1(new_n647), .A2(new_n649), .A3(new_n653), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT59), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n967), .B1(new_n961), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n972), .B1(new_n945), .B2(new_n974), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G63));
  NAND2_X1  g792(.A1(new_n683), .A2(new_n684), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n435), .A2(new_n341), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n980), .B(new_n983), .C1(new_n943), .C2(new_n933), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n928), .B2(new_n934), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n967), .B(new_n984), .C1(new_n986), .C2(new_n501), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(KEYINPUT124), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n983), .B1(new_n943), .B2(new_n933), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n959), .B1(new_n989), .B2(new_n500), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT123), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT61), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n990), .A2(new_n993), .A3(new_n984), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n988), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n988), .B2(new_n994), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(G66));
  OAI21_X1  g811(.A(G953), .B1(new_n450), .B2(new_n315), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n901), .B2(G953), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n954), .B1(G898), .B2(new_n448), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G69));
  NOR2_X1   g815(.A1(new_n598), .A2(new_n601), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n593), .B2(new_n595), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(new_n398), .Z(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n819), .A2(new_n826), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n774), .A2(new_n709), .A3(new_n733), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n840), .A2(new_n871), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n815), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1007), .A2(new_n792), .A3(new_n794), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n448), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(G900), .B2(new_n448), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT125), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1005), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n728), .A2(new_n1007), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n817), .B(new_n776), .C1(new_n658), .C2(new_n673), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1006), .B1(new_n726), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n448), .A3(new_n1005), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n448), .B1(G227), .B2(G900), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1017), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1026), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1025), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1028), .B1(new_n1016), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1027), .A2(new_n1030), .ZN(G72));
  XNOR2_X1  g845(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n756), .A2(new_n341), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n1032), .B(new_n1033), .Z(new_n1034));
  INV_X1    g848(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1035), .B1(new_n1024), .B2(new_n918), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n602), .A2(new_n577), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT127), .Z(new_n1038));
  NAND3_X1  g852(.A1(new_n1036), .A2(new_n570), .A3(new_n1038), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1035), .B1(new_n1040), .B2(new_n918), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1038), .A2(new_n570), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n959), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n944), .ZN(new_n1045));
  INV_X1    g859(.A(new_n618), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1034), .B1(new_n1046), .B2(new_n662), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1044), .B1(new_n1045), .B2(new_n1047), .ZN(G57));
endmodule


