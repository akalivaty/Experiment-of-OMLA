

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U325 ( .A(n377), .B(n376), .ZN(n531) );
  XNOR2_X1 U326 ( .A(n375), .B(KEYINPUT114), .ZN(n376) );
  XNOR2_X1 U327 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U328 ( .A(n335), .B(n314), .ZN(n318) );
  XOR2_X1 U329 ( .A(n328), .B(n327), .Z(n561) );
  XNOR2_X1 U330 ( .A(n561), .B(KEYINPUT84), .ZN(n548) );
  XNOR2_X1 U331 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U332 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(G1GAT), .B(KEYINPUT77), .Z(n349) );
  XOR2_X1 U334 ( .A(G22GAT), .B(G155GAT), .Z(n419) );
  XOR2_X1 U335 ( .A(G15GAT), .B(G127GAT), .Z(n448) );
  XOR2_X1 U336 ( .A(n419), .B(n448), .Z(n294) );
  NAND2_X1 U337 ( .A1(G231GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n349), .B(n295), .ZN(n306) );
  XOR2_X1 U340 ( .A(KEYINPUT15), .B(KEYINPUT85), .Z(n301) );
  XNOR2_X1 U341 ( .A(G57GAT), .B(KEYINPUT78), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n296), .B(KEYINPUT13), .ZN(n333) );
  XOR2_X1 U343 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n298) );
  XNOR2_X1 U344 ( .A(G71GAT), .B(G64GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n333), .B(n299), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U348 ( .A(G8GAT), .B(G183GAT), .Z(n378) );
  XOR2_X1 U349 ( .A(n302), .B(n378), .Z(n304) );
  XNOR2_X1 U350 ( .A(G211GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U352 ( .A(n306), .B(n305), .Z(n476) );
  INV_X1 U353 ( .A(n476), .ZN(n583) );
  XNOR2_X1 U354 ( .A(G50GAT), .B(KEYINPUT81), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n307), .B(G162GAT), .ZN(n432) );
  XOR2_X1 U356 ( .A(G92GAT), .B(G218GAT), .Z(n309) );
  XNOR2_X1 U357 ( .A(G36GAT), .B(G190GAT), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n381) );
  XNOR2_X1 U359 ( .A(n432), .B(n381), .ZN(n328) );
  XOR2_X1 U360 ( .A(G85GAT), .B(KEYINPUT80), .Z(n311) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G106GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n335) );
  NAND2_X1 U363 ( .A1(G232GAT), .A2(G233GAT), .ZN(n313) );
  INV_X1 U364 ( .A(G134GAT), .ZN(n312) );
  XOR2_X1 U365 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n316) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(G29GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U368 ( .A(KEYINPUT76), .B(n317), .Z(n363) );
  XNOR2_X1 U369 ( .A(n318), .B(n363), .ZN(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n320) );
  XNOR2_X1 U371 ( .A(KEYINPUT11), .B(KEYINPUT83), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U373 ( .A(KEYINPUT82), .B(KEYINPUT68), .Z(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U378 ( .A(KEYINPUT36), .B(n548), .ZN(n493) );
  NOR2_X1 U379 ( .A1(n583), .A2(n493), .ZN(n331) );
  XOR2_X1 U380 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n329) );
  XNOR2_X1 U381 ( .A(KEYINPUT69), .B(n329), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n345) );
  XNOR2_X1 U383 ( .A(G176GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n332), .B(G64GAT), .ZN(n385) );
  XOR2_X1 U385 ( .A(n385), .B(n333), .Z(n337) );
  XNOR2_X1 U386 ( .A(G78GAT), .B(KEYINPUT79), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n334), .B(G148GAT), .ZN(n420) );
  XNOR2_X1 U388 ( .A(n420), .B(n335), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n344) );
  XOR2_X1 U390 ( .A(G120GAT), .B(G71GAT), .Z(n449) );
  XOR2_X1 U391 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n339) );
  XNOR2_X1 U392 ( .A(G92GAT), .B(KEYINPUT31), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U394 ( .A(n449), .B(n340), .Z(n342) );
  NAND2_X1 U395 ( .A1(G230GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U397 ( .A(n344), .B(n343), .Z(n578) );
  NAND2_X1 U398 ( .A1(n345), .A2(n578), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n346), .B(KEYINPUT113), .ZN(n366) );
  XOR2_X1 U400 ( .A(KEYINPUT74), .B(KEYINPUT72), .Z(n348) );
  XNOR2_X1 U401 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U403 ( .A(G50GAT), .B(G36GAT), .Z(n351) );
  XNOR2_X1 U404 ( .A(n349), .B(KEYINPUT75), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U406 ( .A(n353), .B(n352), .Z(n355) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U409 ( .A(G15GAT), .B(G197GAT), .Z(n357) );
  XNOR2_X1 U410 ( .A(G22GAT), .B(G141GAT), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U412 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U413 ( .A(KEYINPUT73), .B(KEYINPUT30), .Z(n361) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G113GAT), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U417 ( .A(n365), .B(n364), .Z(n507) );
  INV_X1 U418 ( .A(n507), .ZN(n573) );
  NAND2_X1 U419 ( .A1(n366), .A2(n573), .ZN(n374) );
  INV_X1 U420 ( .A(n561), .ZN(n371) );
  XNOR2_X1 U421 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n368) );
  XOR2_X1 U422 ( .A(KEYINPUT41), .B(n578), .Z(n564) );
  NOR2_X1 U423 ( .A1(n573), .A2(n564), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  NAND2_X1 U425 ( .A1(n583), .A2(n369), .ZN(n370) );
  NOR2_X1 U426 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT47), .B(n372), .ZN(n373) );
  NAND2_X1 U428 ( .A1(n374), .A2(n373), .ZN(n377) );
  XOR2_X1 U429 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n375) );
  XOR2_X1 U430 ( .A(KEYINPUT97), .B(n378), .Z(n380) );
  NAND2_X1 U431 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U433 ( .A(n382), .B(n381), .Z(n387) );
  XOR2_X1 U434 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n384) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n384), .B(n383), .ZN(n443) );
  XNOR2_X1 U437 ( .A(n443), .B(n385), .ZN(n386) );
  XNOR2_X1 U438 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U439 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n389) );
  XNOR2_X1 U440 ( .A(KEYINPUT91), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(n390), .ZN(n424) );
  INV_X1 U443 ( .A(n424), .ZN(n391) );
  XOR2_X1 U444 ( .A(n392), .B(n391), .Z(n484) );
  INV_X1 U445 ( .A(n484), .ZN(n521) );
  XOR2_X1 U446 ( .A(n521), .B(KEYINPUT121), .Z(n393) );
  NOR2_X1 U447 ( .A1(n531), .A2(n393), .ZN(n394) );
  XNOR2_X1 U448 ( .A(KEYINPUT54), .B(n394), .ZN(n417) );
  XOR2_X1 U449 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n396) );
  XNOR2_X1 U450 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U452 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n398) );
  XNOR2_X1 U453 ( .A(G127GAT), .B(KEYINPUT94), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U456 ( .A(G148GAT), .B(G155GAT), .Z(n402) );
  XNOR2_X1 U457 ( .A(G120GAT), .B(G162GAT), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U460 ( .A(n405), .B(KEYINPUT6), .Z(n409) );
  XOR2_X1 U461 ( .A(KEYINPUT92), .B(KEYINPUT3), .Z(n407) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n431) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(n431), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT0), .B(KEYINPUT86), .Z(n411) );
  XNOR2_X1 U467 ( .A(G113GAT), .B(G134GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n450) );
  XOR2_X1 U469 ( .A(G85GAT), .B(n450), .Z(n413) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U472 ( .A(G29GAT), .B(n414), .Z(n415) );
  XOR2_X1 U473 ( .A(n416), .B(n415), .Z(n480) );
  INV_X1 U474 ( .A(n480), .ZN(n532) );
  NAND2_X1 U475 ( .A1(n417), .A2(n532), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n418), .B(KEYINPUT65), .ZN(n572) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U480 ( .A(n424), .B(n423), .Z(n436) );
  XOR2_X1 U481 ( .A(G204GAT), .B(KEYINPUT24), .Z(n426) );
  XNOR2_X1 U482 ( .A(G218GAT), .B(G106GAT), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U484 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n428) );
  XNOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT93), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n470) );
  NAND2_X1 U491 ( .A1(n572), .A2(n470), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n437), .B(KEYINPUT55), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n438), .B(KEYINPUT122), .ZN(n456) );
  XOR2_X1 U494 ( .A(KEYINPUT67), .B(G190GAT), .Z(n440) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(G99GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n455) );
  XOR2_X1 U497 ( .A(G183GAT), .B(KEYINPUT88), .Z(n442) );
  XNOR2_X1 U498 ( .A(KEYINPUT87), .B(KEYINPUT20), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n447) );
  XOR2_X1 U500 ( .A(G176GAT), .B(n443), .Z(n445) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U507 ( .A(n455), .B(n454), .Z(n524) );
  INV_X1 U508 ( .A(n524), .ZN(n537) );
  NAND2_X1 U509 ( .A1(n456), .A2(n537), .ZN(n569) );
  NOR2_X1 U510 ( .A1(n569), .A2(n548), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n458) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n457) );
  XOR2_X1 U513 ( .A(KEYINPUT102), .B(KEYINPUT34), .Z(n482) );
  AND2_X1 U514 ( .A1(n507), .A2(n578), .ZN(n497) );
  NAND2_X1 U515 ( .A1(n484), .A2(n537), .ZN(n461) );
  XOR2_X1 U516 ( .A(KEYINPUT99), .B(n461), .Z(n462) );
  NAND2_X1 U517 ( .A1(n470), .A2(n462), .ZN(n463) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n463), .Z(n467) );
  XOR2_X1 U519 ( .A(n521), .B(KEYINPUT98), .Z(n464) );
  XNOR2_X1 U520 ( .A(n464), .B(KEYINPUT27), .ZN(n534) );
  NOR2_X1 U521 ( .A1(n537), .A2(n470), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n465), .B(KEYINPUT26), .ZN(n571) );
  NAND2_X1 U523 ( .A1(n534), .A2(n571), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U525 ( .A(KEYINPUT100), .B(n468), .Z(n469) );
  NAND2_X1 U526 ( .A1(n469), .A2(n532), .ZN(n475) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT71), .ZN(n471) );
  XOR2_X1 U528 ( .A(n471), .B(KEYINPUT28), .Z(n527) );
  INV_X1 U529 ( .A(n527), .ZN(n535) );
  NOR2_X1 U530 ( .A1(n537), .A2(n535), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n534), .A2(n472), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n480), .A2(n473), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n494) );
  NAND2_X1 U534 ( .A1(n548), .A2(n476), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT16), .B(n477), .ZN(n478) );
  NOR2_X1 U536 ( .A1(n494), .A2(n478), .ZN(n508) );
  NAND2_X1 U537 ( .A1(n497), .A2(n508), .ZN(n479) );
  XNOR2_X1 U538 ( .A(KEYINPUT101), .B(n479), .ZN(n490) );
  NAND2_X1 U539 ( .A1(n490), .A2(n480), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  XOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT103), .Z(n486) );
  NAND2_X1 U543 ( .A1(n490), .A2(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n488) );
  NAND2_X1 U546 ( .A1(n490), .A2(n537), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n489), .ZN(G1326GAT) );
  XOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT105), .Z(n492) );
  NAND2_X1 U550 ( .A1(n490), .A2(n535), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  NOR2_X1 U552 ( .A1(n493), .A2(n494), .ZN(n495) );
  NAND2_X1 U553 ( .A1(n495), .A2(n583), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n496), .B(KEYINPUT37), .ZN(n518) );
  NAND2_X1 U555 ( .A1(n497), .A2(n518), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n498), .B(KEYINPUT38), .ZN(n504) );
  NOR2_X1 U557 ( .A1(n504), .A2(n532), .ZN(n500) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n504), .A2(n521), .ZN(n501) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n501), .Z(G1329GAT) );
  NOR2_X1 U562 ( .A1(n524), .A2(n504), .ZN(n502) );
  XOR2_X1 U563 ( .A(KEYINPUT40), .B(n502), .Z(n503) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NOR2_X1 U565 ( .A1(n504), .A2(n527), .ZN(n505) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n505), .Z(n506) );
  XNOR2_X1 U567 ( .A(KEYINPUT106), .B(n506), .ZN(G1331GAT) );
  NOR2_X1 U568 ( .A1(n564), .A2(n507), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n508), .A2(n517), .ZN(n514) );
  NOR2_X1 U570 ( .A1(n532), .A2(n514), .ZN(n509) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT42), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n521), .A2(n514), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(G1333GAT) );
  NOR2_X1 U576 ( .A1(n524), .A2(n514), .ZN(n513) );
  XOR2_X1 U577 ( .A(G71GAT), .B(n513), .Z(G1334GAT) );
  NOR2_X1 U578 ( .A1(n527), .A2(n514), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n526) );
  NOR2_X1 U582 ( .A1(n532), .A2(n526), .ZN(n519) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n519), .Z(n520) );
  XNOR2_X1 U584 ( .A(KEYINPUT108), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n526), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n526), .ZN(n525) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U591 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U593 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  NOR2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n551) );
  NOR2_X1 U596 ( .A1(n535), .A2(n551), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U598 ( .A(KEYINPUT115), .B(n538), .Z(n547) );
  NOR2_X1 U599 ( .A1(n573), .A2(n547), .ZN(n539) );
  XOR2_X1 U600 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  NOR2_X1 U601 ( .A1(n564), .A2(n547), .ZN(n541) );
  XNOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n544) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n546) );
  NOR2_X1 U608 ( .A1(n583), .A2(n547), .ZN(n545) );
  XOR2_X1 U609 ( .A(n546), .B(n545), .Z(G1342GAT) );
  NOR2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  INV_X1 U613 ( .A(n551), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n552), .A2(n571), .ZN(n560) );
  NOR2_X1 U615 ( .A1(n573), .A2(n560), .ZN(n554) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  NOR2_X1 U618 ( .A1(n564), .A2(n560), .ZN(n556) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n583), .A2(n560), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT120), .B(n558), .Z(n559) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NOR2_X1 U627 ( .A1(n573), .A2(n569), .ZN(n563) );
  XOR2_X1 U628 ( .A(G169GAT), .B(n563), .Z(G1348GAT) );
  NOR2_X1 U629 ( .A1(n569), .A2(n564), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n566) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NOR2_X1 U634 ( .A1(n583), .A2(n569), .ZN(n570) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n570), .Z(G1350GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n585) );
  NOR2_X1 U637 ( .A1(n585), .A2(n573), .ZN(n577) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n585), .A2(n578), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  NOR2_X1 U649 ( .A1(n493), .A2(n585), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

