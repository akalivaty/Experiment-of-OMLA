

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U322 ( .A(n325), .B(n324), .ZN(n527) );
  XNOR2_X1 U323 ( .A(n438), .B(n437), .ZN(n535) );
  XNOR2_X1 U324 ( .A(KEYINPUT118), .B(KEYINPUT47), .ZN(n430) );
  XNOR2_X1 U325 ( .A(n431), .B(n430), .ZN(n436) );
  XNOR2_X1 U326 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n437) );
  XNOR2_X1 U327 ( .A(n448), .B(n367), .ZN(n368) );
  NOR2_X1 U328 ( .A1(n522), .A2(n451), .ZN(n457) );
  XNOR2_X1 U329 ( .A(n369), .B(n368), .ZN(n463) );
  INV_X1 U330 ( .A(G211GAT), .ZN(n454) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(n579) );
  XNOR2_X1 U332 ( .A(n576), .B(n370), .ZN(n563) );
  XOR2_X1 U333 ( .A(n475), .B(KEYINPUT28), .Z(n529) );
  XNOR2_X1 U334 ( .A(n454), .B(KEYINPUT126), .ZN(n455) );
  XNOR2_X1 U335 ( .A(n456), .B(n455), .ZN(G1354GAT) );
  INV_X1 U336 ( .A(KEYINPUT123), .ZN(n453) );
  XOR2_X1 U337 ( .A(G211GAT), .B(KEYINPUT21), .Z(n291) );
  XNOR2_X1 U338 ( .A(G197GAT), .B(G218GAT), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n291), .B(n290), .ZN(n444) );
  XOR2_X1 U340 ( .A(G141GAT), .B(G22GAT), .Z(n385) );
  XOR2_X1 U341 ( .A(n444), .B(n385), .Z(n293) );
  NAND2_X1 U342 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U344 ( .A(n294), .B(G204GAT), .Z(n297) );
  XNOR2_X1 U345 ( .A(G50GAT), .B(KEYINPUT78), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n295), .B(G162GAT), .ZN(n405) );
  XNOR2_X1 U347 ( .A(n405), .B(KEYINPUT22), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U349 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n299) );
  XNOR2_X1 U350 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(n301), .B(n300), .Z(n306) );
  XNOR2_X1 U353 ( .A(G106GAT), .B(G78GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n302), .B(G148GAT), .ZN(n366) );
  XOR2_X1 U355 ( .A(G155GAT), .B(KEYINPUT3), .Z(n304) );
  XNOR2_X1 U356 ( .A(KEYINPUT2), .B(KEYINPUT93), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n334) );
  XNOR2_X1 U358 ( .A(n366), .B(n334), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n475) );
  XOR2_X1 U360 ( .A(G183GAT), .B(KEYINPUT89), .Z(n308) );
  XNOR2_X1 U361 ( .A(KEYINPUT20), .B(KEYINPUT67), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n325) );
  XOR2_X1 U363 ( .A(KEYINPUT87), .B(G134GAT), .Z(n310) );
  XNOR2_X1 U364 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U366 ( .A(G113GAT), .B(n311), .Z(n338) );
  XOR2_X1 U367 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n313) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n445) );
  XOR2_X1 U370 ( .A(G176GAT), .B(n445), .Z(n315) );
  NAND2_X1 U371 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n338), .B(n316), .ZN(n323) );
  XOR2_X1 U374 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n318) );
  XNOR2_X1 U375 ( .A(G15GAT), .B(G99GAT), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U377 ( .A(n319), .B(G190GAT), .Z(n321) );
  XOR2_X1 U378 ( .A(G120GAT), .B(G71GAT), .Z(n355) );
  XNOR2_X1 U379 ( .A(G43GAT), .B(n355), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  NOR2_X1 U382 ( .A1(n475), .A2(n527), .ZN(n327) );
  XNOR2_X1 U383 ( .A(KEYINPUT26), .B(KEYINPUT101), .ZN(n326) );
  XOR2_X1 U384 ( .A(n327), .B(n326), .Z(n551) );
  XOR2_X1 U385 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n329) );
  XNOR2_X1 U386 ( .A(KEYINPUT4), .B(KEYINPUT98), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U388 ( .A(KEYINPUT94), .B(KEYINPUT1), .Z(n331) );
  XNOR2_X1 U389 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U391 ( .A(n333), .B(n332), .Z(n340) );
  XOR2_X1 U392 ( .A(n334), .B(KEYINPUT6), .Z(n336) );
  NAND2_X1 U393 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n348) );
  XOR2_X1 U397 ( .A(G57GAT), .B(G120GAT), .Z(n342) );
  XNOR2_X1 U398 ( .A(G141GAT), .B(G1GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U400 ( .A(G85GAT), .B(G162GAT), .Z(n344) );
  XNOR2_X1 U401 ( .A(G29GAT), .B(G148GAT), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U403 ( .A(n346), .B(n345), .Z(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n522) );
  INV_X1 U405 ( .A(KEYINPUT72), .ZN(n349) );
  NAND2_X1 U406 ( .A1(n349), .A2(KEYINPUT13), .ZN(n352) );
  INV_X1 U407 ( .A(KEYINPUT13), .ZN(n350) );
  NAND2_X1 U408 ( .A1(n350), .A2(KEYINPUT72), .ZN(n351) );
  NAND2_X1 U409 ( .A1(n352), .A2(n351), .ZN(n354) );
  XNOR2_X1 U410 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n423) );
  XOR2_X1 U412 ( .A(n423), .B(n355), .Z(n357) );
  NAND2_X1 U413 ( .A1(G230GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U415 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n359) );
  XNOR2_X1 U416 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n358) );
  XOR2_X1 U417 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n369) );
  XOR2_X1 U419 ( .A(G92GAT), .B(KEYINPUT75), .Z(n363) );
  XNOR2_X1 U420 ( .A(G204GAT), .B(G64GAT), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(n364), .ZN(n448) );
  XNOR2_X1 U423 ( .A(G99GAT), .B(G85GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n365), .B(KEYINPUT74), .ZN(n400) );
  XNOR2_X1 U425 ( .A(n366), .B(n400), .ZN(n367) );
  INV_X1 U426 ( .A(n463), .ZN(n576) );
  XNOR2_X1 U427 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n370) );
  XOR2_X1 U428 ( .A(KEYINPUT69), .B(KEYINPUT71), .Z(n372) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U431 ( .A(n373), .B(KEYINPUT30), .Z(n381) );
  XOR2_X1 U432 ( .A(G113GAT), .B(G197GAT), .Z(n375) );
  XNOR2_X1 U433 ( .A(G36GAT), .B(G50GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U435 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n377) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(G8GAT), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U440 ( .A(G15GAT), .B(G1GAT), .Z(n414) );
  XOR2_X1 U441 ( .A(n382), .B(n414), .Z(n387) );
  XOR2_X1 U442 ( .A(G29GAT), .B(G43GAT), .Z(n384) );
  XNOR2_X1 U443 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n406) );
  XNOR2_X1 U445 ( .A(n406), .B(n385), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n570) );
  NOR2_X1 U447 ( .A1(n563), .A2(n570), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n388), .B(KEYINPUT46), .ZN(n429) );
  XOR2_X1 U449 ( .A(KEYINPUT79), .B(KEYINPUT11), .Z(n390) );
  XNOR2_X1 U450 ( .A(KEYINPUT66), .B(KEYINPUT80), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U452 ( .A(KEYINPUT9), .B(KEYINPUT68), .Z(n392) );
  XNOR2_X1 U453 ( .A(G134GAT), .B(G92GAT), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U455 ( .A(n394), .B(n393), .Z(n399) );
  XOR2_X1 U456 ( .A(KEYINPUT81), .B(KEYINPUT10), .Z(n396) );
  NAND2_X1 U457 ( .A1(G232GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U459 ( .A(G106GAT), .B(n397), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n404) );
  XOR2_X1 U461 ( .A(G36GAT), .B(G190GAT), .Z(n439) );
  XOR2_X1 U462 ( .A(n439), .B(KEYINPUT82), .Z(n402) );
  XNOR2_X1 U463 ( .A(G218GAT), .B(n400), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U465 ( .A(n404), .B(n403), .Z(n408) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n465) );
  INV_X1 U468 ( .A(n465), .ZN(n560) );
  XOR2_X1 U469 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n410) );
  XNOR2_X1 U470 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n418) );
  XOR2_X1 U472 ( .A(G155GAT), .B(G78GAT), .Z(n412) );
  XNOR2_X1 U473 ( .A(G127GAT), .B(G71GAT), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U475 ( .A(n413), .B(G211GAT), .Z(n416) );
  XNOR2_X1 U476 ( .A(G22GAT), .B(n414), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n427) );
  XOR2_X1 U479 ( .A(KEYINPUT15), .B(KEYINPUT86), .Z(n420) );
  NAND2_X1 U480 ( .A1(G231GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U482 ( .A(G8GAT), .B(G183GAT), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n421), .B(KEYINPUT83), .ZN(n442) );
  XOR2_X1 U484 ( .A(n422), .B(n442), .Z(n425) );
  XNOR2_X1 U485 ( .A(G64GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n568) );
  NAND2_X1 U488 ( .A1(n560), .A2(n568), .ZN(n428) );
  OR2_X1 U489 ( .A1(n429), .A2(n428), .ZN(n431) );
  XOR2_X1 U490 ( .A(KEYINPUT36), .B(n465), .Z(n580) );
  NOR2_X1 U491 ( .A1(n580), .A2(n568), .ZN(n432) );
  XNOR2_X1 U492 ( .A(KEYINPUT45), .B(n432), .ZN(n433) );
  NAND2_X1 U493 ( .A1(n433), .A2(n570), .ZN(n434) );
  NOR2_X1 U494 ( .A1(n434), .A2(n463), .ZN(n435) );
  NOR2_X1 U495 ( .A1(n436), .A2(n435), .ZN(n438) );
  XOR2_X1 U496 ( .A(KEYINPUT99), .B(n439), .Z(n441) );
  NAND2_X1 U497 ( .A1(G226GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U499 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n467) );
  NOR2_X1 U503 ( .A1(n535), .A2(n467), .ZN(n450) );
  XOR2_X1 U504 ( .A(n450), .B(KEYINPUT54), .Z(n451) );
  NAND2_X1 U505 ( .A1(n551), .A2(n457), .ZN(n452) );
  NOR2_X1 U506 ( .A1(n579), .A2(n568), .ZN(n456) );
  NAND2_X1 U507 ( .A1(n457), .A2(n475), .ZN(n458) );
  XNOR2_X1 U508 ( .A(n458), .B(KEYINPUT55), .ZN(n459) );
  NAND2_X1 U509 ( .A1(n459), .A2(n527), .ZN(n567) );
  NOR2_X1 U510 ( .A1(n560), .A2(n567), .ZN(n460) );
  XNOR2_X1 U511 ( .A(G190GAT), .B(n460), .ZN(n462) );
  INV_X1 U512 ( .A(KEYINPUT58), .ZN(n461) );
  XNOR2_X1 U513 ( .A(n462), .B(n461), .ZN(G1351GAT) );
  XOR2_X1 U514 ( .A(KEYINPUT34), .B(KEYINPUT105), .Z(n483) );
  NOR2_X1 U515 ( .A1(n463), .A2(n570), .ZN(n464) );
  XNOR2_X1 U516 ( .A(n464), .B(KEYINPUT77), .ZN(n496) );
  NOR2_X1 U517 ( .A1(n465), .A2(n568), .ZN(n466) );
  XNOR2_X1 U518 ( .A(n466), .B(KEYINPUT16), .ZN(n480) );
  INV_X1 U519 ( .A(n467), .ZN(n525) );
  NAND2_X1 U520 ( .A1(n527), .A2(n525), .ZN(n468) );
  NAND2_X1 U521 ( .A1(n468), .A2(n475), .ZN(n469) );
  XNOR2_X1 U522 ( .A(n469), .B(KEYINPUT102), .ZN(n470) );
  XNOR2_X1 U523 ( .A(n470), .B(KEYINPUT25), .ZN(n472) );
  XNOR2_X1 U524 ( .A(n525), .B(KEYINPUT27), .ZN(n476) );
  AND2_X1 U525 ( .A1(n476), .A2(n551), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U527 ( .A1(n473), .A2(n522), .ZN(n474) );
  XNOR2_X1 U528 ( .A(n474), .B(KEYINPUT103), .ZN(n479) );
  NAND2_X1 U529 ( .A1(n476), .A2(n522), .ZN(n549) );
  NOR2_X1 U530 ( .A1(n529), .A2(n549), .ZN(n538) );
  XNOR2_X1 U531 ( .A(n538), .B(KEYINPUT100), .ZN(n477) );
  INV_X1 U532 ( .A(n527), .ZN(n536) );
  NAND2_X1 U533 ( .A1(n477), .A2(n536), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n491) );
  NAND2_X1 U535 ( .A1(n480), .A2(n491), .ZN(n509) );
  NOR2_X1 U536 ( .A1(n496), .A2(n509), .ZN(n481) );
  XNOR2_X1 U537 ( .A(KEYINPUT104), .B(n481), .ZN(n489) );
  NAND2_X1 U538 ( .A1(n489), .A2(n522), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n489), .A2(n525), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(KEYINPUT106), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .Z(n488) );
  NAND2_X1 U545 ( .A1(n489), .A2(n527), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n489), .A2(n529), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  NAND2_X1 U550 ( .A1(n568), .A2(n491), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT107), .B(n492), .Z(n493) );
  NOR2_X1 U552 ( .A1(n580), .A2(n493), .ZN(n495) );
  XNOR2_X1 U553 ( .A(KEYINPUT108), .B(KEYINPUT37), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(n521) );
  NOR2_X1 U555 ( .A1(n496), .A2(n521), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n497), .B(KEYINPUT38), .ZN(n505) );
  NAND2_X1 U557 ( .A1(n505), .A2(n522), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n505), .A2(n525), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n500), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT110), .ZN(n504) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n502) );
  NAND2_X1 U563 ( .A1(n505), .A2(n527), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1330GAT) );
  XOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT111), .Z(n507) );
  NAND2_X1 U567 ( .A1(n529), .A2(n505), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  INV_X1 U570 ( .A(n563), .ZN(n508) );
  NAND2_X1 U571 ( .A1(n570), .A2(n508), .ZN(n520) );
  NOR2_X1 U572 ( .A1(n520), .A2(n509), .ZN(n516) );
  NAND2_X1 U573 ( .A1(n516), .A2(n522), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n525), .A2(n516), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(KEYINPUT112), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  XOR2_X1 U578 ( .A(G71GAT), .B(KEYINPUT113), .Z(n515) );
  NAND2_X1 U579 ( .A1(n516), .A2(n527), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT114), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U582 ( .A1(n516), .A2(n529), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  XOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT115), .Z(n524) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n530) );
  NAND2_X1 U587 ( .A1(n530), .A2(n522), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n530), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n530), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(KEYINPUT116), .ZN(n534) );
  XOR2_X1 U594 ( .A(KEYINPUT117), .B(KEYINPUT44), .Z(n532) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n546) );
  NOR2_X1 U600 ( .A1(n570), .A2(n546), .ZN(n539) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  NOR2_X1 U602 ( .A1(n546), .A2(n563), .ZN(n543) );
  XOR2_X1 U603 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n541) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n568), .A2(n546), .ZN(n544) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(n544), .Z(n545) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  NOR2_X1 U610 ( .A1(n560), .A2(n546), .ZN(n548) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n535), .A2(n549), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT121), .B(n552), .Z(n559) );
  NOR2_X1 U616 ( .A1(n570), .A2(n559), .ZN(n553) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT122), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n557) );
  NOR2_X1 U621 ( .A1(n563), .A2(n559), .ZN(n556) );
  XOR2_X1 U622 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U623 ( .A1(n568), .A2(n559), .ZN(n558) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NOR2_X1 U627 ( .A1(n570), .A2(n567), .ZN(n562) );
  XOR2_X1 U628 ( .A(G169GAT), .B(n562), .Z(G1348GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n567), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(n566), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n579), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT124), .B(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n579), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

