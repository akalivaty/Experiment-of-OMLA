//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G234));
  NAND2_X1  g026(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n468), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  XOR2_X1   g049(.A(KEYINPUT69), .B(G2105), .Z(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n464), .A3(G137), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n464), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n464), .A2(new_n468), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n480), .A2(G124), .B1(new_n481), .B2(G136), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n475), .C2(G112), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  AND2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NOR2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n469), .B(new_n470), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n475), .A2(new_n464), .A3(new_n491), .A4(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n486), .B2(new_n487), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n490), .B2(new_n492), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT70), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G62), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(new_n515), .B1(G75), .B2(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(KEYINPUT71), .A3(G62), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n513), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(new_n520), .A2(KEYINPUT72), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n524), .A2(G543), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT73), .B(G51), .Z(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n513), .A2(new_n520), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n532), .A2(new_n535), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  XOR2_X1   g116(.A(KEYINPUT74), .B(G52), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n530), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n513), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G651), .B1(new_n534), .B2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  AOI22_X1  g125(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n508), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT75), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n554), .B2(new_n533), .ZN(new_n555));
  INV_X1    g130(.A(G43), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n552), .A2(KEYINPUT75), .B1(new_n556), .B2(new_n529), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND4_X1  g138(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n528), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n566), .A2(new_n567), .A3(new_n508), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n566), .B2(new_n508), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n534), .A2(G91), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(new_n570), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(new_n522), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n516), .A2(new_n517), .ZN(new_n574));
  OAI211_X1 g149(.A(KEYINPUT77), .B(new_n573), .C1(new_n574), .C2(new_n508), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n576), .B1(new_n518), .B2(new_n522), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n575), .A2(new_n577), .ZN(G303));
  OAI21_X1  g153(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  INV_X1    g155(.A(G49), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n579), .B1(new_n580), .B2(new_n533), .C1(new_n529), .C2(new_n581), .ZN(G288));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n511), .B2(new_n512), .ZN(new_n584));
  AND2_X1   g159(.A1(G73), .A2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n511), .B2(new_n512), .ZN(new_n588));
  AND2_X1   g163(.A1(G48), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n520), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n534), .A2(G85), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT78), .B(G47), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n592), .B1(new_n508), .B2(new_n593), .C1(new_n529), .C2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n513), .A2(new_n520), .A3(G92), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n530), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n545), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n597), .B1(new_n598), .B2(new_n610), .ZN(G284));
  AOI21_X1  g186(.A(new_n597), .B1(new_n598), .B2(new_n610), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT80), .Z(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G280));
  INV_X1    g192(.A(new_n608), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT81), .B(G559), .Z(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(G860), .B2(new_n619), .ZN(G148));
  INV_X1    g195(.A(new_n558), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n609), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n619), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n624), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n464), .A2(new_n473), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n480), .A2(G123), .B1(new_n481), .B2(G135), .ZN(new_n632));
  OAI221_X1 g207(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n475), .C2(G111), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n629), .A2(new_n630), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n650), .A2(KEYINPUT83), .A3(new_n638), .ZN(new_n651));
  AOI21_X1  g226(.A(KEYINPUT83), .B1(new_n650), .B2(new_n638), .ZN(new_n652));
  OAI221_X1 g227(.A(G14), .B1(new_n638), .B2(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  INV_X1    g237(.A(new_n655), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n671), .A2(new_n672), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n675), .A3(new_n673), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n678), .B(new_n680), .C1(new_n675), .C2(new_n679), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n669), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n684), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n668), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  NAND3_X1  g269(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT25), .Z(new_n696));
  AOI22_X1  g271(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(new_n475), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n481), .A2(G139), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n702), .B2(G33), .ZN(new_n704));
  INV_X1    g279(.A(G2072), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT90), .Z(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G19), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT88), .Z(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n558), .B2(new_n708), .ZN(new_n711));
  INV_X1    g286(.A(G1341), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n702), .A2(G27), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G164), .B2(new_n702), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n707), .B(new_n713), .C1(G2078), .C2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT24), .ZN(new_n718));
  INV_X1    g293(.A(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n718), .B2(new_n719), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G160), .B2(new_n702), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G2084), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT93), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n618), .A2(new_n708), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G4), .B2(new_n708), .ZN(new_n726));
  INV_X1    g301(.A(G1348), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n702), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n702), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT29), .ZN(new_n730));
  OAI22_X1  g305(.A1(new_n726), .A2(new_n727), .B1(new_n730), .B2(G2090), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n702), .A2(G32), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G141), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT91), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT92), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n480), .A2(G129), .B1(G105), .B2(new_n473), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n732), .B1(new_n740), .B2(new_n702), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT27), .Z(new_n742));
  AOI211_X1 g317(.A(new_n724), .B(new_n731), .C1(new_n742), .C2(G1996), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n708), .A2(G20), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT23), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n615), .B2(new_n708), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G1956), .Z(new_n747));
  OAI211_X1 g322(.A(new_n743), .B(new_n747), .C1(G1996), .C2(new_n742), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n704), .A2(new_n705), .ZN(new_n749));
  NOR2_X1   g324(.A1(G168), .A2(new_n708), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n708), .B2(G21), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT30), .B(G28), .ZN(new_n754));
  OR2_X1    g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n754), .A2(new_n702), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n634), .B2(new_n702), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n722), .B2(G2084), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n751), .A2(new_n752), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n749), .A2(new_n753), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n726), .A2(new_n727), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n708), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n708), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1961), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n730), .A2(G2090), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n702), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  AND3_X1   g343(.A1(new_n471), .A2(new_n464), .A3(G128), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT89), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n475), .A2(G116), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n771), .A2(new_n773), .B1(G140), .B2(new_n481), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(new_n702), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n762), .A2(new_n765), .A3(new_n766), .A4(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n716), .A2(G2078), .ZN(new_n781));
  OR3_X1    g356(.A1(new_n761), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n717), .A2(new_n748), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G6), .A2(G16), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n586), .A2(new_n590), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  INV_X1    g362(.A(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n708), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n708), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1971), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n708), .A2(G23), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n579), .B1(new_n580), .B2(new_n533), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G49), .B2(new_n530), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n793), .B1(new_n795), .B2(new_n708), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n789), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1986), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n702), .A2(G25), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n471), .A2(new_n464), .A3(G119), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT87), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n475), .A2(G107), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n807), .A2(new_n809), .B1(G131), .B2(new_n481), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n804), .B1(new_n812), .B2(new_n702), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n800), .A2(new_n801), .A3(new_n803), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT36), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n783), .A2(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n618), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  INV_X1    g396(.A(G67), .ZN(new_n822));
  INV_X1    g397(.A(G80), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n545), .A2(new_n822), .B1(new_n823), .B2(new_n510), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT95), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n826), .B1(new_n823), .B2(new_n510), .C1(new_n545), .C2(new_n822), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n825), .A2(G651), .A3(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n530), .A2(G55), .B1(G93), .B2(new_n534), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n558), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n555), .B2(new_n557), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n821), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  AOI21_X1  g411(.A(G860), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n832), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(G145));
  NAND2_X1  g416(.A1(new_n775), .A2(new_n501), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n775), .A2(new_n501), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n740), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(new_n739), .A3(new_n842), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n700), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n811), .B(new_n628), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n480), .A2(G130), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT96), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n481), .A2(G142), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n475), .A2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n850), .B(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n845), .A2(new_n847), .A3(new_n701), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n849), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n849), .A2(new_n858), .ZN(new_n862));
  INV_X1    g437(.A(new_n857), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT97), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n866), .A3(new_n863), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n477), .B(new_n634), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n484), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n864), .A2(new_n872), .A3(new_n859), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n871), .A2(KEYINPUT40), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT40), .B1(new_n871), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(G395));
  XNOR2_X1  g454(.A(G290), .B(G288), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  XNOR2_X1  g458(.A(G166), .B(new_n785), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n886), .B1(new_n885), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n834), .B(new_n623), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n894));
  NAND2_X1  g469(.A1(G299), .A2(new_n608), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n568), .A2(new_n569), .B1(G91), .B2(new_n534), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n600), .A2(new_n601), .B1(G651), .B2(new_n606), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n565), .A4(new_n603), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n895), .B2(new_n898), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n894), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n895), .A2(new_n898), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n894), .B1(new_n904), .B2(KEYINPUT41), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n893), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n892), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n908), .B1(new_n893), .B2(new_n907), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n891), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n902), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n900), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n905), .B1(new_n918), .B2(new_n894), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT100), .B1(new_n919), .B2(new_n892), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n890), .A2(new_n920), .A3(new_n911), .A4(new_n909), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT102), .ZN(new_n922));
  INV_X1    g497(.A(new_n912), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n890), .A4(new_n920), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n891), .B(KEYINPUT103), .C1(new_n912), .C2(new_n913), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n916), .A2(new_n922), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(G868), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n832), .A2(new_n609), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(G295));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n929), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  NAND2_X1  g507(.A1(G168), .A2(G171), .ZN(new_n933));
  NAND2_X1  g508(.A1(G286), .A2(G301), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n834), .A2(new_n935), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n831), .A2(new_n833), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n936), .A2(new_n937), .A3(new_n904), .ZN(new_n938));
  INV_X1    g513(.A(new_n936), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n834), .A2(new_n940), .A3(new_n935), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n938), .B1(new_n943), .B2(new_n907), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n885), .A2(new_n887), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n834), .A2(new_n935), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT104), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n937), .A2(new_n940), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n936), .A2(new_n904), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n939), .A2(new_n949), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n952), .A2(new_n953), .B1(new_n954), .B2(new_n918), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n874), .B1(new_n955), .B2(new_n946), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n948), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT43), .B1(new_n944), .B2(new_n946), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n945), .B1(new_n944), .B2(new_n959), .ZN(new_n960));
  AOI211_X1 g535(.A(KEYINPUT105), .B(new_n938), .C1(new_n943), .C2(new_n907), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n874), .B(new_n958), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n932), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n948), .A2(new_n956), .A3(KEYINPUT43), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n874), .B(new_n947), .C1(new_n960), .C2(new_n961), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n966), .B2(new_n932), .ZN(G397));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n504), .B2(G1384), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n476), .A2(G40), .A3(new_n474), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n465), .A2(new_n475), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT106), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n775), .B(new_n778), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n976), .B2(new_n740), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n978), .A2(new_n740), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n812), .A2(new_n814), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT126), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n981), .A2(new_n983), .B1(new_n778), .B2(new_n776), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n811), .B(new_n814), .Z(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n975), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n974), .A2(G1986), .A3(G290), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT48), .ZN(new_n989));
  OAI22_X1  g564(.A1(new_n984), .A2(new_n974), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n979), .A2(new_n740), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n975), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n978), .A2(KEYINPUT127), .A3(KEYINPUT46), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT127), .B1(new_n978), .B2(KEYINPUT46), .ZN(new_n994));
  OAI221_X1 g569(.A(new_n992), .B1(KEYINPUT46), .B2(new_n978), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n995), .A2(KEYINPUT47), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(KEYINPUT47), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT70), .B1(new_n493), .B2(new_n500), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n502), .B(new_n499), .C1(new_n490), .C2(new_n492), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(new_n973), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n504), .A2(G1384), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT113), .B(G2084), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n968), .A2(G1384), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n503), .B2(new_n505), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n969), .A2(new_n973), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n752), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(G168), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G8), .ZN(new_n1016));
  AOI21_X1  g591(.A(G168), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT51), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(new_n1019), .A3(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT122), .B(G1961), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1010), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1026));
  INV_X1    g601(.A(G2078), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n973), .A4(new_n969), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1025), .B1(new_n1028), .B2(KEYINPUT121), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1013), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1027), .A4(new_n1026), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1024), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n973), .B1(new_n504), .B2(new_n1011), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n503), .B2(new_n505), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(KEYINPUT45), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1025), .B1(new_n1037), .B2(G2078), .ZN(new_n1038));
  AOI21_X1  g613(.A(G301), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n575), .A2(G8), .A3(new_n577), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(KEYINPUT55), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n575), .A2(G8), .A3(new_n577), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G2090), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1003), .A2(new_n1049), .A3(new_n1007), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1034), .B1(new_n1002), .B2(new_n968), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT107), .B(G1971), .Z(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(G8), .B(new_n1048), .C1(new_n1050), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1005), .A2(new_n973), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n795), .A2(G1976), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(G8), .A4(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1057), .A2(G8), .A3(new_n1058), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1057), .A2(G8), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT109), .B1(new_n785), .B2(new_n788), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT109), .ZN(new_n1065));
  NOR3_X1   g640(.A1(G305), .A2(new_n1065), .A3(G1981), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT110), .B1(new_n785), .B2(new_n788), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n1069));
  NAND3_X1  g644(.A1(G305), .A2(new_n1069), .A3(G1981), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT111), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1063), .B1(new_n1072), .B2(KEYINPUT49), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT111), .B(new_n1074), .C1(new_n1067), .C2(new_n1071), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1062), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G8), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1052), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1037), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n973), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1006), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT112), .B(new_n973), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1082), .A2(new_n1049), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1077), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1054), .B(new_n1076), .C1(new_n1048), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1018), .A2(new_n1089), .A3(new_n1020), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1022), .A2(new_n1039), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G288), .A2(G1976), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1067), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1076), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1094), .A2(new_n1063), .B1(new_n1095), .B2(new_n1054), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(G8), .A3(G168), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1087), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1097), .ZN(new_n1101));
  OAI21_X1  g676(.A(G8), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1101), .A2(new_n1103), .A3(new_n1054), .A4(new_n1076), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1096), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1091), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1348), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1057), .A2(G2067), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n618), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n565), .B2(KEYINPUT115), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G299), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n896), .B(new_n565), .C1(KEYINPUT115), .C2(KEYINPUT57), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(G2072), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1035), .B(new_n1117), .C1(new_n1036), .C2(KEYINPUT45), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT117), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1051), .A2(new_n1120), .A3(new_n1117), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT114), .B(G1956), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1119), .A2(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1115), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1127), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1109), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1127), .A2(new_n1128), .A3(new_n1113), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1124), .B2(new_n1113), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1124), .A2(new_n1113), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1134), .B1(new_n1137), .B2(new_n1131), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n618), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n976), .B(new_n1035), .C1(new_n1036), .C2(KEYINPUT45), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(new_n712), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1057), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1142), .B1(new_n1147), .B2(new_n558), .ZN(new_n1148));
  AOI211_X1 g723(.A(KEYINPUT59), .B(new_n621), .C1(new_n1143), .C2(new_n1146), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1141), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1139), .A2(new_n608), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1140), .B1(new_n1151), .B2(new_n1109), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1136), .A2(new_n1138), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1038), .A2(G301), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n475), .B1(new_n466), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n465), .A2(KEYINPUT123), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n971), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n969), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT124), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1160), .A2(new_n969), .A3(new_n1163), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n1025), .B(G2078), .C1(new_n501), .C2(new_n1010), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(new_n1023), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1156), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1155), .B1(new_n1039), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1033), .A2(G301), .A3(new_n1038), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n1051), .B2(new_n1027), .ZN(new_n1172));
  OAI21_X1  g747(.A(G171), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1173), .A3(KEYINPUT54), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1170), .A2(new_n1021), .A3(new_n1088), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1133), .A2(new_n1154), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1106), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(G290), .B(G1986), .Z(new_n1180));
  OAI211_X1 g755(.A(new_n981), .B(new_n986), .C1(new_n974), .C2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n998), .B1(new_n1179), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g757(.A1(new_n871), .A2(new_n876), .ZN(new_n1184));
  NOR2_X1   g758(.A1(G227), .A2(new_n462), .ZN(new_n1185));
  AND3_X1   g759(.A1(new_n693), .A2(new_n653), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1187), .A2(new_n966), .ZN(G308));
  AND2_X1   g762(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n1189));
  OAI211_X1 g763(.A(new_n1184), .B(new_n1186), .C1(new_n1189), .C2(new_n964), .ZN(G225));
endmodule


