//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n209), .B1(new_n213), .B2(new_n214), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT70), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT70), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G1), .ZN(new_n247));
  NAND4_X1  g0047(.A1(new_n245), .A2(new_n247), .A3(G13), .A4(G20), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G116), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n210), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n245), .A2(new_n247), .A3(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n248), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n249), .B1(new_n255), .B2(G116), .ZN(new_n256));
  AOI21_X1  g0056(.A(G20), .B1(G33), .B2(G283), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G97), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT92), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT92), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G116), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n250), .A2(new_n210), .B1(G20), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(KEYINPUT20), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT20), .B1(new_n264), .B2(new_n266), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n256), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G179), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G264), .A4(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n273), .A2(new_n275), .A3(G257), .A4(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G303), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT72), .ZN(new_n282));
  INV_X1    g0082(.A(new_n210), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n286), .A2(KEYINPUT72), .A3(new_n210), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n272), .B1(new_n281), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n271), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n286), .A2(new_n210), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT70), .B(G1), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT68), .B(G41), .ZN(new_n295));
  OAI211_X1 g0095(.A(G45), .B(new_n294), .C1(new_n295), .C2(KEYINPUT5), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT5), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G41), .ZN(new_n298));
  OAI211_X1 g0098(.A(G270), .B(new_n293), .C1(new_n296), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT87), .B1(new_n297), .B2(G41), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT87), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT5), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(KEYINPUT68), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT68), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G41), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n297), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n245), .A2(new_n247), .A3(G45), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT86), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT5), .B1(new_n309), .B2(new_n311), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n245), .A2(new_n247), .A3(G45), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT86), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n308), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT91), .B1(new_n300), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n316), .A2(new_n319), .ZN(new_n322));
  INV_X1    g0122(.A(new_n308), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT91), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n299), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n291), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n270), .A2(G169), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n281), .A2(new_n288), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n328), .B1(new_n331), .B2(KEYINPUT21), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n330), .ZN(new_n333));
  INV_X1    g0133(.A(new_n329), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT21), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT93), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT93), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(new_n337), .A3(KEYINPUT21), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n332), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT77), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n244), .B(G274), .C1(new_n286), .C2(new_n210), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT69), .B(G45), .Z(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n295), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n280), .A2(G222), .A3(new_n277), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n280), .A2(G223), .A3(G1698), .ZN(new_n345));
  INV_X1    g0145(.A(G77), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n280), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n347), .B2(new_n288), .ZN(new_n348));
  INV_X1    g0148(.A(G45), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n305), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT71), .B1(new_n294), .B2(new_n350), .ZN(new_n351));
  AND4_X1   g0151(.A1(KEYINPUT71), .A2(new_n350), .A3(new_n245), .A4(new_n247), .ZN(new_n352));
  OAI211_X1 g0152(.A(G226), .B(new_n293), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT73), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT8), .B(G58), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n258), .A2(G20), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G150), .ZN(new_n360));
  NOR2_X1   g0160(.A1(G20), .A2(G33), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n357), .A2(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G50), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n211), .B1(new_n201), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n251), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n248), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n364), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n251), .B1(new_n294), .B2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G50), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT73), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n372), .B1(new_n354), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n356), .B(new_n371), .C1(new_n355), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT76), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n370), .A2(new_n368), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n366), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT9), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(new_n377), .A3(new_n366), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT9), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT10), .ZN(new_n386));
  INV_X1    g0186(.A(G200), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n348), .B2(new_n353), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n348), .A2(new_n353), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(G190), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n386), .B1(new_n385), .B2(new_n390), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n375), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n280), .A2(G232), .A3(new_n277), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n280), .A2(G238), .A3(G1698), .ZN(new_n396));
  INV_X1    g0196(.A(G107), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n395), .B(new_n396), .C1(new_n397), .C2(new_n280), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n288), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n342), .A2(new_n295), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(new_n302), .A3(new_n244), .ZN(new_n401));
  OAI211_X1 g0201(.A(G244), .B(new_n293), .C1(new_n351), .C2(new_n352), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n272), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n357), .B1(KEYINPUT74), .B2(new_n362), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(KEYINPUT74), .B2(new_n362), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT15), .B(G87), .Z(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n358), .B1(G20), .B2(G77), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n252), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n369), .A2(G77), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G77), .B2(new_n248), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n404), .B(new_n413), .C1(G169), .C2(new_n403), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n399), .A2(G190), .A3(new_n401), .A4(new_n402), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n412), .B(new_n415), .C1(new_n403), .C2(new_n387), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT75), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n340), .B1(new_n394), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n420), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n419), .B1(new_n414), .B2(new_n416), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n383), .B1(new_n381), .B2(new_n382), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n390), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT10), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n391), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n425), .A2(KEYINPUT77), .A3(new_n430), .A4(new_n375), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n359), .A2(new_n346), .B1(new_n364), .B2(new_n362), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n215), .A2(new_n211), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n251), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  XOR2_X1   g0235(.A(new_n435), .B(KEYINPUT11), .Z(new_n436));
  NAND3_X1  g0236(.A1(new_n367), .A2(KEYINPUT12), .A3(new_n216), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n369), .A2(G68), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n248), .A2(G68), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n437), .B(new_n438), .C1(KEYINPUT12), .C2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n443));
  INV_X1    g0243(.A(G97), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n280), .A2(new_n277), .ZN(new_n445));
  INV_X1    g0245(.A(G226), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n443), .B1(new_n258), .B2(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n288), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n401), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n293), .B1(new_n351), .B2(new_n352), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(new_n217), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT13), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n343), .B1(new_n447), .B2(new_n288), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n450), .A2(new_n217), .ZN(new_n454));
  XOR2_X1   g0254(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(G179), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n453), .B2(new_n454), .ZN(new_n459));
  OAI21_X1  g0259(.A(G169), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n460), .B2(KEYINPUT14), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT14), .ZN(new_n462));
  INV_X1    g0262(.A(new_n455), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n449), .B2(new_n451), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n456), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n462), .B1(new_n465), .B2(G169), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n442), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(G200), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n452), .A2(G190), .A3(new_n456), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n441), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT82), .ZN(new_n472));
  OAI21_X1  g0272(.A(G232), .B1(new_n286), .B2(new_n210), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n350), .A2(new_n245), .A3(new_n247), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n294), .A2(KEYINPUT71), .A3(new_n350), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n472), .B1(new_n478), .B2(new_n343), .ZN(new_n479));
  INV_X1    g0279(.A(new_n473), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n351), .B2(new_n352), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(KEYINPUT82), .A3(new_n401), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n280), .A2(G226), .A3(G1698), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n280), .A2(G223), .A3(new_n277), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G87), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT81), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n288), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n479), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n387), .ZN(new_n490));
  INV_X1    g0290(.A(G190), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n479), .A2(new_n482), .A3(new_n491), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n248), .A2(new_n357), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n369), .B2(new_n357), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n201), .B1(new_n215), .B2(G58), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n211), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT7), .B1(new_n280), .B2(G20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n273), .A2(new_n275), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT7), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n211), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n503), .A3(new_n215), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n361), .A2(G159), .ZN(new_n505));
  AND2_X1   g0305(.A1(KEYINPUT65), .A2(G68), .ZN(new_n506));
  NOR2_X1   g0306(.A1(KEYINPUT65), .A2(G68), .ZN(new_n507));
  OAI21_X1  g0307(.A(G58), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n202), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(KEYINPUT80), .A3(G20), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n499), .A2(new_n504), .A3(new_n505), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT16), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n252), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n280), .A2(KEYINPUT7), .A3(G20), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n502), .B1(new_n501), .B2(new_n211), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT79), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(G20), .B1(new_n273), .B2(new_n275), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n502), .ZN(new_n519));
  OAI21_X1  g0319(.A(G68), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n211), .B1(new_n508), .B2(new_n202), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(KEYINPUT80), .B1(G159), .B2(new_n361), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n522), .A2(KEYINPUT16), .A3(new_n499), .A4(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n496), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n493), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(G179), .B1(new_n487), .B2(new_n288), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n479), .A2(new_n482), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT83), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n489), .A2(new_n373), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n479), .A2(new_n482), .A3(new_n530), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT18), .B1(new_n536), .B2(new_n526), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n513), .A2(new_n525), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n495), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n479), .A2(new_n482), .A3(new_n530), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n534), .B1(new_n489), .B2(new_n373), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT18), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .A4(new_n532), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n493), .A2(KEYINPUT17), .A3(new_n526), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n529), .A2(new_n537), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n471), .B1(KEYINPUT84), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n545), .A2(KEYINPUT84), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n432), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n270), .B1(new_n333), .B2(G200), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n491), .B2(new_n333), .ZN(new_n550));
  XNOR2_X1  g0350(.A(KEYINPUT89), .B(G87), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT90), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT90), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n554), .A2(new_n556), .B1(new_n211), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n280), .A2(new_n211), .A3(G68), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n359), .A2(new_n444), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(KEYINPUT19), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n251), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n407), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n367), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n255), .A2(G87), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n280), .A2(G244), .A3(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G116), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(new_n568), .C1(new_n445), .C2(new_n217), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n288), .ZN(new_n570));
  INV_X1    g0370(.A(G250), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n292), .B1(new_n318), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n294), .A2(G45), .A3(new_n301), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(KEYINPUT88), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT88), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n318), .A2(new_n571), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(new_n573), .A3(new_n293), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT88), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n574), .B1(new_n288), .B2(new_n569), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G190), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n566), .A2(new_n578), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G283), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n273), .A2(new_n275), .A3(G250), .A4(G1698), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(new_n277), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT4), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n288), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(G257), .B(new_n293), .C1(new_n296), .C2(new_n298), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n324), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  XNOR2_X1  g0395(.A(G97), .B(G107), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT85), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(KEYINPUT6), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n598), .B1(KEYINPUT6), .B2(new_n444), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n596), .ZN(new_n602));
  OAI22_X1  g0402(.A1(new_n602), .A2(new_n211), .B1(new_n346), .B2(new_n362), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n500), .A2(new_n503), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n397), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n251), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n248), .A2(G97), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n255), .B2(G97), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n324), .A2(G190), .A3(new_n592), .A4(new_n593), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n595), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n577), .A2(new_n373), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n583), .A2(new_n272), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n562), .A2(new_n564), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n254), .A2(new_n563), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n317), .A2(new_n318), .A3(new_n298), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n292), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(G257), .B1(new_n322), .B2(new_n323), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(new_n272), .A3(new_n592), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n594), .A2(new_n373), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n606), .A2(new_n608), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n585), .A2(new_n610), .A3(new_n615), .A4(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n273), .A2(new_n275), .A3(new_n211), .A4(G87), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT22), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT22), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n280), .A2(new_n626), .A3(new_n211), .A4(G87), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n568), .A2(G20), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT94), .B1(new_n211), .B2(G107), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT23), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT23), .ZN(new_n632));
  OAI211_X1 g0432(.A(KEYINPUT94), .B(new_n632), .C1(new_n211), .C2(G107), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n629), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT24), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT24), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n628), .A2(new_n637), .A3(new_n634), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n252), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n367), .A2(KEYINPUT25), .A3(new_n397), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT25), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n248), .B2(G107), .ZN(new_n642));
  AOI22_X1  g0442(.A1(G107), .A2(new_n255), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n280), .A2(G257), .A3(G1698), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n280), .A2(G250), .A3(new_n277), .ZN(new_n647));
  NAND2_X1  g0447(.A1(G33), .A2(G294), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n288), .ZN(new_n650));
  OAI211_X1 g0450(.A(G264), .B(new_n293), .C1(new_n296), .C2(new_n298), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n387), .B1(new_n652), .B2(new_n320), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n324), .A2(new_n491), .A3(new_n651), .A4(new_n650), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n645), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n652), .A2(new_n272), .A3(new_n320), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(G169), .B1(new_n652), .B2(new_n320), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n636), .A2(new_n638), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n251), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n658), .A2(new_n659), .B1(new_n661), .B2(new_n643), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT95), .B1(new_n656), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n659), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n664), .A2(new_n657), .B1(new_n639), .B2(new_n644), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n645), .A2(new_n655), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT95), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n623), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  AND4_X1   g0469(.A1(new_n339), .A2(new_n548), .A3(new_n550), .A4(new_n669), .ZN(G372));
  INV_X1    g0470(.A(new_n375), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n467), .A2(new_n414), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n470), .A3(new_n529), .A4(new_n544), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n537), .A2(new_n543), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n430), .B(KEYINPUT97), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n548), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n585), .A3(new_n615), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n578), .A2(KEYINPUT96), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT96), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n577), .A2(new_n683), .A3(G200), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n682), .A2(new_n584), .A3(new_n566), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(new_n679), .A4(new_n615), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n681), .A2(new_n615), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n333), .A2(new_n334), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT21), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n689), .A2(new_n690), .B1(new_n327), .B2(new_n291), .ZN(new_n691));
  INV_X1    g0491(.A(new_n338), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n337), .B1(new_n331), .B2(KEYINPUT21), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n691), .B(new_n665), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n610), .A2(new_n622), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n666), .A3(new_n615), .A4(new_n685), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n688), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n677), .B1(new_n678), .B2(new_n698), .ZN(G369));
  OAI21_X1  g0499(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n211), .A2(G13), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n294), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n271), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n339), .A2(new_n550), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n663), .A2(new_n668), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n645), .B2(new_n706), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n665), .A2(new_n706), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT98), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n711), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n715), .ZN(new_n718));
  INV_X1    g0518(.A(new_n706), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n339), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n718), .A2(new_n720), .B1(new_n662), .B2(new_n706), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n717), .A2(new_n721), .ZN(G399));
  AND3_X1   g0522(.A1(new_n554), .A2(new_n265), .A3(new_n556), .ZN(new_n723));
  INV_X1    g0523(.A(new_n207), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n312), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n214), .B2(new_n726), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT99), .B(KEYINPUT28), .Z(new_n729));
  XNOR2_X1  g0529(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n694), .A2(new_n697), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n615), .B1(new_n680), .B2(KEYINPUT26), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n685), .A2(new_n615), .A3(new_n679), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(new_n733), .B2(KEYINPUT26), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n719), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n698), .A2(KEYINPUT29), .A3(new_n719), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n669), .A2(new_n339), .A3(new_n550), .A4(new_n706), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n594), .A2(new_n577), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n272), .B1(new_n652), .B2(new_n320), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n333), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n321), .A2(new_n326), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n289), .A2(new_n650), .A3(new_n651), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n618), .A3(new_n583), .A4(new_n592), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n577), .A2(new_n290), .A3(new_n652), .ZN(new_n750));
  INV_X1    g0550(.A(new_n594), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n327), .A3(KEYINPUT30), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n744), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n719), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT31), .B1(new_n753), .B2(new_n719), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n739), .B1(new_n740), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n737), .A2(new_n738), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n730), .B1(new_n758), .B2(G1), .ZN(G364));
  INV_X1    g0559(.A(new_n711), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n244), .B1(new_n701), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n725), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G330), .B2(new_n710), .ZN(new_n765));
  INV_X1    g0565(.A(new_n763), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n210), .B1(G20), .B2(new_n373), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n211), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n491), .A3(G200), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n769), .A2(new_n771), .B1(new_n772), .B2(new_n279), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n770), .A2(new_n491), .A3(new_n387), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n280), .B1(new_n775), .B2(G329), .ZN(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n491), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n211), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n776), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(G20), .A2(G179), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT101), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n491), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G200), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n773), .B(new_n780), .C1(G311), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n782), .A2(G190), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n387), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G326), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n783), .A2(new_n387), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT33), .B(G317), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G322), .A2(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n785), .A2(new_n788), .A3(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n280), .B1(new_n772), .B2(new_n551), .C1(new_n397), .C2(new_n771), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT103), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT102), .B(KEYINPUT32), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  OR3_X1    g0597(.A1(new_n774), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n779), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G97), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n796), .B1(new_n774), .B2(new_n797), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G58), .B2(new_n789), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G50), .A2(new_n787), .B1(new_n784), .B2(G77), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n790), .A2(G68), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n795), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n768), .B1(new_n793), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n767), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT100), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n724), .A2(new_n501), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G355), .A2(new_n814), .B1(new_n265), .B2(new_n724), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n242), .A2(new_n349), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n724), .A2(new_n280), .ZN(new_n817));
  INV_X1    g0617(.A(new_n342), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n214), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n815), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n766), .B(new_n807), .C1(new_n813), .C2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT104), .Z(new_n822));
  INV_X1    g0622(.A(new_n810), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n710), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n765), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  OR2_X1    g0626(.A1(new_n414), .A2(new_n719), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n416), .B1(new_n412), .B2(new_n706), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n414), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n698), .B2(new_n719), .ZN(new_n831));
  INV_X1    g0631(.A(new_n830), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n696), .B1(new_n339), .B2(new_n665), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n706), .B(new_n832), .C1(new_n833), .C2(new_n688), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n740), .A2(new_n756), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G330), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n763), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n835), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G137), .A2(new_n787), .B1(new_n790), .B2(G150), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  INV_X1    g0641(.A(new_n789), .ZN(new_n842));
  INV_X1    g0642(.A(new_n784), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n840), .B1(new_n841), .B2(new_n842), .C1(new_n797), .C2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT34), .Z(new_n845));
  INV_X1    g0645(.A(G68), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n364), .A2(new_n772), .B1(new_n771), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT106), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  INV_X1    g0649(.A(G58), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n280), .B1(new_n774), .B2(new_n849), .C1(new_n779), .C2(new_n850), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n845), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G283), .A2(new_n790), .B1(new_n787), .B2(G303), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n265), .B2(new_n843), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT105), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n789), .A2(G294), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n280), .B1(new_n775), .B2(G311), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n857), .A2(new_n800), .ZN(new_n858));
  INV_X1    g0658(.A(new_n772), .ZN(new_n859));
  INV_X1    g0659(.A(new_n771), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n859), .A2(G107), .B1(new_n860), .B2(G87), .ZN(new_n861));
  AND4_X1   g0661(.A1(new_n855), .A2(new_n856), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n767), .B1(new_n852), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n767), .A2(new_n808), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n766), .B1(new_n346), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n863), .B(new_n865), .C1(new_n809), .C2(new_n832), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n839), .A2(new_n866), .ZN(G384));
  INV_X1    g0667(.A(KEYINPUT35), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n265), .B(new_n213), .C1(new_n602), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n602), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n869), .A2(KEYINPUT107), .B1(KEYINPUT35), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(KEYINPUT107), .B2(new_n869), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT36), .Z(new_n873));
  NAND4_X1  g0673(.A1(new_n508), .A2(G50), .A3(G77), .A4(new_n202), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n364), .A2(G68), .ZN(new_n875));
  AOI211_X1 g0675(.A(G13), .B(new_n294), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n674), .A2(new_n705), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n834), .A2(new_n827), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n467), .B(new_n470), .C1(new_n441), .C2(new_n706), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n468), .A2(new_n469), .A3(new_n441), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n460), .A2(KEYINPUT14), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n465), .A2(new_n462), .A3(G169), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(new_n884), .A3(new_n457), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n442), .B(new_n719), .C1(new_n882), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n518), .B1(new_n500), .B2(new_n503), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n524), .B(new_n499), .C1(new_n890), .C2(new_n520), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n512), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n499), .A2(new_n505), .A3(new_n510), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n520), .B1(new_n604), .B2(KEYINPUT79), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n512), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n251), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT108), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n252), .B1(new_n891), .B2(new_n512), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n496), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n705), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n545), .A2(KEYINPUT109), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT109), .B1(new_n545), .B2(new_n903), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n525), .B1(new_n899), .B2(KEYINPUT108), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n896), .A2(new_n897), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n495), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n536), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n909), .A2(new_n910), .B1(new_n526), .B2(new_n493), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n705), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n906), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n539), .A2(new_n541), .A3(new_n532), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n539), .A2(new_n705), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n914), .A2(new_n906), .A3(new_n915), .A4(new_n527), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n904), .A2(new_n905), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n545), .A2(new_n903), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT109), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n545), .A2(KEYINPUT109), .A3(new_n903), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n527), .B1(new_n901), .B2(new_n536), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT37), .B1(new_n926), .B2(new_n903), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n916), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(KEYINPUT38), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n920), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n878), .B1(new_n889), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n545), .A2(new_n539), .A3(new_n705), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n914), .A2(new_n527), .A3(new_n915), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n916), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n918), .B2(new_n919), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n885), .A2(new_n442), .A3(new_n706), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n920), .A2(new_n929), .A3(KEYINPUT39), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n931), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n548), .B1(new_n737), .B2(new_n738), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n677), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n945), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n830), .B1(new_n881), .B2(new_n886), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n836), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT40), .B1(new_n930), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n836), .A2(new_n949), .A3(KEYINPUT40), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n951), .B1(new_n938), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n548), .A2(new_n836), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n739), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n294), .B2(new_n701), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n948), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n877), .B1(new_n958), .B2(new_n959), .ZN(G367));
  NAND2_X1  g0760(.A1(new_n621), .A2(new_n719), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n695), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n679), .A2(new_n719), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n718), .A2(new_n720), .A3(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT42), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n622), .B1(new_n962), .B2(new_n665), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n706), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(KEYINPUT42), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n566), .A2(new_n706), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n685), .A3(new_n615), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n615), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT110), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n970), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n976), .B1(new_n970), .B2(new_n978), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n964), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n717), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n981), .B(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n725), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n718), .B(new_n720), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(new_n711), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n711), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n758), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n721), .A2(new_n995), .A3(new_n964), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n721), .B2(new_n964), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT112), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n996), .A2(new_n997), .B1(new_n716), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n721), .A2(new_n964), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n716), .A2(new_n998), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1004), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n999), .A2(new_n1006), .A3(new_n1002), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n994), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n987), .B1(new_n1008), .B2(new_n992), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n985), .B1(new_n1009), .B2(new_n761), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n813), .B1(new_n207), .B2(new_n563), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n817), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n234), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n763), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G283), .A2(new_n784), .B1(new_n790), .B2(G294), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n787), .ZN(new_n1016));
  XOR2_X1   g0816(.A(KEYINPUT113), .B(G311), .Z(new_n1017));
  OAI221_X1 g0817(.A(new_n1015), .B1(new_n279), .B2(new_n842), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n859), .A2(G116), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT46), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n771), .A2(new_n444), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n280), .B(new_n1021), .C1(G317), .C2(new_n775), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(new_n397), .C2(new_n779), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n790), .A2(G159), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n860), .A2(G77), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(KEYINPUT114), .B(G137), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n501), .B1(new_n775), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n799), .A2(G68), .B1(new_n859), .B2(G58), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G50), .A2(new_n784), .B1(new_n789), .B2(G150), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n841), .B2(new_n1016), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1018), .A2(new_n1023), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1014), .B1(new_n1033), .B2(new_n767), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n974), .A2(new_n823), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1010), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(G387));
  INV_X1    g0839(.A(new_n991), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n713), .A2(new_n715), .A3(new_n810), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n817), .B1(new_n230), .B2(new_n342), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n814), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n723), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n357), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n723), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1044), .A2(new_n1048), .B1(new_n397), .B2(new_n724), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n763), .B1(new_n1049), .B2(new_n812), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n787), .A2(G159), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT115), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n789), .A2(G50), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n563), .A2(new_n779), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n280), .B1(new_n774), .B2(new_n360), .C1(new_n444), .C2(new_n771), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(G77), .C2(new_n859), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n357), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G68), .A2(new_n784), .B1(new_n790), .B2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1052), .A2(new_n1053), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G303), .A2(new_n784), .B1(new_n789), .B2(G317), .ZN(new_n1060));
  INV_X1    g0860(.A(G322), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n790), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1016), .C1(new_n1062), .C2(new_n1017), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n779), .A2(new_n769), .B1(new_n772), .B2(new_n777), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n280), .B1(new_n775), .B2(G326), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n265), .C2(new_n771), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT49), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1059), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1050), .B1(new_n1072), .B2(new_n767), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1040), .A2(new_n762), .B1(new_n1041), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n994), .A2(new_n725), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1040), .A2(new_n758), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(G393));
  AOI21_X1  g0877(.A(new_n761), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n982), .A2(new_n810), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n239), .A2(new_n1012), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n813), .B1(new_n444), .B2(new_n207), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n763), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n779), .A2(new_n346), .ZN(new_n1083));
  INV_X1    g0883(.A(G87), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n280), .B1(new_n774), .B2(new_n841), .C1(new_n1084), .C2(new_n771), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(new_n215), .C2(new_n859), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n364), .B2(new_n1062), .C1(new_n357), .C2(new_n843), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G150), .A2(new_n787), .B1(new_n789), .B2(G159), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT51), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G311), .A2(new_n789), .B1(new_n787), .B2(G317), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n774), .A2(new_n1061), .B1(new_n772), .B2(new_n769), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n784), .A2(G294), .B1(KEYINPUT116), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n501), .B1(new_n771), .B2(new_n397), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G116), .B2(new_n799), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n790), .A2(G303), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1092), .A2(KEYINPUT116), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1087), .A2(new_n1089), .B1(new_n1091), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1082), .B1(new_n1099), .B2(new_n767), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1078), .B1(new_n1079), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1007), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1006), .B1(new_n999), .B2(new_n1002), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n993), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1005), .A2(new_n994), .A3(new_n1007), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n725), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1101), .A2(new_n1106), .ZN(G390));
  NAND3_X1  g0907(.A1(new_n757), .A2(new_n832), .A3(new_n887), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n942), .B1(new_n879), .B2(new_n887), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n940), .B2(new_n943), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n827), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n735), .B2(new_n829), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n938), .B(new_n941), .C1(new_n1113), .C2(new_n888), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1109), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n940), .A2(new_n943), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1110), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n1114), .A3(new_n1108), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n548), .A2(new_n757), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n946), .A2(new_n677), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n887), .B1(new_n757), .B2(new_n832), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n879), .B1(new_n1109), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1124), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n1113), .A3(new_n1108), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1121), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1116), .A2(new_n1120), .A3(new_n1128), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n725), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1116), .A2(new_n1120), .A3(new_n762), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1117), .A2(new_n808), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n864), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n763), .B1(new_n1057), .B2(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n501), .B1(new_n774), .B2(new_n777), .C1(new_n846), .C2(new_n771), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1083), .B(new_n1137), .C1(G87), .C2(new_n859), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n784), .A2(G97), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n790), .A2(G107), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G116), .A2(new_n789), .B1(new_n787), .B2(G283), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G128), .A2(new_n787), .B1(new_n789), .B2(G132), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT118), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n799), .A2(G159), .B1(new_n775), .B2(G125), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT53), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n772), .A2(new_n360), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n790), .A2(new_n1026), .B1(new_n784), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n280), .B1(new_n771), .B2(new_n364), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT117), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1149), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1142), .B1(new_n1144), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1136), .B1(new_n1156), .B2(new_n767), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1134), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1132), .A2(new_n1133), .A3(new_n1158), .ZN(G378));
  NAND2_X1  g0959(.A1(new_n676), .A2(new_n375), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n902), .B1(new_n381), .B2(new_n382), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1161), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n676), .A2(new_n375), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n918), .A2(new_n919), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT38), .B1(new_n925), .B2(new_n928), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n950), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT40), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n739), .B1(new_n952), .B2(new_n938), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT121), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n923), .A2(new_n924), .B1(new_n916), .B2(new_n927), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n936), .B1(new_n1175), .B2(KEYINPUT38), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n836), .A2(new_n949), .A3(KEYINPUT40), .ZN(new_n1177));
  OAI21_X1  g0977(.A(G330), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT121), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n951), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1167), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n951), .B2(new_n1178), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1166), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1165), .B(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1181), .A2(new_n945), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1123), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1131), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n945), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n836), .A2(new_n949), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n920), .B2(new_n929), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1173), .B(KEYINPUT121), .C1(KEYINPUT40), .C2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1184), .B1(new_n1182), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1167), .B1(new_n1194), .B2(new_n1179), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1189), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1186), .A2(new_n1188), .A3(new_n1196), .A4(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n945), .A2(KEYINPUT122), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1181), .A2(new_n1198), .A3(new_n1185), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT122), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n931), .B2(new_n944), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1199), .A2(new_n1202), .B1(new_n1187), .B2(new_n1131), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n725), .B(new_n1197), .C1(new_n1203), .C2(KEYINPUT57), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1167), .A2(new_n808), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n779), .A2(new_n360), .B1(new_n772), .B2(new_n1150), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G125), .A2(new_n787), .B1(new_n789), .B2(G128), .ZN(new_n1207));
  INV_X1    g1007(.A(G137), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1207), .B1(new_n1208), .B2(new_n843), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1206), .B(new_n1209), .C1(G132), .C2(new_n790), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G33), .B(G41), .C1(new_n775), .C2(G124), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n797), .B2(new_n771), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT120), .Z(new_n1216));
  NAND3_X1  g1016(.A1(new_n1212), .A2(new_n1213), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n787), .A2(G116), .B1(G68), .B2(new_n799), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT119), .Z(new_n1219));
  NAND2_X1  g1019(.A1(new_n859), .A2(G77), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n860), .A2(G58), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n775), .A2(G283), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n312), .A2(new_n280), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G97), .B2(new_n790), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n397), .B2(new_n842), .C1(new_n563), .C2(new_n843), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT58), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n364), .B1(G33), .B2(G41), .C1(new_n312), .C2(new_n280), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1227), .A2(KEYINPUT58), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1217), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n767), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n864), .A2(new_n364), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1205), .A2(new_n763), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1236), .B2(new_n762), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1204), .A2(new_n1237), .ZN(G375));
  NAND3_X1  g1038(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1129), .A2(new_n1239), .A3(new_n987), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n762), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n763), .B1(G68), .B2(new_n1135), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1025), .A2(new_n501), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT123), .Z(new_n1245));
  NOR2_X1   g1045(.A1(new_n772), .A2(new_n444), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1246), .B(new_n1054), .C1(G303), .C2(new_n775), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(new_n769), .C2(new_n842), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G107), .A2(new_n784), .B1(new_n790), .B2(G116), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n777), .B2(new_n1016), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n789), .A2(new_n1026), .B1(new_n790), .B2(new_n1151), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n849), .B2(new_n1016), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n784), .A2(G150), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n501), .B1(new_n775), .B2(G128), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n799), .A2(G50), .B1(new_n859), .B2(G159), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1221), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1248), .A2(new_n1250), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1243), .B1(new_n1257), .B2(new_n767), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n887), .B2(new_n809), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1242), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1240), .A2(new_n1261), .ZN(G381));
  OR3_X1    g1062(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(G378), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(new_n1204), .A4(new_n1237), .ZN(G407));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G375), .C2(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT127), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1010), .B2(new_n1037), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1104), .A2(new_n758), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n762), .B1(new_n1274), .B2(new_n987), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G390), .B(new_n1036), .C1(new_n1275), .C2(new_n985), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(G393), .B(new_n825), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1273), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1268), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT60), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1239), .B1(new_n1128), .B2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .A4(KEYINPUT60), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1284), .A2(new_n725), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(G384), .A3(new_n1261), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1286), .B2(new_n1261), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1204), .A2(G378), .A3(new_n1237), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1186), .A2(new_n1196), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT124), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1186), .A2(new_n1196), .A3(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n762), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1235), .B1(new_n1203), .B2(new_n987), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G378), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1281), .B(new_n1290), .C1(new_n1291), .C2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1186), .A2(new_n1294), .A3(new_n1196), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1294), .B1(new_n1186), .B2(new_n1196), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n761), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1236), .A2(new_n987), .A3(new_n1188), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1234), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1265), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1204), .A2(G378), .A3(new_n1237), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1268), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1268), .A2(G2897), .ZN(new_n1310));
  INV_X1    g1110(.A(G384), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1311), .B1(new_n1312), .B2(new_n1260), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1287), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1310), .B1(new_n1314), .B2(KEYINPUT125), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT125), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1310), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n1316), .B(new_n1317), .C1(new_n1313), .C2(new_n1287), .ZN(new_n1318));
  OAI22_X1  g1118(.A1(new_n1315), .A2(new_n1318), .B1(KEYINPUT125), .B2(new_n1314), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1301), .B1(new_n1309), .B2(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1300), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1280), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT126), .B1(new_n1309), .B2(new_n1319), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1281), .B1(new_n1291), .B2(new_n1298), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1317), .B1(new_n1290), .B2(new_n1316), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1314), .A2(KEYINPUT125), .A3(new_n1310), .ZN(new_n1327));
  AOI22_X1  g1127(.A1(new_n1326), .A2(new_n1327), .B1(new_n1316), .B2(new_n1290), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1325), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1299), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1324), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1280), .B(new_n1301), .C1(new_n1299), .C2(new_n1331), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1271), .B1(new_n1323), .B2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1328), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1309), .A2(new_n1338), .A3(new_n1290), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1322), .A3(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1280), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1342), .B(KEYINPUT127), .C1(new_n1334), .C2(new_n1333), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1336), .A2(new_n1343), .ZN(G405));
  XNOR2_X1  g1144(.A(G375), .B(G378), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1290), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1346), .B(new_n1280), .ZN(G402));
endmodule


