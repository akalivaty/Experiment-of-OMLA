//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n542, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT65), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n463), .A2(new_n468), .A3(G137), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT64), .Z(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  XOR2_X1   g051(.A(KEYINPUT3), .B(G2104), .Z(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n463), .A2(new_n468), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n469), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR4_X1   g066(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n491), .A4(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(new_n468), .A3(G138), .A4(new_n469), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n496), .B(KEYINPUT67), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n463), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n494), .A2(new_n499), .ZN(G164));
  AND2_X1   g075(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n502));
  OAI21_X1  g077(.A(G651), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  OAI211_X1 g082(.A(KEYINPUT69), .B(G651), .C1(new_n501), .C2(new_n502), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n505), .A2(G543), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n505), .A2(new_n511), .A3(new_n507), .A4(new_n508), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT70), .B(G88), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  NAND4_X1  g092(.A1(new_n505), .A2(G89), .A3(new_n507), .A4(new_n508), .ZN(new_n518));
  NAND2_X1  g093(.A1(G63), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n511), .ZN(new_n521));
  INV_X1    g096(.A(new_n509), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n523), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  AOI22_X1  g103(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n506), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n530), .B1(new_n509), .B2(new_n531), .C1(new_n532), .C2(new_n514), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  INV_X1    g109(.A(G43), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n509), .A2(new_n535), .B1(new_n506), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n514), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  AND3_X1   g116(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G36), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G188));
  AOI22_X1  g121(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n506), .ZN(new_n548));
  INV_X1    g123(.A(new_n514), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G91), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n509), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(new_n553), .B2(G53), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  NOR4_X1   g130(.A1(new_n509), .A2(new_n552), .A3(KEYINPUT9), .A4(new_n555), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n548), .B(new_n550), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT73), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n559), .A2(KEYINPUT72), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n553), .A2(new_n551), .A3(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n563), .A2(new_n564), .A3(new_n548), .A4(new_n550), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n558), .A2(new_n565), .ZN(G299));
  OR2_X1    g141(.A1(new_n513), .A2(new_n516), .ZN(G303));
  OAI21_X1  g142(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n568));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n514), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G49), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n509), .A2(new_n571), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n570), .A2(new_n572), .ZN(G288));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n509), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n549), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XOR2_X1   g153(.A(KEYINPUT5), .B(G543), .Z(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(KEYINPUT74), .A3(G651), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n506), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n576), .A2(new_n577), .A3(new_n586), .ZN(G305));
  AND2_X1   g162(.A1(new_n549), .A2(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n509), .A2(new_n589), .B1(new_n506), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n549), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n514), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n579), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n595), .A2(new_n598), .B1(G651), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n522), .A2(G54), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n594), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n594), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  MUX2_X1   g182(.A(G286), .B(G299), .S(new_n607), .Z(G280));
  XOR2_X1   g183(.A(G280), .B(KEYINPUT75), .Z(G297));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n604), .B1(new_n610), .B2(G860), .ZN(G148));
  NOR2_X1   g186(.A1(new_n540), .A2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n595), .A2(new_n598), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n601), .A2(G651), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n613), .A2(new_n610), .A3(new_n603), .A4(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n602), .A2(KEYINPUT76), .A3(new_n610), .A4(new_n603), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G868), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT77), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n483), .A2(G123), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT78), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(KEYINPUT79), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(KEYINPUT79), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n627), .C1(G111), .C2(new_n469), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n485), .A2(G135), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n477), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n471), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n632), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2443), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(KEYINPUT81), .ZN(new_n662));
  INV_X1    g237(.A(new_n658), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n657), .A3(new_n665), .ZN(new_n666));
  OAI221_X1 g241(.A(new_n660), .B1(new_n661), .B2(new_n662), .C1(new_n664), .C2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n631), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT83), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT82), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n673), .A2(new_n676), .A3(new_n680), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT87), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n688), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G35), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n695), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT29), .Z(new_n698));
  INV_X1    g273(.A(G2090), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT99), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n483), .A2(G129), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n485), .A2(G141), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT97), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n471), .A2(G105), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n702), .A2(new_n703), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G32), .B(new_n708), .S(G29), .Z(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT27), .B(G1996), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n695), .A2(G26), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n483), .A2(G128), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n485), .A2(G140), .ZN(new_n716));
  OR2_X1    g291(.A1(G104), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(new_n695), .ZN(new_n721));
  INV_X1    g296(.A(G2067), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G19), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n540), .B2(new_n724), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(G1341), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n711), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G168), .A2(new_n724), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n724), .B2(G21), .ZN(new_n730));
  INV_X1    g305(.A(G1966), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n695), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n695), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n733), .C1(G2078), .C2(new_n735), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n701), .A2(new_n728), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n695), .B1(new_n738), .B2(G28), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(KEYINPUT98), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(KEYINPUT98), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n740), .B(new_n741), .C1(new_n738), .C2(G28), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n630), .A2(new_n695), .ZN(new_n743));
  INV_X1    g318(.A(G2072), .ZN(new_n744));
  OR2_X1    g319(.A1(G29), .A2(G33), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n485), .A2(G139), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT25), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n633), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n746), .B(new_n749), .C1(new_n469), .C2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(new_n695), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n742), .B(new_n743), .C1(new_n744), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G5), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G171), .B2(G16), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G1961), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n735), .A2(G2078), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n752), .A2(new_n744), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT96), .Z(new_n759));
  NAND4_X1  g334(.A1(new_n753), .A2(new_n756), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  OR2_X1    g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT24), .A2(G34), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n762), .A2(new_n695), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G160), .B2(new_n695), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT95), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n724), .A2(G4), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n604), .B2(new_n724), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G1348), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n761), .A2(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n698), .A2(new_n699), .B1(new_n766), .B2(new_n761), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n760), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n737), .B(new_n774), .C1(G1961), .C2(new_n755), .ZN(new_n775));
  AND3_X1   g350(.A1(new_n724), .A2(KEYINPUT23), .A3(G20), .ZN(new_n776));
  AOI21_X1  g351(.A(KEYINPUT23), .B1(new_n724), .B2(G20), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n776), .B(new_n777), .C1(G299), .C2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1956), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT31), .B(G11), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n695), .A2(G25), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n483), .A2(G119), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n485), .A2(G131), .ZN(new_n785));
  OR2_X1    g360(.A1(G95), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(new_n695), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT35), .B(G1991), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n790), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n724), .A2(G24), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n592), .B2(new_n724), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT88), .B(G1986), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n724), .A2(G23), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n570), .A2(new_n572), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n724), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT33), .Z(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G1976), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(G1976), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n724), .A2(G6), .ZN(new_n804));
  INV_X1    g379(.A(G305), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n724), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT32), .B(G1981), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT90), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n724), .A2(G22), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G166), .B2(new_n724), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT91), .B(G1971), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n802), .A2(new_n803), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n793), .B(new_n797), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT92), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n815), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n818), .B1(new_n817), .B2(new_n819), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n781), .B(new_n782), .C1(new_n820), .C2(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  NAND2_X1  g398(.A1(G80), .A2(G543), .ZN(new_n824));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n579), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G651), .ZN(new_n827));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n509), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n514), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(G860), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n604), .A2(G559), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n559), .A2(G93), .A3(new_n511), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT68), .B(KEYINPUT6), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT69), .B1(new_n838), .B2(G651), .ZN(new_n839));
  INV_X1    g414(.A(new_n508), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n841), .A2(G55), .A3(G543), .A4(new_n507), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n837), .A2(new_n842), .A3(new_n843), .A4(new_n827), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT100), .B1(new_n829), .B2(new_n831), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n540), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n844), .A2(new_n845), .A3(new_n540), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n836), .B(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n833), .B1(new_n851), .B2(G860), .ZN(G145));
  NAND2_X1  g427(.A1(new_n483), .A2(G130), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n485), .A2(G142), .ZN(new_n854));
  NOR2_X1   g429(.A1(G106), .A2(G2105), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(new_n469), .B2(G118), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n853), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(new_n635), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n789), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n708), .B(new_n719), .ZN(new_n860));
  XNOR2_X1  g435(.A(G164), .B(KEYINPUT101), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n751), .B(KEYINPUT102), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n751), .A2(KEYINPUT102), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n859), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT103), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n864), .A2(new_n866), .A3(new_n859), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(new_n859), .C1(new_n864), .C2(new_n866), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n630), .B(new_n480), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n489), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n867), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n558), .A2(new_n565), .A3(new_n604), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n604), .B1(new_n558), .B2(new_n565), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n604), .ZN(new_n884));
  NAND2_X1  g459(.A1(G299), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n558), .A2(new_n565), .A3(new_n604), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n844), .A2(new_n845), .A3(new_n540), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n540), .B1(new_n844), .B2(new_n845), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT104), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n848), .B2(new_n849), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n890), .A2(new_n892), .A3(new_n619), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT104), .B1(new_n888), .B2(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n848), .A2(new_n891), .A3(new_n849), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n894), .A2(new_n895), .B1(new_n617), .B2(new_n618), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n883), .B(new_n887), .C1(new_n893), .C2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n881), .A2(new_n882), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n619), .B1(new_n890), .B2(new_n892), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n894), .A2(new_n895), .A3(new_n617), .A4(new_n618), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n904), .A2(KEYINPUT105), .A3(new_n887), .A4(new_n883), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n899), .A2(new_n908), .A3(new_n903), .A4(new_n905), .ZN(new_n909));
  XNOR2_X1  g484(.A(G288), .B(G166), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n592), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(new_n799), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G290), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(G305), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n907), .A2(new_n909), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n907), .B2(new_n909), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n917), .A2(new_n918), .A3(new_n607), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n829), .A2(new_n831), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(G868), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT106), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n918), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n907), .A2(new_n909), .A3(new_n916), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(G868), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n927), .ZN(G295));
  NAND2_X1  g503(.A1(new_n922), .A2(new_n927), .ZN(G331));
  NAND4_X1  g504(.A1(G301), .A2(new_n521), .A3(new_n523), .A4(new_n526), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(G286), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n930), .B(new_n931), .C1(new_n888), .C2(new_n889), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n930), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n849), .A3(new_n848), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n900), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n883), .A2(new_n887), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n932), .A3(KEYINPUT107), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(KEYINPUT107), .B2(new_n932), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n915), .B(new_n935), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n916), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n883), .A2(new_n887), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n934), .A2(new_n932), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n946), .A2(new_n947), .B1(new_n900), .B2(new_n938), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n939), .B(new_n940), .C1(new_n948), .C2(new_n915), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n949), .B2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n941), .A2(KEYINPUT108), .A3(new_n954), .A4(new_n943), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n943), .A2(new_n939), .A3(new_n954), .A4(new_n940), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n952), .B1(new_n961), .B2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n708), .B(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n719), .B(new_n722), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n791), .B2(new_n788), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n789), .A2(new_n792), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1986), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n592), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT110), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n971), .B(new_n974), .C1(new_n972), .C2(new_n592), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n494), .B2(new_n499), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n473), .A2(G40), .A3(new_n479), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n980), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT45), .B(new_n976), .C1(new_n494), .C2(new_n499), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1971), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n989), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n980), .B1(new_n991), .B2(KEYINPUT112), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n977), .A2(new_n994), .A3(KEYINPUT50), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n988), .B(new_n990), .C1(new_n996), .C2(G2090), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n998));
  NAND2_X1  g573(.A1(G303), .A2(G8), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI211_X1 g576(.A(KEYINPUT113), .B(KEYINPUT55), .C1(G303), .C2(G8), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n997), .A2(G8), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1976), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G288), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1009), .A2(KEYINPUT117), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT117), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n799), .A2(G1976), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT114), .B(G8), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1013), .B(new_n1014), .C1(new_n980), .C2(new_n977), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1981), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n576), .A2(new_n577), .A3(new_n1017), .A4(new_n586), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT118), .B(G86), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n514), .A2(new_n1019), .B1(new_n506), .B2(new_n584), .ZN(new_n1020));
  OAI21_X1  g595(.A(G1981), .B1(new_n1020), .B2(new_n575), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT49), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n977), .A2(new_n980), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1014), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1022), .A2(new_n1023), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1025), .A2(new_n1028), .A3(KEYINPUT120), .A4(new_n1030), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1016), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n993), .A2(new_n983), .A3(new_n991), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1037), .A2(new_n699), .B1(new_n986), .B2(new_n985), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1005), .B1(new_n1038), .B2(new_n1027), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1026), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1040), .A2(KEYINPUT115), .A3(new_n1014), .A4(new_n1013), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1015), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1043), .A3(KEYINPUT52), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT116), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1041), .A2(new_n1043), .A3(new_n1046), .A4(KEYINPUT52), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1007), .A2(new_n1035), .A3(new_n1039), .A4(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT56), .B(G2072), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n979), .A2(new_n983), .A3(new_n984), .A4(new_n1050), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1051), .A2(KEYINPUT123), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1036), .A2(new_n779), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(KEYINPUT123), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n557), .B(KEYINPUT57), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n996), .A2(new_n770), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1026), .B(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G2067), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1057), .B1(new_n1062), .B2(new_n884), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1056), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1062), .A2(KEYINPUT60), .A3(new_n884), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n996), .A2(new_n770), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(KEYINPUT60), .C1(G2067), .C2(new_n1060), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1074), .A3(new_n604), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1057), .A2(new_n1065), .A3(KEYINPUT61), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1069), .A2(new_n1070), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT58), .B(G1341), .Z(new_n1078));
  NAND2_X1  g653(.A1(new_n1060), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n985), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n964), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n847), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT59), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1066), .B1(new_n1077), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n992), .A2(new_n761), .A3(new_n993), .A4(new_n995), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n985), .A2(new_n731), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1027), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G168), .A2(new_n1027), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1087), .A2(KEYINPUT51), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G8), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1088), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1090), .A2(new_n1093), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G2078), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n1080), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1961), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n996), .ZN(new_n1099));
  XOR2_X1   g674(.A(G301), .B(KEYINPUT54), .Z(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n478), .B(KEYINPUT125), .Z(new_n1102));
  AOI211_X1 g677(.A(new_n1101), .B(G2078), .C1(new_n1102), .C2(G2105), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n473), .A2(G40), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(new_n979), .A3(new_n984), .A4(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1099), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1080), .A2(KEYINPUT53), .A3(new_n1096), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1100), .B1(new_n1099), .B2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1095), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1084), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1095), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1094), .A2(new_n1088), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1093), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(new_n1089), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT62), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1099), .A2(new_n1107), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1112), .A2(G171), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1049), .B1(new_n1110), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1007), .A2(new_n1035), .A3(new_n1048), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1087), .A2(G168), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(KEYINPUT122), .A3(new_n1039), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1049), .B2(new_n1121), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n997), .A2(G8), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1005), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1120), .A2(KEYINPUT63), .A3(new_n1122), .A4(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n799), .A2(new_n1008), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1018), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1028), .B(KEYINPUT121), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1035), .A2(new_n1048), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1007), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n982), .B1(new_n1119), .B2(new_n1139), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n967), .A2(new_n969), .B1(G2067), .B2(new_n719), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1141), .A2(new_n981), .ZN(new_n1142));
  INV_X1    g717(.A(new_n966), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n981), .B1(new_n1143), .B2(new_n708), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT46), .ZN(new_n1145));
  INV_X1    g720(.A(new_n981), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(G1996), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n981), .A2(KEYINPUT46), .A3(new_n964), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT47), .Z(new_n1150));
  NOR2_X1   g725(.A1(new_n974), .A2(new_n1146), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n970), .A2(new_n981), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n1142), .B(new_n1150), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1140), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g731(.A(G319), .ZN(new_n1158));
  OR2_X1    g732(.A1(G227), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OR2_X1    g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1162));
  AND3_X1   g736(.A1(new_n693), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g737(.A(G401), .B1(new_n875), .B2(new_n877), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n1163), .A2(new_n950), .A3(new_n1164), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


