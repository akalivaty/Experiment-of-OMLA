//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT68), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT69), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G101), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(G125), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n476), .B1(new_n484), .B2(new_n485), .ZN(G160));
  AOI21_X1  g061(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n487));
  AOI22_X1  g062(.A1(G124), .A2(new_n487), .B1(new_n473), .B2(G136), .ZN(new_n488));
  INV_X1    g063(.A(G100), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n489), .A2(new_n467), .A3(KEYINPUT72), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT72), .B1(new_n489), .B2(new_n467), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G112), .B2(new_n467), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT73), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n467), .B2(G114), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT74), .A3(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(G126), .A2(new_n487), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT76), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n504), .B(new_n505), .C1(new_n478), .C2(new_n477), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(KEYINPUT75), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n467), .A2(G138), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n471), .B2(new_n472), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n511), .B2(new_n505), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n504), .B(new_n509), .C1(new_n478), .C2(new_n477), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT4), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n502), .B(new_n508), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  OR2_X1    g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G50), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n522), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n526), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n531), .B1(new_n532), .B2(new_n524), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n521), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n524), .A2(new_n543), .B1(new_n526), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n521), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n524), .A2(new_n549), .B1(new_n526), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(KEYINPUT78), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(KEYINPUT78), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT79), .Z(G188));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n526), .A2(KEYINPUT9), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n526), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(new_n519), .ZN(new_n568));
  XNOR2_X1  g143(.A(KEYINPUT80), .B(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n524), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n570), .A2(G651), .B1(new_n571), .B2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n566), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  OAI21_X1  g149(.A(KEYINPUT81), .B1(new_n537), .B2(new_n539), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n535), .A2(new_n536), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n531), .B1(new_n524), .B2(new_n532), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(new_n579), .A3(new_n538), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n526), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n519), .A2(new_n523), .A3(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT82), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n526), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G49), .ZN(new_n590));
  INV_X1    g165(.A(new_n587), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n584), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n588), .A2(new_n593), .ZN(G288));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  INV_X1    g170(.A(G48), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n524), .A2(new_n595), .B1(new_n526), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n517), .B2(new_n518), .ZN(new_n599));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n521), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  INV_X1    g182(.A(G47), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n524), .A2(new_n607), .B1(new_n526), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n519), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n521), .B1(new_n613), .B2(KEYINPUT83), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(KEYINPUT83), .B2(new_n613), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n519), .A2(new_n523), .A3(G92), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n589), .A2(G54), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n612), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n612), .B1(new_n620), .B2(G868), .ZN(G321));
  NOR2_X1   g197(.A1(G299), .A2(G868), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n581), .B2(G868), .ZN(G297));
  AOI21_X1  g199(.A(new_n623), .B1(new_n581), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n620), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n620), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n471), .A2(new_n472), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n464), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT84), .B(G2100), .Z(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n473), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n487), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n467), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n637), .A2(new_n638), .A3(new_n644), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT17), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT85), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n668), .B(new_n665), .C1(new_n661), .C2(new_n663), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n661), .A3(new_n663), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n681), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n678), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(KEYINPUT88), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(KEYINPUT88), .ZN(new_n688));
  AOI211_X1 g263(.A(new_n683), .B(new_n685), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(G1971), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G6), .A2(G16), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n603), .B2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n697), .A2(G23), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n586), .A2(new_n587), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n697), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n701), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT90), .B(G29), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT91), .ZN(new_n720));
  AOI22_X1  g295(.A1(G119), .A2(new_n487), .B1(new_n473), .B2(G131), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n717), .B1(new_n722), .B2(new_n716), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n697), .A2(G24), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n610), .B2(new_n697), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1986), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n712), .A2(new_n713), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n714), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT36), .Z(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G33), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n738));
  NAND3_X1  g313(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n473), .A2(G139), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n632), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n740), .B(new_n741), .C1(new_n467), .C2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT97), .Z(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2072), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n697), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n697), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT102), .Z(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n736), .A2(G32), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n473), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT26), .Z(new_n754));
  INV_X1    g329(.A(G129), .ZN(new_n755));
  INV_X1    g330(.A(new_n487), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n752), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(new_n736), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT100), .Z(new_n760));
  OAI221_X1 g335(.A(new_n746), .B1(G1961), .B2(new_n749), .C1(new_n750), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n716), .A2(G35), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n716), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G2090), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n620), .A2(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G4), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(G1348), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n697), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT23), .Z(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  NOR2_X1   g348(.A1(G164), .A2(new_n715), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G27), .B2(new_n715), .ZN(new_n775));
  INV_X1    g350(.A(G2078), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n769), .A2(new_n773), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n697), .A2(G21), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G168), .B2(new_n697), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n760), .A2(new_n750), .B1(new_n781), .B2(G1966), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n749), .A2(G1961), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n782), .B(new_n783), .C1(new_n768), .C2(new_n767), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n761), .A2(new_n765), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n764), .A2(G2090), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n697), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n556), .B2(new_n697), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1341), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n715), .A2(G26), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT28), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n473), .A2(G140), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT95), .Z(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n795));
  INV_X1    g370(.A(G116), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(G2105), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G128), .B2(new_n487), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n792), .B1(new_n800), .B2(new_n736), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G2067), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT31), .B(G11), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT101), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(G28), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n736), .B1(new_n805), .B2(G28), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n804), .B1(new_n806), .B2(new_n807), .C1(new_n643), .C2(new_n715), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n801), .B2(G2067), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n781), .A2(G1966), .ZN(new_n810));
  NAND2_X1  g385(.A1(G160), .A2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT24), .B(G34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n715), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT98), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G2084), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n802), .A2(new_n809), .A3(new_n810), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT99), .Z(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n785), .A2(new_n786), .A3(new_n790), .A4(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n735), .B1(new_n824), .B2(new_n825), .ZN(G311));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  INV_X1    g402(.A(new_n735), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(G150));
  NOR2_X1   g404(.A1(new_n619), .A2(new_n626), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n521), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n524), .A2(new_n835), .B1(new_n526), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n552), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n838), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n839), .B1(new_n555), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n832), .B(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n838), .A2(new_n844), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  XOR2_X1   g424(.A(G162), .B(new_n643), .Z(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(G160), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n799), .B(G164), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n758), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n744), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n743), .B2(new_n853), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n722), .B(new_n634), .Z(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n487), .A2(G130), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT105), .ZN(new_n861));
  AOI211_X1 g436(.A(new_n859), .B(new_n861), .C1(G142), .C2(new_n473), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n856), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n855), .A2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n851), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(new_n851), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n869), .A3(new_n864), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g448(.A(new_n603), .B(new_n707), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n876));
  NAND2_X1  g451(.A1(G303), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(G166), .A2(KEYINPUT106), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(G290), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(G290), .B1(new_n877), .B2(new_n878), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n874), .A3(new_n879), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT108), .Z(new_n888));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT107), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n841), .B(new_n628), .Z(new_n894));
  OR2_X1    g469(.A1(new_n619), .A2(G299), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n619), .A2(G299), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n895), .A2(KEYINPUT41), .A3(new_n896), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n898), .B1(new_n901), .B2(new_n894), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n893), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G868), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n838), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n838), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n581), .A2(G171), .ZN(new_n908));
  NOR2_X1   g483(.A1(G168), .A2(G171), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n841), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G301), .B1(new_n575), .B2(new_n580), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n838), .B1(new_n553), .B2(new_n554), .ZN(new_n913));
  OAI22_X1  g488(.A1(new_n912), .A2(new_n909), .B1(new_n913), .B2(new_n839), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(KEYINPUT109), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n841), .A2(new_n908), .A3(new_n916), .A4(new_n910), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n901), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n897), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n919), .A3(new_n914), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n918), .A2(new_n891), .A3(new_n890), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n871), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n918), .A2(new_n920), .B1(new_n891), .B2(new_n890), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n907), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n911), .A2(new_n914), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n901), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT110), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n901), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n897), .B1(new_n915), .B2(new_n917), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n929), .B(new_n931), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n892), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n922), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n926), .B1(new_n938), .B2(new_n925), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n925), .A3(new_n937), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n922), .B2(new_n923), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT112), .B1(new_n942), .B2(new_n907), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n944), .B(KEYINPUT44), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n939), .B1(new_n943), .B2(new_n945), .ZN(G397));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n512), .A2(new_n514), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n487), .A2(G126), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n499), .A2(new_n501), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n508), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n947), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(G137), .A2(new_n473), .B1(new_n466), .B2(new_n469), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT70), .B1(new_n481), .B2(G2105), .ZN(new_n956));
  AOI211_X1 g531(.A(new_n483), .B(new_n467), .C1(new_n479), .C2(new_n480), .ZN(new_n957));
  OAI211_X1 g532(.A(G40), .B(new_n955), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n722), .B(new_n724), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT114), .ZN(new_n961));
  INV_X1    g536(.A(G2067), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n799), .B(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n757), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n959), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1986), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n968), .A3(new_n610), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n967), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n959), .A2(new_n964), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  INV_X1    g550(.A(new_n963), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n959), .B1(new_n976), .B2(new_n757), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  NAND2_X1  g554(.A1(new_n722), .A2(new_n724), .ZN(new_n980));
  OAI22_X1  g555(.A1(new_n966), .A2(new_n980), .B1(G2067), .B2(new_n799), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n973), .B(new_n979), .C1(new_n959), .C2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n958), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n515), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n954), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n515), .A2(new_n988), .A3(new_n947), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n983), .A3(new_n989), .ZN(new_n990));
  OAI22_X1  g565(.A1(new_n986), .A2(G1966), .B1(G2084), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G8), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(G168), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(KEYINPUT51), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n997));
  INV_X1    g572(.A(G168), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(G8), .C1(new_n991), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT125), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n991), .B2(new_n994), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n991), .A2(new_n1000), .A3(new_n994), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n996), .B(new_n999), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n707), .A2(G1976), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1005), .B(G8), .C1(new_n952), .C2(new_n958), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT116), .B(G1976), .Z(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(G288), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n1012));
  OAI21_X1  g587(.A(G1981), .B1(new_n597), .B2(new_n602), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n571), .A2(G86), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n589), .A2(G48), .ZN(new_n1015));
  INV_X1    g590(.A(G1981), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n601), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT117), .B(KEYINPUT49), .Z(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1012), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g596(.A(KEYINPUT118), .B(new_n1019), .C1(new_n1013), .C2(new_n1017), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1021), .A2(new_n1022), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1024));
  INV_X1    g599(.A(new_n952), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n983), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G8), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1010), .B(new_n1011), .C1(new_n1024), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n986), .A2(G1971), .B1(G2090), .B2(new_n990), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(G166), .B2(new_n993), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1030), .A2(new_n1035), .A3(G8), .A4(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n515), .A2(new_n988), .A3(new_n947), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n988), .B1(new_n515), .B2(new_n947), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n958), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1040), .A2(new_n1041), .B1(new_n985), .B2(new_n700), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1033), .B(new_n1031), .C1(new_n1042), .C2(new_n993), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1029), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n985), .B2(G2078), .ZN(new_n1047));
  INV_X1    g622(.A(G1961), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n990), .A2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1046), .A2(G2078), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n986), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(G301), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1004), .A2(new_n1045), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT127), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(G301), .A3(new_n1052), .ZN(new_n1058));
  AND4_X1   g633(.A1(G40), .A2(new_n955), .A3(new_n482), .A4(new_n1051), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n954), .A2(new_n1059), .A3(new_n984), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1047), .A2(new_n1049), .A3(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1061), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT126), .B1(new_n1061), .B2(G171), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT54), .B(new_n1058), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1061), .A2(G171), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1053), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1064), .A2(new_n1003), .A3(new_n1067), .A4(new_n1045), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n952), .A2(new_n958), .A3(G2067), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT60), .B(new_n1071), .C1(new_n1040), .C2(G1348), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n1075));
  AOI211_X1 g650(.A(new_n1075), .B(new_n1070), .C1(new_n990), .C2(new_n768), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n620), .B1(new_n1076), .B2(KEYINPUT123), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1072), .A2(new_n1073), .A3(new_n619), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1070), .B1(new_n990), .B2(new_n768), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(KEYINPUT60), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1069), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  INV_X1    g658(.A(G1956), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n990), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT56), .B(G2072), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n954), .A2(new_n983), .A3(new_n984), .A4(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1085), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1088), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1083), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1085), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(KEYINPUT61), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1099), .B(KEYINPUT122), .Z(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n952), .B2(new_n958), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT120), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n954), .A2(new_n964), .A3(new_n983), .A4(new_n984), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n1102), .C1(new_n952), .C2(new_n958), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n556), .ZN(new_n1109));
  NOR2_X1   g684(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1101), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1110), .B(new_n1100), .C1(new_n1108), .C2(new_n556), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1093), .B(new_n1098), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1076), .A2(KEYINPUT123), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT123), .B(new_n620), .C1(new_n1080), .C2(KEYINPUT60), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n619), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1081), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(KEYINPUT124), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1082), .A2(new_n1115), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1080), .A2(new_n619), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1097), .B1(new_n1123), .B2(new_n1092), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1068), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1037), .A2(new_n1028), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G288), .A2(G1976), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1017), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1027), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n991), .A2(G8), .A3(new_n581), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1134), .A2(new_n1044), .A3(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1132), .B(KEYINPUT119), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT63), .B1(new_n1137), .B2(new_n1045), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1131), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1057), .B1(new_n1125), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1131), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1135), .B1(new_n1134), .B2(new_n1044), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(new_n1045), .A3(KEYINPUT63), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1124), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1114), .B1(new_n1146), .B2(new_n1069), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1147), .B2(new_n1121), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT127), .B(new_n1144), .C1(new_n1148), .C2(new_n1068), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1056), .B1(new_n1140), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n959), .A2(G1986), .A3(G290), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n969), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT113), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n967), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n982), .B1(new_n1150), .B2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g730(.A1(G227), .A2(new_n461), .A3(G401), .A4(G229), .ZN(new_n1157));
  NAND3_X1  g731(.A1(new_n872), .A2(new_n1157), .A3(new_n942), .ZN(G225));
  INV_X1    g732(.A(G225), .ZN(G308));
endmodule


