//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n203), .A2(G50), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n209), .B1(new_n213), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G58), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n210), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  OAI22_X1  g0049(.A1(new_n249), .A2(new_n216), .B1(new_n211), .B2(G68), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G50), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n246), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT11), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n257), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n202), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT12), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n246), .B1(new_n260), .B2(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n257), .A2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G68), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n256), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  OAI211_X1 g0071(.A(G232), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT73), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n247), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT73), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(G232), .A4(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G97), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(G226), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n273), .A2(new_n279), .A3(new_n280), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G1), .A3(G13), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(new_n285), .A3(G274), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n285), .A2(G238), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT74), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT74), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n287), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT13), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n287), .A2(new_n301), .A3(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n269), .B1(new_n303), .B2(G200), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n287), .A2(new_n301), .A3(new_n298), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n287), .B2(new_n298), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT75), .B1(new_n307), .B2(G190), .ZN(new_n308));
  AND4_X1   g0108(.A1(KEYINPUT75), .A2(new_n300), .A3(G190), .A4(new_n302), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n304), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(KEYINPUT76), .B(new_n304), .C1(new_n308), .C2(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT14), .B1(new_n307), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n303), .A2(new_n317), .A3(G169), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n316), .B(new_n318), .C1(new_n319), .C2(new_n303), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n269), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(new_n322), .B(KEYINPUT77), .Z(new_n323));
  INV_X1    g0123(.A(G226), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G1698), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G223), .B2(G1698), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT78), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n247), .A2(KEYINPUT78), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT3), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(new_n275), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n286), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G232), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n285), .A2(new_n292), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n291), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(G169), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G223), .A2(G1698), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n324), .B2(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n247), .A2(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n327), .A2(G33), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n274), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n344), .B2(new_n271), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n285), .B1(new_n345), .B2(new_n332), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n346), .A2(G179), .A3(new_n337), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT80), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n334), .A2(new_n319), .A3(new_n338), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n315), .B1(new_n346), .B2(new_n337), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT80), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT8), .B(G58), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n257), .B2(G20), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n263), .A2(new_n354), .B1(new_n355), .B2(new_n266), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n201), .A2(new_n202), .ZN(new_n357));
  NOR2_X1   g0157(.A1(G58), .A2(G68), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n251), .A2(G159), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT78), .B(G33), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n211), .B(new_n275), .C1(new_n363), .C2(new_n274), .ZN(new_n364));
  OAI21_X1  g0164(.A(G68), .B1(new_n364), .B2(KEYINPUT7), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n342), .A2(new_n343), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n271), .B1(new_n367), .B2(KEYINPUT3), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n366), .B1(new_n368), .B2(new_n211), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT16), .B(new_n362), .C1(new_n365), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n246), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n363), .B2(new_n274), .ZN(new_n373));
  AOI21_X1  g0173(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n275), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(G68), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n361), .B1(new_n376), .B2(KEYINPUT79), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT79), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(G68), .C1(new_n373), .C2(new_n375), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT16), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n356), .B1(new_n371), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n353), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT18), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT18), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n353), .A2(new_n384), .A3(new_n381), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n334), .A2(new_n386), .A3(new_n338), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n346), .B2(new_n337), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n356), .B(new_n390), .C1(new_n371), .C2(new_n380), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n371), .A2(new_n380), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n394), .A2(KEYINPUT17), .A3(new_n356), .A4(new_n390), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n383), .A2(new_n385), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n277), .A2(G223), .A3(G1698), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n277), .A2(new_n281), .ZN(new_n399));
  INV_X1    g0199(.A(G222), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n398), .B1(new_n216), .B2(new_n277), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n286), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n291), .C1(new_n324), .C2(new_n336), .ZN(new_n403));
  INV_X1    g0203(.A(new_n246), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT67), .ZN(new_n406));
  INV_X1    g0206(.A(new_n354), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n248), .B1(G150), .B2(new_n251), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n266), .A2(G50), .A3(new_n267), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G50), .B2(new_n262), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n403), .A2(G200), .B1(new_n412), .B2(KEYINPUT9), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n412), .A2(KEYINPUT9), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(new_n386), .C2(new_n403), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT10), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n412), .B1(new_n403), .B2(new_n315), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G179), .B2(new_n403), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n277), .A2(G238), .A3(G1698), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n422), .B1(new_n218), .B2(new_n277), .C1(new_n399), .C2(new_n335), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n285), .B1(new_n423), .B2(KEYINPUT69), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(KEYINPUT69), .B2(new_n423), .ZN(new_n425));
  INV_X1    g0225(.A(new_n291), .ZN(new_n426));
  INV_X1    g0226(.A(new_n336), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(G244), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G200), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n407), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT70), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT15), .B(G87), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n249), .ZN(new_n434));
  INV_X1    g0234(.A(new_n433), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(KEYINPUT70), .A3(new_n248), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n431), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n246), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT71), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n216), .B1(new_n257), .B2(G20), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n263), .A2(new_n216), .B1(new_n266), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n430), .A2(KEYINPUT72), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT72), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(new_n441), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n388), .B1(new_n425), .B2(new_n428), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n442), .B(new_n446), .C1(new_n386), .C2(new_n429), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n429), .A2(new_n315), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n425), .A2(new_n319), .A3(new_n428), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n397), .A2(new_n421), .A3(new_n447), .A4(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n323), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n257), .A2(G33), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n262), .A2(new_n404), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n266), .A2(KEYINPUT83), .A3(new_n453), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(G107), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n260), .A2(new_n218), .A3(new_n261), .ZN(new_n459));
  XOR2_X1   g0259(.A(new_n459), .B(KEYINPUT25), .Z(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT93), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT93), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n211), .A2(G107), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT92), .A2(KEYINPUT23), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT92), .A2(KEYINPUT23), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n367), .A2(G116), .ZN(new_n470));
  OAI221_X1 g0270(.A(new_n469), .B1(new_n468), .B2(new_n466), .C1(new_n470), .C2(G20), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n211), .B(G87), .C1(new_n344), .C2(new_n271), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT91), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n275), .B1(new_n363), .B2(new_n274), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(KEYINPUT91), .A3(new_n211), .A4(G87), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(KEYINPUT22), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n270), .A2(new_n271), .ZN(new_n478));
  INV_X1    g0278(.A(G87), .ZN(new_n479));
  OR4_X1    g0279(.A1(KEYINPUT22), .A2(new_n478), .A3(G20), .A4(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n471), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n246), .B1(new_n481), .B2(KEYINPUT24), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  AOI211_X1 g0283(.A(new_n483), .B(new_n471), .C1(new_n477), .C2(new_n480), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n465), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT94), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G250), .A2(G1698), .ZN(new_n487));
  INV_X1    g0287(.A(G257), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(G1698), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n344), .B2(new_n271), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n367), .A2(G294), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n285), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n288), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n289), .A2(G1), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G264), .A3(new_n285), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n486), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G274), .ZN(new_n502));
  INV_X1    g0302(.A(new_n210), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n284), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(new_n496), .A3(new_n495), .A4(new_n497), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n475), .A2(new_n489), .B1(G294), .B2(new_n367), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT94), .B(new_n499), .C1(new_n506), .C2(new_n285), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n501), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n505), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n492), .A2(new_n500), .A3(new_n509), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n508), .A2(new_n319), .B1(new_n510), .B2(new_n315), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n485), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n388), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n386), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n515), .B(new_n465), .C1(new_n484), .C2(new_n482), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n262), .A2(G97), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n456), .A2(new_n457), .ZN(new_n520));
  INV_X1    g0320(.A(G97), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT82), .ZN(new_n523));
  OAI211_X1 g0323(.A(KEYINPUT7), .B(new_n374), .C1(new_n367), .C2(KEYINPUT3), .ZN(new_n524));
  INV_X1    g0324(.A(new_n375), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n218), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n527), .A2(KEYINPUT81), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(KEYINPUT81), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n521), .A2(new_n218), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(G97), .A3(new_n218), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n211), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n252), .A2(new_n216), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n526), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n523), .B1(new_n537), .B2(new_n404), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n535), .A2(new_n536), .ZN(new_n539));
  OAI211_X1 g0339(.A(KEYINPUT82), .B(new_n246), .C1(new_n539), .C2(new_n526), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n522), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n217), .A2(G1698), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT4), .B1(new_n475), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(KEYINPUT4), .A2(G244), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n281), .B(new_n544), .C1(new_n270), .C2(new_n271), .ZN(new_n545));
  OAI211_X1 g0345(.A(G250), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT84), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT84), .ZN(new_n551));
  INV_X1    g0351(.A(new_n542), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n330), .B2(new_n275), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n550), .B(new_n551), .C1(new_n553), .C2(KEYINPUT4), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n286), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n498), .A2(new_n285), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n505), .B1(new_n556), .B2(new_n488), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(G179), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n541), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n315), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n555), .A2(new_n386), .A3(new_n558), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n550), .B1(new_n553), .B2(KEYINPUT4), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n285), .B1(new_n564), .B2(KEYINPUT84), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n557), .B1(new_n565), .B2(new_n554), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n563), .B1(new_n566), .B2(G200), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n561), .A2(new_n562), .B1(new_n541), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT88), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n504), .A2(new_n497), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n285), .B(G250), .C1(G1), .C2(new_n289), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G238), .A2(G1698), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n217), .B2(G1698), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n344), .B2(new_n271), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n470), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n577), .B2(new_n286), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n570), .B1(new_n578), .B2(G190), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n285), .B1(new_n576), .B2(new_n470), .ZN(new_n580));
  NOR4_X1   g0380(.A1(new_n580), .A2(KEYINPUT87), .A3(new_n386), .A4(new_n573), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n569), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n262), .A2(new_n435), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n211), .B(G68), .C1(new_n344), .C2(new_n271), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n248), .A2(new_n586), .A3(G97), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n531), .A2(new_n479), .B1(new_n280), .B2(new_n211), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n586), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(KEYINPUT86), .B(new_n584), .C1(new_n590), .C2(new_n404), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT86), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n404), .B1(new_n585), .B2(new_n589), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n583), .ZN(new_n594));
  INV_X1    g0394(.A(new_n520), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n591), .A2(new_n594), .B1(new_n595), .B2(G87), .ZN(new_n596));
  INV_X1    g0396(.A(new_n573), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n475), .A2(new_n575), .B1(G116), .B2(new_n367), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(G190), .C1(new_n598), .C2(new_n285), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT87), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n578), .A2(new_n570), .A3(G190), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT88), .ZN(new_n602));
  INV_X1    g0402(.A(new_n578), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n582), .A2(new_n596), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n591), .A2(new_n594), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n595), .A2(new_n435), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n603), .A2(new_n315), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n578), .A2(new_n319), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(G257), .A2(G1698), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n219), .B2(G1698), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n344), .B2(new_n271), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n478), .A2(G303), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n286), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n498), .A2(G270), .A3(new_n285), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n505), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT89), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n285), .B1(new_n615), .B2(new_n616), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT89), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(G190), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(G20), .B1(G33), .B2(G283), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n247), .A2(G97), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G116), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n245), .A2(new_n210), .B1(G20), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT20), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n629), .A2(new_n630), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT90), .B1(new_n627), .B2(new_n628), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n633), .B(KEYINPUT20), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n632), .B1(new_n266), .B2(new_n453), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n263), .A2(G116), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n634), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n618), .A2(KEYINPUT89), .A3(new_n621), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n624), .B1(new_n623), .B2(new_n620), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(G200), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n626), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n641), .A2(G169), .A3(new_n644), .A4(new_n643), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n640), .A2(new_n639), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT20), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n637), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n315), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n655), .A2(KEYINPUT21), .A3(new_n644), .A4(new_n643), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n623), .A2(new_n620), .A3(new_n319), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n641), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n646), .A2(new_n649), .A3(new_n656), .A4(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n612), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n452), .A2(new_n517), .A3(new_n568), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT95), .ZN(G372));
  INV_X1    g0462(.A(new_n541), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n566), .A2(new_n319), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n562), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n665), .A2(new_n612), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n665), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT96), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n580), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n598), .A2(KEYINPUT96), .A3(new_n285), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n597), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n315), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n608), .A2(new_n673), .A3(new_n610), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(G200), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n600), .A2(new_n601), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n596), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT97), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n674), .B2(new_n677), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n668), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n667), .B1(new_n681), .B2(new_n666), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n674), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n649), .A2(new_n656), .A3(new_n658), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n512), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n686), .A2(new_n568), .A3(new_n516), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n679), .A2(new_n680), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n684), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n452), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n310), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n321), .B1(new_n693), .B2(new_n450), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n391), .B(KEYINPUT17), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n353), .A2(new_n384), .A3(new_n381), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n384), .B1(new_n353), .B2(new_n381), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT98), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n417), .B1(new_n700), .B2(KEYINPUT98), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n420), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n692), .A2(new_n703), .ZN(G369));
  NAND3_X1  g0504(.A1(new_n257), .A2(new_n211), .A3(G13), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n642), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n685), .A2(new_n646), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n685), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n485), .A2(new_n710), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n517), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n512), .B2(new_n711), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n485), .A2(new_n511), .A3(new_n711), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n685), .A2(new_n710), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n517), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n207), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G1), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n531), .A2(new_n479), .A3(new_n632), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n729), .A2(new_n730), .B1(new_n214), .B2(new_n728), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n691), .A2(new_n733), .A3(new_n711), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n665), .A2(new_n612), .A3(KEYINPUT26), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n681), .B2(KEYINPUT26), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n710), .B1(new_n690), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n734), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G330), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n517), .A2(new_n568), .A3(new_n660), .A4(new_n711), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n643), .A2(new_n644), .A3(new_n319), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n559), .A3(new_n508), .A4(new_n672), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n657), .A2(new_n501), .A3(new_n507), .A4(new_n578), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(new_n559), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n501), .A2(new_n507), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n623), .A2(new_n620), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n748), .A2(G179), .A3(new_n578), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n566), .A2(new_n747), .A3(new_n749), .A4(KEYINPUT30), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n743), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n752));
  AOI21_X1  g0552(.A(KEYINPUT31), .B1(new_n751), .B2(new_n710), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n740), .B1(new_n741), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n739), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n732), .B1(new_n758), .B2(G1), .ZN(G364));
  AND2_X1   g0559(.A1(new_n211), .A2(G13), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n257), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n727), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n717), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G330), .B2(new_n715), .ZN(new_n765));
  INV_X1    g0565(.A(new_n763), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n726), .A2(new_n478), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G355), .B1(new_n632), .B2(new_n726), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n243), .A2(new_n289), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n475), .A2(new_n726), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G45), .B2(new_n214), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n210), .B1(G20), .B2(new_n315), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT99), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n766), .B1(new_n772), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(KEYINPUT100), .ZN(new_n781));
  INV_X1    g0581(.A(new_n776), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n211), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n386), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n218), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n211), .A2(new_n319), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n386), .A2(G179), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n211), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n789), .A2(new_n201), .B1(new_n521), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n787), .A2(new_n388), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n785), .B(new_n792), .C1(G50), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G190), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n783), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT101), .B(KEYINPUT32), .Z(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(G159), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n797), .B2(G159), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(G87), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n786), .A2(new_n386), .A3(G200), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n277), .B1(new_n804), .B2(new_n202), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n786), .A2(new_n795), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(G77), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n794), .A2(new_n799), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G322), .ZN(new_n810));
  INV_X1    g0610(.A(new_n793), .ZN(new_n811));
  INV_X1    g0611(.A(G326), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n789), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n784), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G283), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n804), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n277), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G311), .A2(new_n807), .B1(new_n797), .B2(G329), .ZN(new_n819));
  INV_X1    g0619(.A(new_n791), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(G294), .B1(new_n802), .B2(G303), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n815), .A2(new_n818), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n782), .B1(new_n809), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n780), .A2(KEYINPUT100), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n775), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n781), .B(new_n825), .C1(new_n715), .C2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n765), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n691), .A2(new_n711), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n450), .A2(new_n710), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n444), .A2(new_n710), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n447), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(new_n450), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n830), .B(new_n834), .Z(new_n835));
  AOI21_X1  g0635(.A(new_n763), .B1(new_n835), .B2(new_n756), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n756), .B2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(G303), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n811), .A2(new_n838), .B1(new_n784), .B2(new_n479), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G294), .B2(new_n788), .ZN(new_n840));
  INV_X1    g0640(.A(G311), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n806), .A2(new_n632), .B1(new_n796), .B2(new_n841), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n277), .B(new_n842), .C1(G283), .C2(new_n816), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n820), .A2(G97), .B1(new_n802), .B2(G107), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n840), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n816), .A2(G150), .B1(new_n807), .B2(G159), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n788), .A2(G143), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n811), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n368), .B1(G132), .B2(new_n797), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n791), .A2(new_n201), .B1(new_n801), .B2(new_n253), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n784), .A2(new_n202), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n849), .A2(new_n850), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n782), .B1(new_n858), .B2(KEYINPUT102), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(KEYINPUT102), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n776), .A2(new_n773), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n766), .B1(new_n216), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(new_n834), .C2(new_n774), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n837), .A2(new_n863), .ZN(G384));
  NAND2_X1  g0664(.A1(new_n532), .A2(new_n534), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n632), .B(new_n213), .C1(new_n865), .C2(KEYINPUT35), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(KEYINPUT35), .B2(new_n865), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT36), .Z(new_n868));
  NOR3_X1   g0668(.A1(new_n214), .A2(new_n216), .A3(new_n357), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT103), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n869), .A2(KEYINPUT103), .B1(new_n253), .B2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n257), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n708), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n699), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n368), .A2(new_n366), .A3(new_n211), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n364), .A2(KEYINPUT7), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(G68), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n879), .B2(new_n362), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n356), .B1(new_n371), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n874), .ZN(new_n882));
  INV_X1    g0682(.A(new_n352), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n351), .B1(new_n349), .B2(new_n350), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n356), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n370), .A2(new_n246), .ZN(new_n887));
  INV_X1    g0687(.A(new_n880), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n882), .B(new_n391), .C1(new_n885), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n381), .A2(new_n874), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n382), .A2(new_n892), .A3(new_n893), .A4(new_n391), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n882), .B1(new_n699), .B2(new_n695), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n876), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n882), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n396), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n891), .A2(new_n894), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n893), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n396), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n382), .A2(new_n391), .A3(new_n893), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n894), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT106), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n897), .B(new_n901), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT39), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n907), .ZN(new_n912));
  NOR2_X1   g0712(.A1(KEYINPUT106), .A2(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n320), .A2(new_n269), .A3(new_n711), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n875), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n269), .A2(new_n710), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n321), .A2(new_n310), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n320), .B1(new_n312), .B2(new_n313), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n686), .A2(new_n568), .A3(new_n516), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n674), .B1(new_n924), .B2(new_n688), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n711), .B(new_n834), .C1(new_n925), .C2(new_n682), .ZN(new_n926));
  INV_X1    g0726(.A(new_n831), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT104), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n897), .B2(new_n901), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n899), .B2(new_n900), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n911), .A2(new_n933), .A3(KEYINPUT105), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n928), .A2(KEYINPUT104), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n918), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n738), .A2(new_n452), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(new_n703), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n741), .A2(new_n754), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n922), .A2(new_n941), .A3(new_n834), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n934), .B2(new_n932), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n903), .A2(new_n906), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n876), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n940), .B1(new_n945), .B2(new_n901), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n946), .A3(KEYINPUT107), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT107), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT40), .B1(new_n911), .B2(new_n907), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n922), .A2(new_n941), .A3(new_n834), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n940), .A2(new_n943), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n452), .A2(new_n941), .ZN(new_n954));
  OAI21_X1  g0754(.A(G330), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n953), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n939), .A2(new_n956), .B1(new_n257), .B2(new_n760), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n939), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n873), .B1(new_n957), .B2(new_n958), .ZN(G367));
  OAI21_X1  g0759(.A(new_n568), .B1(new_n541), .B2(new_n711), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n668), .A2(new_n710), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(new_n724), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n665), .B1(new_n960), .B2(new_n512), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n963), .A2(KEYINPUT42), .B1(new_n711), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(KEYINPUT42), .B2(new_n963), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n596), .A2(new_n711), .ZN(new_n968));
  MUX2_X1   g0768(.A(new_n688), .B(new_n674), .S(new_n968), .Z(new_n969));
  OAI21_X1  g0769(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n967), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n721), .A2(new_n962), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n972), .B(new_n973), .Z(new_n974));
  INV_X1    g0774(.A(KEYINPUT109), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n724), .A2(new_n722), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n962), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT44), .Z(new_n978));
  NOR2_X1   g0778(.A1(new_n962), .A2(new_n976), .ZN(new_n979));
  XNOR2_X1  g0779(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n721), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n978), .A2(new_n721), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n724), .B1(new_n720), .B2(new_n723), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(new_n716), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n739), .A2(new_n989), .A3(new_n756), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n975), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n990), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n992), .A2(KEYINPUT109), .A3(new_n985), .A4(new_n984), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n757), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n727), .B(KEYINPUT41), .Z(new_n995));
  OAI21_X1  g0795(.A(new_n761), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n974), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n770), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n235), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n777), .B1(new_n207), .B2(new_n433), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n763), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(G159), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n804), .A2(new_n1002), .B1(new_n806), .B2(new_n253), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n478), .B(new_n1003), .C1(G137), .C2(new_n797), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n788), .A2(G150), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n791), .A2(new_n202), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G77), .B2(new_n814), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n793), .A2(G143), .B1(new_n802), .B2(G58), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n788), .A2(G303), .B1(new_n814), .B2(G97), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n841), .B2(new_n811), .ZN(new_n1011));
  INV_X1    g0811(.A(G283), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n791), .A2(new_n218), .B1(new_n806), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1011), .B1(KEYINPUT110), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(KEYINPUT110), .B2(new_n1013), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n816), .A2(G294), .B1(new_n797), .B2(G317), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT46), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n801), .B2(new_n632), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n802), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n368), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1009), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT47), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1001), .B1(new_n1022), .B2(new_n776), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT111), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n969), .A2(new_n775), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n997), .A2(new_n1027), .ZN(G387));
  NAND2_X1  g0828(.A1(new_n757), .A2(new_n988), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n727), .A3(new_n990), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n720), .A2(new_n826), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n767), .A2(new_n730), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(G107), .B2(new_n207), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n231), .A2(new_n289), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n354), .A2(G50), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT50), .ZN(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n730), .C1(G68), .C2(G77), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n998), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1033), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n763), .B1(new_n1039), .B2(new_n778), .ZN(new_n1040));
  XOR2_X1   g0840(.A(KEYINPUT112), .B(G150), .Z(new_n1041));
  OAI22_X1  g0841(.A1(new_n1041), .A2(new_n796), .B1(new_n806), .B2(new_n202), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n407), .B2(new_n816), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n793), .A2(G159), .B1(new_n802), .B2(G77), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n435), .A2(new_n820), .B1(new_n788), .B2(G50), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n368), .B1(G97), .B2(new_n814), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(G294), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n791), .A2(new_n1012), .B1(new_n801), .B2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n816), .A2(G311), .B1(new_n807), .B2(G303), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n788), .A2(G317), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n810), .C2(new_n811), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n1053), .B2(new_n1052), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT49), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n368), .B1(new_n812), .B2(new_n796), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G116), .B2(new_n814), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1047), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1040), .B1(new_n1061), .B2(new_n776), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n989), .A2(new_n762), .B1(new_n1031), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1030), .A2(new_n1063), .ZN(G393));
  NAND2_X1  g0864(.A1(new_n991), .A2(new_n993), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n728), .B1(new_n986), .B2(new_n990), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n986), .A2(new_n761), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n962), .A2(new_n775), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n202), .A2(new_n801), .B1(new_n784), .B2(new_n479), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n368), .B(new_n1070), .C1(G143), .C2(new_n797), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT113), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G150), .A2(new_n793), .B1(new_n788), .B2(G159), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n791), .A2(new_n216), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n804), .A2(new_n253), .B1(new_n806), .B2(new_n354), .ZN(new_n1076));
  OR4_X1    g0876(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G311), .A2(new_n788), .B1(new_n793), .B2(G317), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT52), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n806), .A2(new_n1048), .B1(new_n796), .B2(new_n810), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n277), .B(new_n1080), .C1(G303), .C2(new_n816), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n801), .A2(new_n1012), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n785), .B(new_n1082), .C1(G116), .C2(new_n820), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n782), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n240), .A2(new_n770), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n776), .B(new_n775), .C1(G97), .C2(new_n726), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n766), .B(new_n1085), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1068), .B1(new_n1069), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1067), .A2(new_n1089), .ZN(G390));
  XNOR2_X1  g0890(.A(new_n916), .B(KEYINPUT114), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n912), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n833), .A2(new_n450), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n831), .B1(new_n737), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1094), .B2(new_n923), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n909), .A2(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n928), .B2(new_n917), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n755), .A2(new_n834), .A3(new_n922), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n755), .A2(new_n834), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n923), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1094), .A2(new_n1103), .A3(new_n1098), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1098), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n926), .A2(new_n927), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n452), .A2(new_n755), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n937), .A2(new_n1110), .A3(new_n703), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n727), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1096), .A2(new_n773), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n806), .A2(new_n521), .B1(new_n796), .B2(new_n1048), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n277), .B(new_n1117), .C1(G107), .C2(new_n816), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n793), .A2(G283), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1075), .B1(G116), .B2(new_n788), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n854), .B1(G87), .B2(new_n802), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(G128), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n811), .A2(new_n1123), .B1(new_n1002), .B2(new_n791), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G132), .B2(new_n788), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1041), .A2(new_n801), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n797), .A2(G125), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n816), .A2(G137), .B1(new_n807), .B2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n277), .B1(new_n784), .B2(new_n253), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT116), .Z(new_n1134));
  OAI21_X1  g0934(.A(new_n1122), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n776), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n861), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n763), .B1(new_n407), .B2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT115), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT117), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1101), .A2(new_n762), .B1(new_n1116), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1115), .A2(new_n1142), .ZN(G378));
  INV_X1    g0943(.A(KEYINPUT119), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1096), .A2(new_n916), .B1(new_n699), .B2(new_n874), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n934), .A2(new_n932), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1106), .A2(new_n922), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT104), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1145), .B1(new_n1149), .B2(new_n929), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n943), .A2(new_n940), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n947), .A2(new_n951), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(G330), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n416), .A2(new_n419), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n874), .B1(new_n409), .B2(new_n411), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT55), .Z(new_n1156));
  XOR2_X1   g0956(.A(new_n1154), .B(new_n1156), .Z(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1154), .B(new_n1156), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1158), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1153), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n952), .A2(G330), .A3(new_n1163), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1150), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1149), .A2(new_n929), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1165), .A2(new_n1166), .B1(new_n1168), .B2(new_n918), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1144), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1163), .B1(new_n952), .B2(G330), .ZN(new_n1171));
  AND4_X1   g0971(.A1(G330), .A2(new_n1151), .A3(new_n1152), .A4(new_n1163), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n936), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1150), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(KEYINPUT119), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1111), .B1(new_n1101), .B2(new_n1112), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1173), .A2(KEYINPUT57), .A3(new_n1174), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n727), .B1(new_n1180), .B2(new_n1177), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G132), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n804), .A2(new_n1183), .B1(new_n806), .B2(new_n848), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G150), .A2(new_n820), .B1(new_n793), .B2(G125), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n1123), .B2(new_n789), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(new_n802), .C2(new_n1130), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT59), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n814), .A2(G159), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n816), .A2(G97), .B1(new_n797), .B2(G283), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n433), .B2(new_n806), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1006), .B(new_n1195), .C1(G77), .C2(new_n802), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n789), .A2(new_n218), .B1(new_n784), .B2(new_n201), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G116), .B2(new_n793), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1196), .A2(new_n288), .A3(new_n368), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G50), .B1(new_n247), .B2(new_n288), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n475), .B2(G41), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1193), .A2(new_n1201), .A3(new_n1202), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n776), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n766), .B1(new_n253), .B2(new_n861), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n1164), .C2(new_n774), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1176), .B2(new_n762), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1182), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(G375));
  NOR2_X1   g1013(.A1(new_n922), .A2(new_n774), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT120), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n763), .B1(G68), .B2(new_n1137), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n816), .A2(G116), .B1(new_n807), .B2(G107), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1048), .B2(new_n811), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT121), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n478), .B1(new_n796), .B2(new_n838), .C1(new_n216), .C2(new_n784), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n820), .A2(new_n435), .B1(new_n802), .B2(G97), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1012), .B2(new_n789), .ZN(new_n1222));
  OR3_X1    g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT122), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n801), .A2(new_n1002), .B1(new_n796), .B2(new_n1123), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT123), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G50), .A2(new_n820), .B1(new_n788), .B2(G137), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n816), .A2(new_n1130), .B1(new_n807), .B2(G150), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n793), .A2(G132), .B1(new_n814), .B2(G58), .ZN(new_n1229));
  AND4_X1   g1029(.A1(new_n475), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1223), .A2(new_n1224), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1224), .B2(new_n1223), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1216), .B1(new_n1232), .B2(new_n776), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1108), .A2(new_n762), .B1(new_n1215), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n995), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1111), .B2(new_n1109), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(G381));
  AOI21_X1  g1038(.A(new_n1026), .B1(new_n974), .B2(new_n996), .ZN(new_n1239));
  INV_X1    g1039(.A(G378), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1030), .A2(new_n828), .A3(new_n1063), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1212), .A2(new_n1239), .A3(new_n1240), .A4(new_n1242), .ZN(G407));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G343), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1212), .A2(new_n1240), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(G407), .A2(G213), .A3(new_n1246), .ZN(G409));
  AND3_X1   g1047(.A1(new_n1030), .A2(new_n828), .A3(new_n1063), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n828), .B1(new_n1030), .B2(new_n1063), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT125), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT125), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1241), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(G390), .A2(new_n1250), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G390), .B1(new_n1253), .B2(new_n1250), .ZN(new_n1256));
  OAI21_X1  g1056(.A(G387), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n1067), .A3(new_n1089), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n1239), .A3(new_n1254), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1210), .C1(new_n1179), .C2(new_n1181), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1173), .A2(KEYINPUT119), .A3(new_n1174), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT119), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1235), .B(new_n1178), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1173), .A2(new_n762), .A3(new_n1174), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1208), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(KEYINPUT124), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT124), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1269), .A3(new_n1208), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1265), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1240), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1245), .B1(new_n1262), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1112), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1237), .B1(new_n1274), .B2(KEYINPUT60), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1109), .A2(new_n1111), .A3(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n727), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1234), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(G384), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G384), .B(new_n1234), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT62), .B1(new_n1273), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1262), .A2(new_n1272), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1245), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT126), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1288), .B(new_n1245), .C1(new_n1262), .C2(new_n1272), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1283), .A2(KEYINPUT62), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1284), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1245), .A2(G2897), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1280), .A2(new_n1281), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1293), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1261), .B1(new_n1292), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1288), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1273), .A2(KEYINPUT126), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1283), .A2(KEYINPUT63), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT127), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1261), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1299), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1273), .B2(new_n1283), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1273), .A2(new_n1296), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT127), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1290), .A2(new_n1313), .A3(new_n1305), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1307), .A2(new_n1312), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1301), .A2(new_n1315), .ZN(G405));
  NAND2_X1  g1116(.A1(G375), .A2(new_n1240), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1262), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1283), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1317), .A2(new_n1262), .A3(new_n1282), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1261), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1319), .A2(new_n1308), .A3(new_n1320), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(G402));
endmodule


