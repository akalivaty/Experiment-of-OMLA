

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743;

  NOR2_X1 U360 ( .A1(G237), .A2(G953), .ZN(n488) );
  XNOR2_X1 U361 ( .A(n375), .B(KEYINPUT69), .ZN(n495) );
  INV_X1 U362 ( .A(G953), .ZN(n732) );
  AND2_X2 U363 ( .A1(n401), .A2(n403), .ZN(n408) );
  NOR2_X2 U364 ( .A1(n681), .A2(n682), .ZN(n545) );
  NOR2_X2 U365 ( .A1(n739), .A2(n742), .ZN(n547) );
  NOR2_X2 U366 ( .A1(n372), .A2(n609), .ZN(n578) );
  NOR2_X1 U367 ( .A1(n352), .A2(n359), .ZN(n584) );
  INV_X1 U368 ( .A(G143), .ZN(n373) );
  INV_X1 U369 ( .A(G134), .ZN(n390) );
  NOR2_X2 U370 ( .A1(n645), .A2(n743), .ZN(n618) );
  XNOR2_X1 U371 ( .A(KEYINPUT0), .B(n584), .ZN(n599) );
  AND2_X1 U372 ( .A1(n400), .A2(n399), .ZN(n398) );
  NAND2_X1 U373 ( .A1(n427), .A2(n426), .ZN(n405) );
  NAND2_X1 U374 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U375 ( .A(n495), .B(n390), .ZN(n374) );
  XNOR2_X1 U376 ( .A(n368), .B(n462), .ZN(n729) );
  XNOR2_X1 U377 ( .A(n379), .B(n378), .ZN(n348) );
  XNOR2_X1 U378 ( .A(n381), .B(G107), .ZN(n474) );
  XNOR2_X1 U379 ( .A(n465), .B(G146), .ZN(n368) );
  XNOR2_X1 U380 ( .A(n382), .B(G122), .ZN(n494) );
  INV_X1 U381 ( .A(G125), .ZN(n465) );
  NAND2_X1 U382 ( .A1(n425), .A2(n424), .ZN(n423) );
  INV_X1 U383 ( .A(G902), .ZN(n424) );
  INV_X1 U384 ( .A(n471), .ZN(n425) );
  NAND2_X1 U385 ( .A1(n466), .A2(n622), .ZN(n384) );
  INV_X1 U386 ( .A(G104), .ZN(n382) );
  XNOR2_X1 U387 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n462) );
  NAND2_X1 U388 ( .A1(n663), .A2(n664), .ZN(n372) );
  INV_X1 U389 ( .A(n383), .ZN(n357) );
  NAND2_X1 U390 ( .A1(n388), .A2(n500), .ZN(n386) );
  NOR2_X2 U391 ( .A1(n668), .A2(n592), .ZN(n664) );
  AND2_X1 U392 ( .A1(n542), .A2(n418), .ZN(n683) );
  INV_X1 U393 ( .A(n654), .ZN(n418) );
  XNOR2_X1 U394 ( .A(n536), .B(KEYINPUT110), .ZN(n537) );
  AND2_X1 U395 ( .A1(n607), .A2(n679), .ZN(n538) );
  XOR2_X1 U396 ( .A(G902), .B(KEYINPUT15), .Z(n500) );
  NOR2_X1 U397 ( .A1(n581), .A2(n522), .ZN(n539) );
  NAND2_X1 U398 ( .A1(n701), .A2(n471), .ZN(n427) );
  NAND2_X1 U399 ( .A1(n442), .A2(n448), .ZN(n420) );
  XNOR2_X1 U400 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n478) );
  INV_X1 U401 ( .A(G131), .ZN(n375) );
  XNOR2_X1 U402 ( .A(KEYINPUT11), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U403 ( .A(G143), .B(G113), .ZN(n486) );
  XOR2_X1 U404 ( .A(KEYINPUT100), .B(G140), .Z(n487) );
  XNOR2_X1 U405 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n455) );
  OR2_X1 U406 ( .A1(n423), .A2(n409), .ZN(n404) );
  INV_X1 U407 ( .A(n539), .ZN(n400) );
  AND2_X1 U408 ( .A1(n679), .A2(KEYINPUT19), .ZN(n362) );
  AND2_X1 U409 ( .A1(n383), .A2(n362), .ZN(n358) );
  NAND2_X1 U410 ( .A1(n357), .A2(n356), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n529), .B(n366), .ZN(n365) );
  XNOR2_X1 U412 ( .A(n531), .B(n528), .ZN(n366) );
  XNOR2_X1 U413 ( .A(n441), .B(n339), .ZN(n716) );
  XNOR2_X1 U414 ( .A(n380), .B(n348), .ZN(n441) );
  XNOR2_X1 U415 ( .A(n494), .B(n474), .ZN(n380) );
  XNOR2_X1 U416 ( .A(G128), .B(G119), .ZN(n510) );
  XOR2_X1 U417 ( .A(KEYINPUT23), .B(G110), .Z(n511) );
  XNOR2_X1 U418 ( .A(n509), .B(n729), .ZN(n461) );
  XNOR2_X1 U419 ( .A(KEYINPUT93), .B(KEYINPUT75), .ZN(n505) );
  XOR2_X1 U420 ( .A(KEYINPUT82), .B(KEYINPUT24), .Z(n506) );
  XNOR2_X1 U421 ( .A(n452), .B(n451), .ZN(n450) );
  XNOR2_X1 U422 ( .A(G104), .B(G107), .ZN(n452) );
  XNOR2_X1 U423 ( .A(G146), .B(G101), .ZN(n451) );
  XOR2_X1 U424 ( .A(KEYINPUT89), .B(G110), .Z(n467) );
  XNOR2_X1 U425 ( .A(n541), .B(KEYINPUT39), .ZN(n573) );
  INV_X1 U426 ( .A(n679), .ZN(n445) );
  XNOR2_X1 U427 ( .A(n594), .B(n453), .ZN(n363) );
  INV_X1 U428 ( .A(KEYINPUT22), .ZN(n453) );
  NAND2_X1 U429 ( .A1(n357), .A2(n354), .ZN(n566) );
  NAND2_X1 U430 ( .A1(n361), .A2(n360), .ZN(n359) );
  OR2_X1 U431 ( .A1(n679), .A2(KEYINPUT19), .ZN(n360) );
  NAND2_X1 U432 ( .A1(n385), .A2(n362), .ZN(n361) );
  XNOR2_X1 U433 ( .A(n371), .B(n369), .ZN(n549) );
  XNOR2_X1 U434 ( .A(n370), .B(KEYINPUT111), .ZN(n369) );
  NOR2_X1 U435 ( .A1(n546), .A2(n666), .ZN(n371) );
  INV_X1 U436 ( .A(KEYINPUT28), .ZN(n370) );
  AND2_X1 U437 ( .A1(n351), .A2(n355), .ZN(n350) );
  INV_X1 U438 ( .A(n358), .ZN(n351) );
  NOR2_X1 U439 ( .A1(n631), .A2(G902), .ZN(n498) );
  XNOR2_X1 U440 ( .A(n503), .B(n434), .ZN(n456) );
  XNOR2_X1 U441 ( .A(n504), .B(KEYINPUT94), .ZN(n434) );
  XNOR2_X1 U442 ( .A(n545), .B(n437), .ZN(n678) );
  INV_X1 U443 ( .A(KEYINPUT41), .ZN(n437) );
  NAND2_X1 U444 ( .A1(n683), .A2(KEYINPUT47), .ZN(n561) );
  XOR2_X1 U445 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n490) );
  OR2_X1 U446 ( .A1(G237), .A2(G902), .ZN(n533) );
  XNOR2_X1 U447 ( .A(n501), .B(n433), .ZN(n523) );
  XNOR2_X1 U448 ( .A(n502), .B(KEYINPUT95), .ZN(n433) );
  XOR2_X1 U449 ( .A(KEYINPUT96), .B(KEYINPUT20), .Z(n502) );
  XNOR2_X1 U450 ( .A(n527), .B(G137), .ZN(n446) );
  XNOR2_X1 U451 ( .A(n526), .B(KEYINPUT5), .ZN(n527) );
  XNOR2_X1 U452 ( .A(G116), .B(G146), .ZN(n528) );
  INV_X1 U453 ( .A(KEYINPUT45), .ZN(n457) );
  XNOR2_X1 U454 ( .A(G113), .B(G119), .ZN(n378) );
  XNOR2_X1 U455 ( .A(n377), .B(G101), .ZN(n379) );
  INV_X1 U456 ( .A(KEYINPUT3), .ZN(n377) );
  INV_X1 U457 ( .A(G116), .ZN(n381) );
  AND2_X1 U458 ( .A1(n460), .A2(n741), .ZN(n459) );
  INV_X1 U459 ( .A(n659), .ZN(n460) );
  XNOR2_X1 U460 ( .A(n417), .B(n416), .ZN(n631) );
  XNOR2_X1 U461 ( .A(n496), .B(n729), .ZN(n416) );
  XNOR2_X1 U462 ( .A(n493), .B(n340), .ZN(n417) );
  XNOR2_X1 U463 ( .A(n454), .B(n463), .ZN(n440) );
  NAND2_X2 U464 ( .A1(n408), .A2(n406), .ZN(n663) );
  XOR2_X1 U465 ( .A(KEYINPUT34), .B(KEYINPUT78), .Z(n585) );
  NAND2_X1 U466 ( .A1(n397), .A2(KEYINPUT73), .ZN(n391) );
  XNOR2_X1 U467 ( .A(n499), .B(n419), .ZN(n542) );
  INV_X1 U468 ( .A(KEYINPUT105), .ZN(n419) );
  OR2_X1 U469 ( .A1(n624), .A2(G902), .ZN(n364) );
  NAND2_X1 U470 ( .A1(n353), .A2(n355), .ZN(n352) );
  NOR2_X1 U471 ( .A1(n358), .A2(n582), .ZN(n353) );
  XNOR2_X1 U472 ( .A(n624), .B(KEYINPUT62), .ZN(n625) );
  XNOR2_X1 U473 ( .A(n461), .B(n344), .ZN(n516) );
  XNOR2_X1 U474 ( .A(G134), .B(G122), .ZN(n472) );
  XNOR2_X1 U475 ( .A(n469), .B(n432), .ZN(n447) );
  XNOR2_X1 U476 ( .A(n450), .B(n467), .ZN(n469) );
  XNOR2_X1 U477 ( .A(n468), .B(n470), .ZN(n432) );
  NOR2_X1 U478 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U479 ( .A(n436), .B(n345), .ZN(n742) );
  AND2_X1 U480 ( .A1(n549), .A2(n548), .ZN(n438) );
  NOR2_X1 U481 ( .A1(n558), .A2(n559), .ZN(n443) );
  NAND2_X1 U482 ( .A1(n350), .A2(n349), .ZN(n583) );
  INV_X1 U483 ( .A(n359), .ZN(n349) );
  INV_X1 U484 ( .A(n542), .ZN(n650) );
  AND2_X1 U485 ( .A1(n429), .A2(n430), .ZN(n338) );
  XNOR2_X1 U486 ( .A(n467), .B(KEYINPUT16), .ZN(n339) );
  XOR2_X1 U487 ( .A(n487), .B(n486), .Z(n340) );
  AND2_X1 U488 ( .A1(n431), .A2(n430), .ZN(n341) );
  AND2_X1 U489 ( .A1(n556), .A2(KEYINPUT48), .ZN(n342) );
  INV_X1 U490 ( .A(KEYINPUT1), .ZN(n409) );
  XOR2_X1 U491 ( .A(n532), .B(KEYINPUT109), .Z(n343) );
  XOR2_X1 U492 ( .A(n508), .B(KEYINPUT92), .Z(n344) );
  INV_X1 U493 ( .A(n466), .ZN(n388) );
  XNOR2_X1 U494 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n345) );
  INV_X1 U495 ( .A(KEYINPUT73), .ZN(n399) );
  XNOR2_X1 U496 ( .A(n716), .B(n439), .ZN(n634) );
  XOR2_X1 U497 ( .A(n634), .B(n635), .Z(n346) );
  XOR2_X1 U498 ( .A(n631), .B(n464), .Z(n347) );
  INV_X1 U499 ( .A(KEYINPUT48), .ZN(n448) );
  NOR2_X1 U500 ( .A1(G952), .A2(n732), .ZN(n715) );
  INV_X1 U501 ( .A(n715), .ZN(n430) );
  XNOR2_X1 U502 ( .A(n446), .B(n348), .ZN(n529) );
  INV_X1 U503 ( .A(n385), .ZN(n354) );
  NOR2_X1 U504 ( .A1(n385), .A2(KEYINPUT19), .ZN(n356) );
  NAND2_X1 U505 ( .A1(n363), .A2(n610), .ZN(n614) );
  AND2_X1 U506 ( .A1(n363), .A2(n595), .ZN(n606) );
  XNOR2_X2 U507 ( .A(n364), .B(G472), .ZN(n607) );
  XNOR2_X1 U508 ( .A(n367), .B(n365), .ZN(n624) );
  XNOR2_X2 U509 ( .A(n367), .B(n507), .ZN(n730) );
  XNOR2_X2 U510 ( .A(n376), .B(n374), .ZN(n367) );
  XNOR2_X1 U511 ( .A(n368), .B(n455), .ZN(n454) );
  NOR2_X1 U512 ( .A1(n372), .A2(n666), .ZN(n674) );
  XNOR2_X2 U513 ( .A(n373), .B(G128), .ZN(n475) );
  XNOR2_X2 U514 ( .A(n475), .B(KEYINPUT4), .ZN(n376) );
  XNOR2_X1 U515 ( .A(n376), .B(n440), .ZN(n439) );
  AND2_X1 U516 ( .A1(n411), .A2(n409), .ZN(n407) );
  OR2_X1 U517 ( .A1(n701), .A2(n423), .ZN(n411) );
  XNOR2_X2 U518 ( .A(n730), .B(n447), .ZN(n701) );
  NOR2_X1 U519 ( .A1(n634), .A2(n384), .ZN(n383) );
  NAND2_X1 U520 ( .A1(n634), .A2(n388), .ZN(n387) );
  NOR2_X2 U521 ( .A1(n722), .A2(n389), .ZN(n621) );
  XNOR2_X1 U522 ( .A(n389), .B(n734), .ZN(n733) );
  NAND2_X1 U523 ( .A1(n422), .A2(n459), .ZN(n389) );
  NAND2_X1 U524 ( .A1(n598), .A2(n398), .ZN(n395) );
  NAND2_X1 U525 ( .A1(n392), .A2(n391), .ZN(n562) );
  NAND2_X1 U526 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U527 ( .A1(n540), .A2(n399), .ZN(n393) );
  NAND2_X1 U528 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U529 ( .A(n540), .ZN(n396) );
  NAND2_X1 U530 ( .A1(n598), .A2(n400), .ZN(n397) );
  NAND2_X1 U531 ( .A1(n562), .A2(n435), .ZN(n541) );
  NAND2_X1 U532 ( .A1(n405), .A2(KEYINPUT1), .ZN(n401) );
  NAND2_X1 U533 ( .A1(n402), .A2(n412), .ZN(n421) );
  NAND2_X1 U534 ( .A1(n414), .A2(n415), .ZN(n402) );
  INV_X1 U535 ( .A(n405), .ZN(n410) );
  OR2_X1 U536 ( .A1(n701), .A2(n404), .ZN(n403) );
  NAND2_X1 U537 ( .A1(n410), .A2(n411), .ZN(n548) );
  NAND2_X1 U538 ( .A1(n407), .A2(n410), .ZN(n406) );
  NAND2_X1 U539 ( .A1(n557), .A2(n342), .ZN(n414) );
  XNOR2_X1 U540 ( .A(n547), .B(KEYINPUT46), .ZN(n557) );
  INV_X1 U541 ( .A(n413), .ZN(n415) );
  NAND2_X1 U542 ( .A1(n571), .A2(n572), .ZN(n413) );
  NAND2_X1 U543 ( .A1(n413), .A2(KEYINPUT48), .ZN(n412) );
  NAND2_X1 U544 ( .A1(n421), .A2(n420), .ZN(n422) );
  NAND2_X1 U545 ( .A1(n471), .A2(G902), .ZN(n426) );
  XNOR2_X2 U546 ( .A(n428), .B(n457), .ZN(n722) );
  NAND2_X1 U547 ( .A1(n449), .A2(n458), .ZN(n428) );
  XNOR2_X1 U548 ( .A(n632), .B(n347), .ZN(n429) );
  XNOR2_X1 U549 ( .A(n636), .B(n346), .ZN(n431) );
  NAND2_X1 U550 ( .A1(n705), .A2(G210), .ZN(n636) );
  XNOR2_X2 U551 ( .A(n623), .B(KEYINPUT64), .ZN(n705) );
  NAND2_X1 U552 ( .A1(n435), .A2(n679), .ZN(n682) );
  NOR2_X1 U553 ( .A1(n435), .A2(n679), .ZN(n680) );
  XNOR2_X2 U554 ( .A(n559), .B(KEYINPUT38), .ZN(n435) );
  NAND2_X1 U555 ( .A1(n438), .A2(n678), .ZN(n436) );
  NAND2_X1 U556 ( .A1(n557), .A2(n556), .ZN(n442) );
  XNOR2_X1 U557 ( .A(n443), .B(KEYINPUT36), .ZN(n560) );
  NAND2_X1 U558 ( .A1(n343), .A2(n444), .ZN(n558) );
  NOR2_X1 U559 ( .A1(n542), .A2(n445), .ZN(n444) );
  XNOR2_X1 U560 ( .A(n605), .B(KEYINPUT85), .ZN(n449) );
  XNOR2_X2 U561 ( .A(n517), .B(n456), .ZN(n668) );
  NAND2_X1 U562 ( .A1(n620), .A2(n619), .ZN(n458) );
  XNOR2_X1 U563 ( .A(n703), .B(n702), .ZN(n704) );
  BUF_X1 U564 ( .A(n705), .Z(n711) );
  XNOR2_X2 U565 ( .A(n590), .B(n589), .ZN(n617) );
  AND2_X1 U566 ( .A1(G224), .A2(n732), .ZN(n463) );
  XNOR2_X1 U567 ( .A(KEYINPUT59), .B(KEYINPUT121), .ZN(n464) );
  INV_X1 U568 ( .A(KEYINPUT44), .ZN(n616) );
  XNOR2_X1 U569 ( .A(n538), .B(n537), .ZN(n540) );
  XNOR2_X1 U570 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U571 ( .A(n514), .B(n513), .ZN(n515) );
  INV_X1 U572 ( .A(KEYINPUT63), .ZN(n628) );
  XNOR2_X1 U573 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U574 ( .A(n628), .B(KEYINPUT88), .ZN(n629) );
  XNOR2_X1 U575 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U576 ( .A1(G210), .A2(n533), .ZN(n466) );
  XNOR2_X1 U577 ( .A(G137), .B(G140), .ZN(n507) );
  XNOR2_X1 U578 ( .A(KEYINPUT91), .B(KEYINPUT76), .ZN(n470) );
  NAND2_X1 U579 ( .A1(G227), .A2(n732), .ZN(n468) );
  XNOR2_X1 U580 ( .A(KEYINPUT70), .B(G469), .ZN(n471) );
  XNOR2_X1 U581 ( .A(KEYINPUT104), .B(G478), .ZN(n485) );
  XOR2_X1 U582 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n473) );
  XNOR2_X1 U583 ( .A(n473), .B(n472), .ZN(n483) );
  XOR2_X1 U584 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n477) );
  XNOR2_X1 U585 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U586 ( .A(n477), .B(n476), .ZN(n481) );
  NAND2_X1 U587 ( .A1(n732), .A2(G234), .ZN(n479) );
  XNOR2_X1 U588 ( .A(n479), .B(n478), .ZN(n512) );
  NAND2_X1 U589 ( .A1(n512), .A2(G217), .ZN(n480) );
  XOR2_X1 U590 ( .A(n481), .B(n480), .Z(n482) );
  XNOR2_X1 U591 ( .A(n483), .B(n482), .ZN(n706) );
  NOR2_X1 U592 ( .A1(G902), .A2(n706), .ZN(n484) );
  XNOR2_X1 U593 ( .A(n485), .B(n484), .ZN(n563) );
  XNOR2_X1 U594 ( .A(n488), .B(KEYINPUT72), .ZN(n530) );
  NAND2_X1 U595 ( .A1(n530), .A2(G214), .ZN(n492) );
  XNOR2_X1 U596 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U597 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U599 ( .A(KEYINPUT13), .B(G475), .ZN(n497) );
  XNOR2_X1 U600 ( .A(n498), .B(n497), .ZN(n552) );
  NAND2_X1 U601 ( .A1(n563), .A2(n552), .ZN(n499) );
  XOR2_X1 U602 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n504) );
  INV_X1 U603 ( .A(n500), .ZN(n622) );
  NAND2_X1 U604 ( .A1(G234), .A2(n622), .ZN(n501) );
  NAND2_X1 U605 ( .A1(G217), .A2(n523), .ZN(n503) );
  XNOR2_X1 U606 ( .A(n506), .B(n505), .ZN(n509) );
  INV_X1 U607 ( .A(n507), .ZN(n508) );
  XOR2_X1 U608 ( .A(n511), .B(n510), .Z(n514) );
  NAND2_X1 U609 ( .A1(G221), .A2(n512), .ZN(n513) );
  XNOR2_X1 U610 ( .A(n516), .B(n515), .ZN(n710) );
  NOR2_X1 U611 ( .A1(G902), .A2(n710), .ZN(n517) );
  NAND2_X1 U612 ( .A1(G234), .A2(G237), .ZN(n518) );
  XNOR2_X1 U613 ( .A(n518), .B(KEYINPUT90), .ZN(n519) );
  XNOR2_X1 U614 ( .A(KEYINPUT14), .B(n519), .ZN(n520) );
  NAND2_X1 U615 ( .A1(G952), .A2(n520), .ZN(n693) );
  NOR2_X1 U616 ( .A1(G953), .A2(n693), .ZN(n581) );
  AND2_X1 U617 ( .A1(n520), .A2(G953), .ZN(n521) );
  NAND2_X1 U618 ( .A1(G902), .A2(n521), .ZN(n579) );
  NOR2_X1 U619 ( .A1(G900), .A2(n579), .ZN(n522) );
  NAND2_X1 U620 ( .A1(n523), .A2(G221), .ZN(n524) );
  XNOR2_X1 U621 ( .A(n524), .B(KEYINPUT21), .ZN(n669) );
  NOR2_X1 U622 ( .A1(n539), .A2(n669), .ZN(n525) );
  NAND2_X1 U623 ( .A1(n668), .A2(n525), .ZN(n546) );
  INV_X1 U624 ( .A(KEYINPUT98), .ZN(n526) );
  NAND2_X1 U625 ( .A1(G210), .A2(n530), .ZN(n531) );
  XNOR2_X1 U626 ( .A(n607), .B(KEYINPUT6), .ZN(n609) );
  NOR2_X1 U627 ( .A1(n546), .A2(n609), .ZN(n532) );
  NAND2_X1 U628 ( .A1(G214), .A2(n533), .ZN(n679) );
  NOR2_X1 U629 ( .A1(n663), .A2(n558), .ZN(n534) );
  XNOR2_X1 U630 ( .A(n534), .B(KEYINPUT43), .ZN(n535) );
  NOR2_X1 U631 ( .A1(n566), .A2(n535), .ZN(n659) );
  INV_X1 U632 ( .A(KEYINPUT30), .ZN(n536) );
  XOR2_X1 U633 ( .A(KEYINPUT97), .B(n669), .Z(n592) );
  AND2_X1 U634 ( .A1(n548), .A2(n664), .ZN(n598) );
  INV_X1 U635 ( .A(n566), .ZN(n559) );
  NAND2_X1 U636 ( .A1(n573), .A2(n650), .ZN(n544) );
  XOR2_X1 U637 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n543) );
  XNOR2_X1 U638 ( .A(n544), .B(n543), .ZN(n739) );
  INV_X1 U639 ( .A(n552), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n563), .A2(n564), .ZN(n681) );
  INV_X1 U641 ( .A(n607), .ZN(n666) );
  NAND2_X1 U642 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U643 ( .A1(n550), .A2(n583), .ZN(n553) );
  NAND2_X1 U644 ( .A1(KEYINPUT66), .A2(n553), .ZN(n551) );
  XNOR2_X1 U645 ( .A(n551), .B(KEYINPUT47), .ZN(n555) );
  NOR2_X1 U646 ( .A1(n552), .A2(n563), .ZN(n654) );
  NAND2_X1 U647 ( .A1(n683), .A2(n553), .ZN(n554) );
  NAND2_X1 U648 ( .A1(n555), .A2(n554), .ZN(n556) );
  INV_X1 U649 ( .A(n663), .ZN(n595) );
  XNOR2_X1 U650 ( .A(KEYINPUT87), .B(n595), .ZN(n611) );
  NAND2_X1 U651 ( .A1(n560), .A2(n611), .ZN(n658) );
  XNOR2_X1 U652 ( .A(n658), .B(KEYINPUT84), .ZN(n572) );
  XNOR2_X1 U653 ( .A(KEYINPUT81), .B(n561), .ZN(n569) );
  INV_X1 U654 ( .A(n562), .ZN(n568) );
  NOR2_X1 U655 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U656 ( .A(n565), .B(KEYINPUT108), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n566), .A2(n587), .ZN(n567) );
  NOR2_X1 U658 ( .A1(n568), .A2(n567), .ZN(n648) );
  NOR2_X1 U659 ( .A1(n569), .A2(n648), .ZN(n570) );
  XNOR2_X1 U660 ( .A(n570), .B(KEYINPUT80), .ZN(n571) );
  NAND2_X1 U661 ( .A1(n573), .A2(n654), .ZN(n574) );
  XNOR2_X1 U662 ( .A(KEYINPUT114), .B(n574), .ZN(n741) );
  XNOR2_X1 U663 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n576) );
  INV_X1 U664 ( .A(KEYINPUT107), .ZN(n575) );
  XNOR2_X1 U665 ( .A(n578), .B(n577), .ZN(n660) );
  NOR2_X1 U666 ( .A1(G898), .A2(n579), .ZN(n580) );
  NOR2_X1 U667 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U668 ( .A1(n660), .A2(n599), .ZN(n586) );
  XNOR2_X1 U669 ( .A(n586), .B(n585), .ZN(n588) );
  NAND2_X1 U670 ( .A1(n588), .A2(n587), .ZN(n590) );
  XOR2_X1 U671 ( .A(KEYINPUT35), .B(KEYINPUT77), .Z(n589) );
  NAND2_X1 U672 ( .A1(n617), .A2(KEYINPUT44), .ZN(n591) );
  XNOR2_X1 U673 ( .A(n591), .B(KEYINPUT86), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n681), .A2(n592), .ZN(n593) );
  NAND2_X1 U675 ( .A1(n599), .A2(n593), .ZN(n594) );
  NAND2_X1 U676 ( .A1(n606), .A2(n609), .ZN(n596) );
  NOR2_X1 U677 ( .A1(n668), .A2(n596), .ZN(n638) );
  NAND2_X1 U678 ( .A1(n599), .A2(n674), .ZN(n597) );
  XNOR2_X1 U679 ( .A(n597), .B(KEYINPUT31), .ZN(n655) );
  NAND2_X1 U680 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n607), .A2(n600), .ZN(n641) );
  NOR2_X1 U682 ( .A1(n655), .A2(n641), .ZN(n601) );
  NOR2_X1 U683 ( .A1(n683), .A2(n601), .ZN(n602) );
  NOR2_X1 U684 ( .A1(n638), .A2(n602), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n668), .A2(n606), .ZN(n608) );
  NOR2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n645) );
  XOR2_X1 U688 ( .A(KEYINPUT79), .B(n609), .Z(n610) );
  NAND2_X1 U689 ( .A1(n668), .A2(n611), .ZN(n612) );
  XNOR2_X1 U690 ( .A(KEYINPUT106), .B(n612), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U692 ( .A(KEYINPUT32), .B(n615), .ZN(n743) );
  XNOR2_X1 U693 ( .A(n618), .B(n616), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT2), .ZN(n661) );
  NOR2_X2 U696 ( .A1(n661), .A2(n622), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n705), .A2(G472), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X2 U699 ( .A1(n627), .A2(n715), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(G57) );
  NAND2_X1 U701 ( .A1(G475), .A2(n705), .ZN(n632) );
  XOR2_X1 U702 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n633) );
  XNOR2_X1 U703 ( .A(n338), .B(n633), .ZN(G60) );
  XOR2_X1 U704 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT83), .B(KEYINPUT56), .Z(n637) );
  XNOR2_X1 U706 ( .A(n341), .B(n637), .ZN(G51) );
  XOR2_X1 U707 ( .A(G101), .B(n638), .Z(G3) );
  XOR2_X1 U708 ( .A(G104), .B(KEYINPUT115), .Z(n640) );
  NAND2_X1 U709 ( .A1(n641), .A2(n650), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(G6) );
  XOR2_X1 U711 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n643) );
  NAND2_X1 U712 ( .A1(n641), .A2(n654), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(G107), .B(n644), .ZN(G9) );
  XOR2_X1 U715 ( .A(n645), .B(G110), .Z(G12) );
  XOR2_X1 U716 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  NAND2_X1 U717 ( .A1(n553), .A2(n654), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(G30) );
  XOR2_X1 U719 ( .A(G143), .B(n648), .Z(G45) );
  NAND2_X1 U720 ( .A1(n553), .A2(n650), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n649), .B(G146), .ZN(G48) );
  XOR2_X1 U722 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n652) );
  NAND2_X1 U723 ( .A1(n655), .A2(n650), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(G113), .B(n653), .ZN(G15) );
  NAND2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(G116), .ZN(G18) );
  XOR2_X1 U728 ( .A(G125), .B(KEYINPUT37), .Z(n657) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(G27) );
  XOR2_X1 U730 ( .A(G140), .B(n659), .Z(G42) );
  BUF_X1 U731 ( .A(n660), .Z(n687) );
  NAND2_X1 U732 ( .A1(n687), .A2(n678), .ZN(n697) );
  BUF_X1 U733 ( .A(n661), .Z(n662) );
  NAND2_X1 U734 ( .A1(n732), .A2(n662), .ZN(n695) );
  XNOR2_X1 U735 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n691) );
  XNOR2_X1 U736 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n676) );
  OR2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(KEYINPUT50), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n672) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U741 ( .A(KEYINPUT49), .B(n670), .ZN(n671) );
  NOR2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n689) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  OR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U750 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U751 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U752 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(KEYINPUT53), .ZN(n699) );
  XOR2_X1 U755 ( .A(KEYINPUT120), .B(n699), .Z(G75) );
  NAND2_X1 U756 ( .A1(G469), .A2(n711), .ZN(n703) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n700) );
  NOR2_X1 U758 ( .A1(n715), .A2(n704), .ZN(G54) );
  NAND2_X1 U759 ( .A1(n711), .A2(G478), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n706), .B(KEYINPUT122), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n715), .A2(n709), .ZN(G63) );
  BUF_X1 U762 ( .A(n710), .Z(n713) );
  NAND2_X1 U763 ( .A1(G217), .A2(n711), .ZN(n712) );
  XNOR2_X1 U764 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U765 ( .A1(n715), .A2(n714), .ZN(G66) );
  XNOR2_X1 U766 ( .A(KEYINPUT125), .B(n716), .ZN(n718) );
  NOR2_X1 U767 ( .A1(n732), .A2(G898), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n728) );
  NAND2_X1 U769 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U770 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n720), .A2(G898), .ZN(n721) );
  XNOR2_X1 U772 ( .A(KEYINPUT123), .B(n721), .ZN(n725) );
  NOR2_X1 U773 ( .A1(G953), .A2(n722), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n723), .B(KEYINPUT124), .ZN(n724) );
  NOR2_X1 U775 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U776 ( .A(n726), .B(KEYINPUT126), .Z(n727) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(G69) );
  XOR2_X1 U778 ( .A(n730), .B(n729), .Z(n731) );
  XNOR2_X1 U779 ( .A(KEYINPUT127), .B(n731), .ZN(n734) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(n738) );
  XNOR2_X1 U781 ( .A(G227), .B(n734), .ZN(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(G900), .ZN(n736) );
  NAND2_X1 U783 ( .A1(G953), .A2(n736), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n738), .A2(n737), .ZN(G72) );
  BUF_X1 U785 ( .A(n739), .Z(n740) );
  XOR2_X1 U786 ( .A(G131), .B(n740), .Z(G33) );
  XOR2_X1 U787 ( .A(n617), .B(G122), .Z(G24) );
  XNOR2_X1 U788 ( .A(G134), .B(n741), .ZN(G36) );
  XOR2_X1 U789 ( .A(G137), .B(n742), .Z(G39) );
  XOR2_X1 U790 ( .A(G119), .B(n743), .Z(G21) );
endmodule

