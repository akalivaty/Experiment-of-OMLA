

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U324 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U325 ( .A1(n559), .A2(n558), .ZN(n292) );
  XNOR2_X1 U326 ( .A(KEYINPUT108), .B(KEYINPUT47), .ZN(n408) );
  XNOR2_X1 U327 ( .A(n409), .B(n408), .ZN(n415) );
  XNOR2_X1 U328 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U329 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U330 ( .A(n454), .B(n453), .ZN(n560) );
  XOR2_X1 U331 ( .A(n464), .B(KEYINPUT28), .Z(n530) );
  XNOR2_X1 U332 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G120GAT), .B(G71GAT), .Z(n365) );
  XOR2_X1 U335 ( .A(G15GAT), .B(G127GAT), .Z(n401) );
  XNOR2_X1 U336 ( .A(n365), .B(n401), .ZN(n294) );
  XNOR2_X1 U337 ( .A(G113GAT), .B(G134GAT), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n293), .B(KEYINPUT0), .ZN(n324) );
  XNOR2_X1 U339 ( .A(n294), .B(n324), .ZN(n300) );
  XOR2_X1 U340 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n419) );
  XOR2_X1 U343 ( .A(n419), .B(G176GAT), .Z(n298) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U346 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U347 ( .A(KEYINPUT64), .B(G99GAT), .Z(n302) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U350 ( .A(G183GAT), .B(KEYINPUT82), .Z(n304) );
  XNOR2_X1 U351 ( .A(KEYINPUT83), .B(KEYINPUT20), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n459) );
  NAND2_X1 U355 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XOR2_X1 U356 ( .A(G155GAT), .B(G148GAT), .Z(n310) );
  XNOR2_X1 U357 ( .A(G29GAT), .B(G120GAT), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n312) );
  XOR2_X1 U359 ( .A(G162GAT), .B(G85GAT), .Z(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n330) );
  XOR2_X1 U362 ( .A(KEYINPUT6), .B(KEYINPUT87), .Z(n316) );
  XNOR2_X1 U363 ( .A(KEYINPUT4), .B(KEYINPUT91), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n328) );
  XOR2_X1 U365 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n318) );
  XNOR2_X1 U366 ( .A(G127GAT), .B(KEYINPUT89), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U368 ( .A(G57GAT), .B(KEYINPUT1), .Z(n320) );
  XNOR2_X1 U369 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U371 ( .A(n322), .B(n321), .Z(n326) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n323), .B(KEYINPUT2), .ZN(n439) );
  XNOR2_X1 U374 ( .A(n324), .B(n439), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U376 ( .A(n328), .B(n327), .Z(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n514) );
  XOR2_X1 U378 ( .A(KEYINPUT67), .B(G8GAT), .Z(n332) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(G113GAT), .ZN(n331) );
  XNOR2_X1 U380 ( .A(n332), .B(n331), .ZN(n349) );
  XOR2_X1 U381 ( .A(G197GAT), .B(G141GAT), .Z(n334) );
  XNOR2_X1 U382 ( .A(G169GAT), .B(G22GAT), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n334), .B(n333), .ZN(n336) );
  XOR2_X1 U384 ( .A(G50GAT), .B(G36GAT), .Z(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n345) );
  XNOR2_X1 U386 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n337), .B(KEYINPUT29), .ZN(n338) );
  XOR2_X1 U388 ( .A(n338), .B(KEYINPUT66), .Z(n343) );
  XOR2_X1 U389 ( .A(G29GAT), .B(G43GAT), .Z(n340) );
  XNOR2_X1 U390 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n384) );
  XNOR2_X1 U392 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n341), .B(KEYINPUT70), .ZN(n402) );
  XNOR2_X1 U394 ( .A(n384), .B(n402), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n347) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n556) );
  XNOR2_X1 U400 ( .A(G99GAT), .B(G85GAT), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n350), .B(KEYINPUT72), .ZN(n383) );
  INV_X1 U402 ( .A(n383), .ZN(n351) );
  NAND2_X1 U403 ( .A1(n351), .A2(KEYINPUT33), .ZN(n354) );
  INV_X1 U404 ( .A(KEYINPUT33), .ZN(n352) );
  NAND2_X1 U405 ( .A1(n352), .A2(n383), .ZN(n353) );
  NAND2_X1 U406 ( .A1(n354), .A2(n353), .ZN(n356) );
  NAND2_X1 U407 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U409 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n358) );
  XNOR2_X1 U410 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n357) );
  XOR2_X1 U411 ( .A(n358), .B(n357), .Z(n359) );
  XNOR2_X1 U412 ( .A(n360), .B(n359), .ZN(n368) );
  XOR2_X1 U413 ( .A(G78GAT), .B(G148GAT), .Z(n362) );
  XNOR2_X1 U414 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n440) );
  XOR2_X1 U416 ( .A(G64GAT), .B(G92GAT), .Z(n364) );
  XNOR2_X1 U417 ( .A(G176GAT), .B(G204GAT), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n420) );
  XNOR2_X1 U419 ( .A(n440), .B(n420), .ZN(n366) );
  XOR2_X1 U420 ( .A(G57GAT), .B(KEYINPUT13), .Z(n391) );
  XNOR2_X1 U421 ( .A(n369), .B(n391), .ZN(n575) );
  XNOR2_X1 U422 ( .A(KEYINPUT41), .B(n575), .ZN(n558) );
  AND2_X1 U423 ( .A1(n556), .A2(n558), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n370), .B(KEYINPUT46), .ZN(n387) );
  XOR2_X1 U425 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n372) );
  XNOR2_X1 U426 ( .A(G106GAT), .B(G92GAT), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U428 ( .A(G36GAT), .B(G190GAT), .Z(n421) );
  XOR2_X1 U429 ( .A(KEYINPUT77), .B(n421), .Z(n374) );
  XOR2_X1 U430 ( .A(G50GAT), .B(G162GAT), .Z(n446) );
  XNOR2_X1 U431 ( .A(n446), .B(G218GAT), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U433 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U434 ( .A1(G232GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U436 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n380) );
  XNOR2_X1 U437 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U439 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n553) );
  NOR2_X1 U442 ( .A1(n387), .A2(n553), .ZN(n407) );
  XOR2_X1 U443 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n389) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT15), .B(n390), .ZN(n406) );
  XOR2_X1 U447 ( .A(G8GAT), .B(G183GAT), .Z(n425) );
  XOR2_X1 U448 ( .A(n425), .B(n391), .Z(n393) );
  XNOR2_X1 U449 ( .A(G78GAT), .B(G211GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U451 ( .A(n394), .B(KEYINPUT79), .Z(n399) );
  XOR2_X1 U452 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n396) );
  XNOR2_X1 U453 ( .A(G64GAT), .B(KEYINPUT78), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(G71GAT), .B(n397), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U457 ( .A(G22GAT), .B(G155GAT), .Z(n445) );
  XOR2_X1 U458 ( .A(n400), .B(n445), .Z(n404) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n579) );
  NAND2_X1 U462 ( .A1(n407), .A2(n579), .ZN(n409) );
  XNOR2_X1 U463 ( .A(KEYINPUT36), .B(KEYINPUT99), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n553), .B(n410), .ZN(n585) );
  NOR2_X1 U465 ( .A1(n585), .A2(n579), .ZN(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT45), .B(n411), .ZN(n412) );
  NAND2_X1 U467 ( .A1(n412), .A2(n575), .ZN(n413) );
  NOR2_X1 U468 ( .A1(n556), .A2(n413), .ZN(n414) );
  NOR2_X1 U469 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n416), .B(KEYINPUT48), .ZN(n527) );
  XOR2_X1 U471 ( .A(G211GAT), .B(KEYINPUT21), .Z(n418) );
  XNOR2_X1 U472 ( .A(G197GAT), .B(G218GAT), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n443) );
  XNOR2_X1 U474 ( .A(n419), .B(n443), .ZN(n429) );
  XOR2_X1 U475 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U476 ( .A1(G226GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U478 ( .A(n424), .B(KEYINPUT93), .Z(n427) );
  XNOR2_X1 U479 ( .A(n425), .B(KEYINPUT92), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n517) );
  XOR2_X1 U482 ( .A(KEYINPUT118), .B(n517), .Z(n430) );
  NOR2_X1 U483 ( .A1(n527), .A2(n430), .ZN(n432) );
  INV_X1 U484 ( .A(KEYINPUT54), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n433) );
  NOR2_X1 U486 ( .A1(n514), .A2(n433), .ZN(n569) );
  XOR2_X1 U487 ( .A(G204GAT), .B(KEYINPUT85), .Z(n435) );
  XNOR2_X1 U488 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n450) );
  XOR2_X1 U490 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n437) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U493 ( .A(n438), .B(KEYINPUT24), .Z(n442) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U496 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U499 ( .A(n450), .B(n449), .Z(n464) );
  NAND2_X1 U500 ( .A1(n569), .A2(n464), .ZN(n454) );
  XOR2_X1 U501 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n452) );
  INV_X1 U502 ( .A(KEYINPUT55), .ZN(n451) );
  NOR2_X1 U503 ( .A1(n459), .A2(n560), .ZN(n565) );
  NAND2_X1 U504 ( .A1(n565), .A2(n553), .ZN(n458) );
  XOR2_X1 U505 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n456) );
  INV_X1 U506 ( .A(G190GAT), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n517), .B(KEYINPUT27), .ZN(n466) );
  NAND2_X1 U508 ( .A1(n514), .A2(n466), .ZN(n526) );
  INV_X1 U509 ( .A(n459), .ZN(n559) );
  OR2_X1 U510 ( .A1(n559), .A2(n530), .ZN(n460) );
  NOR2_X1 U511 ( .A1(n526), .A2(n460), .ZN(n471) );
  NAND2_X1 U512 ( .A1(n517), .A2(n559), .ZN(n461) );
  XNOR2_X1 U513 ( .A(KEYINPUT94), .B(n461), .ZN(n462) );
  NAND2_X1 U514 ( .A1(n462), .A2(n464), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n463), .B(KEYINPUT25), .ZN(n468) );
  NOR2_X1 U516 ( .A1(n464), .A2(n559), .ZN(n465) );
  XNOR2_X1 U517 ( .A(KEYINPUT26), .B(n465), .ZN(n568) );
  AND2_X1 U518 ( .A1(n466), .A2(n568), .ZN(n467) );
  NOR2_X1 U519 ( .A1(n468), .A2(n467), .ZN(n469) );
  NOR2_X1 U520 ( .A1(n514), .A2(n469), .ZN(n470) );
  NOR2_X1 U521 ( .A1(n471), .A2(n470), .ZN(n472) );
  XOR2_X1 U522 ( .A(KEYINPUT95), .B(n472), .Z(n487) );
  NOR2_X1 U523 ( .A1(n553), .A2(n579), .ZN(n473) );
  XOR2_X1 U524 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U525 ( .A1(n487), .A2(n474), .ZN(n475) );
  XOR2_X1 U526 ( .A(KEYINPUT96), .B(n475), .Z(n500) );
  NAND2_X1 U527 ( .A1(n556), .A2(n575), .ZN(n476) );
  XNOR2_X1 U528 ( .A(n476), .B(KEYINPUT75), .ZN(n490) );
  INV_X1 U529 ( .A(n490), .ZN(n477) );
  NOR2_X1 U530 ( .A1(n500), .A2(n477), .ZN(n485) );
  NAND2_X1 U531 ( .A1(n485), .A2(n514), .ZN(n481) );
  XOR2_X1 U532 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n479) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U535 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U536 ( .A1(n485), .A2(n517), .ZN(n482) );
  XNOR2_X1 U537 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U539 ( .A1(n485), .A2(n559), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NAND2_X1 U541 ( .A1(n485), .A2(n530), .ZN(n486) );
  XNOR2_X1 U542 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT38), .B(KEYINPUT100), .Z(n492) );
  NOR2_X1 U544 ( .A1(n585), .A2(n487), .ZN(n488) );
  NAND2_X1 U545 ( .A1(n579), .A2(n488), .ZN(n489) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n489), .ZN(n511) );
  NAND2_X1 U547 ( .A1(n490), .A2(n511), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n492), .B(n491), .ZN(n498) );
  NAND2_X1 U549 ( .A1(n514), .A2(n498), .ZN(n494) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  XNOR2_X1 U551 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n498), .A2(n517), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n559), .A2(n498), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n530), .A2(n498), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT101), .B(KEYINPUT42), .Z(n502) );
  INV_X1 U560 ( .A(n556), .ZN(n570) );
  NAND2_X1 U561 ( .A1(n558), .A2(n570), .ZN(n510) );
  NOR2_X1 U562 ( .A1(n500), .A2(n510), .ZN(n507) );
  NAND2_X1 U563 ( .A1(n507), .A2(n514), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n507), .A2(n517), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n559), .A2(n507), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT102), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U572 ( .A1(n507), .A2(n530), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT104), .ZN(n516) );
  INV_X1 U575 ( .A(n510), .ZN(n512) );
  NAND2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT103), .ZN(n523) );
  NAND2_X1 U578 ( .A1(n514), .A2(n523), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n519) );
  NAND2_X1 U581 ( .A1(n523), .A2(n517), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  XOR2_X1 U584 ( .A(G99GAT), .B(KEYINPUT107), .Z(n522) );
  NAND2_X1 U585 ( .A1(n523), .A2(n559), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n530), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT110), .ZN(n532) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n543), .A2(n559), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT109), .B(n528), .Z(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n539), .A2(n556), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n534) );
  NAND2_X1 U598 ( .A1(n539), .A2(n558), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT111), .Z(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  INV_X1 U602 ( .A(n579), .ZN(n566) );
  NAND2_X1 U603 ( .A1(n566), .A2(n539), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U607 ( .A1(n539), .A2(n553), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U609 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT115), .Z(n546) );
  NAND2_X1 U611 ( .A1(n568), .A2(n543), .ZN(n544) );
  XOR2_X1 U612 ( .A(KEYINPUT114), .B(n544), .Z(n552) );
  NAND2_X1 U613 ( .A1(n552), .A2(n556), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U616 ( .A1(n552), .A2(n558), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n566), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n550), .B(KEYINPUT116), .ZN(n551) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(G162GAT), .B(KEYINPUT117), .Z(n555) );
  NAND2_X1 U623 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n565), .A2(n556), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT57), .Z(n562) );
  OR2_X1 U628 ( .A1(n292), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n584) );
  NOR2_X1 U635 ( .A1(n570), .A2(n584), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n584), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT61), .B(KEYINPUT124), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n584), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n583) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

