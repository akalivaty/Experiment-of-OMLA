//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  NAND2_X1  g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT90), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n204), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT91), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT14), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n206), .A2(new_n207), .A3(new_n209), .A4(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G43gat), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  NAND2_X1  g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n206), .A2(new_n209), .A3(new_n212), .A4(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n216), .B2(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n213), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  AND4_X1   g022(.A1(new_n205), .A2(new_n212), .A3(new_n203), .A4(new_n209), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(new_n219), .C1(new_n221), .C2(new_n207), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n230), .A2(G1gat), .ZN(new_n231));
  AOI21_X1  g030(.A(G8gat), .B1(new_n231), .B2(KEYINPUT93), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT92), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OR3_X1    g033(.A1(new_n233), .A2(new_n234), .A3(G1gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(G1gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n231), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n232), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT94), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n226), .B2(KEYINPUT17), .ZN(new_n241));
  AOI211_X1 g040(.A(KEYINPUT94), .B(new_n228), .C1(new_n223), .C2(new_n225), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n229), .B(new_n239), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n239), .A2(new_n226), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n247), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n239), .B(new_n226), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n244), .B(KEYINPUT13), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT11), .ZN(new_n255));
  INV_X1    g054(.A(G169gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G197gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n248), .A2(new_n249), .A3(new_n252), .A4(new_n259), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n265));
  XNOR2_X1  g064(.A(G1gat), .B(G29gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT0), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n270), .A2(KEYINPUT68), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(KEYINPUT68), .ZN(new_n272));
  INV_X1    g071(.A(G120gat), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n273), .A2(G113gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(G113gat), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n271), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT69), .B(G113gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G120gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n275), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n270), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT1), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n277), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n285), .A2(KEYINPUT81), .ZN(new_n286));
  XNOR2_X1  g085(.A(G141gat), .B(G148gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G155gat), .ZN(new_n290));
  INV_X1    g089(.A(G162gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n295), .B2(KEYINPUT2), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n293), .B(new_n295), .C1(new_n287), .C2(KEYINPUT2), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n299), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT80), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n285), .A2(KEYINPUT81), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n286), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n302), .A2(KEYINPUT82), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT82), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n297), .A2(new_n310), .A3(new_n299), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(KEYINPUT4), .A3(new_n285), .ZN(new_n313));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n302), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n285), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n308), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n286), .A2(new_n302), .A3(new_n306), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n321), .A2(new_n317), .ZN(new_n322));
  OAI211_X1 g121(.A(KEYINPUT5), .B(new_n320), .C1(new_n322), .C2(new_n314), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n285), .A2(new_n309), .A3(new_n311), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT83), .B1(new_n324), .B2(KEYINPUT4), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT83), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n312), .A2(new_n326), .A3(new_n318), .A4(new_n285), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n317), .A2(KEYINPUT4), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n315), .A2(KEYINPUT5), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n308), .A3(new_n330), .ZN(new_n331));
  AOI211_X1 g130(.A(new_n265), .B(new_n269), .C1(new_n323), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n320), .A2(KEYINPUT5), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n314), .B1(new_n321), .B2(new_n317), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n269), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n323), .A2(new_n269), .A3(new_n331), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n265), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n332), .B1(new_n339), .B2(KEYINPUT89), .ZN(new_n340));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT22), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT74), .B(G218gat), .ZN(new_n346));
  INV_X1    g145(.A(G211gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(G211gat), .B(G218gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  OR2_X1    g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(KEYINPUT24), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G176gat), .ZN(new_n360));
  OAI221_X1 g159(.A(new_n359), .B1(KEYINPUT24), .B2(new_n358), .C1(new_n256), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT64), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT23), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT25), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(KEYINPUT65), .A3(KEYINPUT25), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n365), .A2(KEYINPUT25), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT27), .B(G183gat), .ZN(new_n372));
  INV_X1    g171(.A(G190gat), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT66), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(KEYINPUT28), .ZN(new_n375));
  OR3_X1    g174(.A1(new_n375), .A2(new_n374), .A3(KEYINPUT28), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n374), .B2(KEYINPUT28), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n256), .A2(new_n360), .A3(KEYINPUT67), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n256), .A2(new_n360), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(KEYINPUT26), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(KEYINPUT26), .B2(new_n378), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n376), .A2(new_n377), .A3(new_n358), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n356), .B1(new_n371), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(KEYINPUT76), .B(KEYINPUT29), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n371), .B2(new_n382), .ZN(new_n386));
  INV_X1    g185(.A(new_n356), .ZN(new_n387));
  OAI22_X1  g186(.A1(KEYINPUT77), .A2(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n383), .A2(KEYINPUT77), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n355), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n382), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n356), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n383), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n383), .A2(new_n395), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n394), .B(new_n354), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n390), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT37), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n344), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n383), .A2(new_n395), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n395), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n402), .A2(new_n403), .B1(new_n356), .B2(new_n393), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n404), .B2(new_n355), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n354), .B1(new_n388), .B2(new_n389), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT38), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n401), .A2(new_n407), .B1(new_n399), .B2(new_n344), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT6), .B1(new_n335), .B2(new_n336), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT89), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n338), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n399), .A2(new_n400), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n398), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n343), .B1(new_n413), .B2(KEYINPUT37), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT38), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n340), .A2(new_n408), .A3(new_n411), .A4(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n354), .A2(new_n384), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n312), .B1(new_n420), .B2(new_n298), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n354), .B1(new_n300), .B2(new_n384), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n300), .A2(new_n384), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT84), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n419), .B1(new_n425), .B2(new_n355), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n354), .B2(new_n392), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n316), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G22gat), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n423), .B2(new_n428), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n418), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n423), .A2(new_n428), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G22gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n417), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT31), .B(G50gat), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n432), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n432), .B2(new_n436), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n329), .A2(new_n308), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(new_n315), .ZN(new_n444));
  AOI211_X1 g243(.A(KEYINPUT87), .B(new_n314), .C1(new_n329), .C2(new_n308), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n321), .A2(new_n314), .A3(new_n317), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n447), .A2(KEYINPUT88), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(KEYINPUT88), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n444), .B2(new_n445), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n269), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT40), .A4(new_n269), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n337), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n390), .A2(new_n398), .A3(new_n460), .A4(new_n344), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n390), .A2(new_n398), .A3(new_n344), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT30), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n344), .B1(new_n390), .B2(new_n398), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n459), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n413), .A2(new_n343), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(KEYINPUT30), .A3(new_n462), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n459), .B1(new_n468), .B2(new_n461), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n416), .B(new_n441), .C1(new_n458), .C2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n430), .A2(new_n431), .A3(new_n418), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n417), .B1(new_n434), .B2(new_n435), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n437), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n432), .A2(new_n436), .A3(new_n438), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n335), .A2(KEYINPUT6), .A3(new_n336), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n339), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n468), .A2(new_n461), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n475), .A2(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n391), .A2(new_n285), .ZN(new_n481));
  INV_X1    g280(.A(new_n285), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n371), .A2(new_n482), .A3(new_n382), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n481), .A2(G227gat), .A3(G233gat), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT32), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G43gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT71), .ZN(new_n489));
  XOR2_X1   g288(.A(G71gat), .B(G99gat), .Z(new_n490));
  XOR2_X1   g289(.A(new_n489), .B(new_n490), .Z(new_n491));
  NAND3_X1  g290(.A1(new_n485), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n483), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n482), .B1(new_n371), .B2(new_n382), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n497), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n493), .B(new_n499), .C1(new_n494), .C2(new_n495), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n491), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n484), .B(KEYINPUT32), .C1(new_n486), .C2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n492), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n492), .B2(new_n503), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n501), .A3(new_n503), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n503), .ZN(new_n511));
  INV_X1    g310(.A(new_n501), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n492), .A2(new_n501), .A3(KEYINPUT73), .A4(new_n503), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n507), .B1(new_n506), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n472), .B1(new_n480), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n478), .A2(new_n479), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n439), .B2(new_n440), .ZN(new_n519));
  INV_X1    g318(.A(new_n507), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(KEYINPUT36), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT85), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n471), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n475), .A2(new_n476), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n504), .A2(new_n505), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n525), .A2(new_n518), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n340), .A2(new_n411), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n470), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n521), .A2(new_n475), .A3(new_n529), .A4(new_n476), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n264), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  OR3_X1    g333(.A1(KEYINPUT95), .A2(G71gat), .A3(G78gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT95), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G57gat), .ZN(new_n539));
  INV_X1    g338(.A(G64gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G57gat), .A2(G64gat), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n541), .A2(KEYINPUT9), .A3(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G71gat), .ZN(new_n545));
  INV_X1    g344(.A(G78gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT9), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n536), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n549));
  AND2_X1   g348(.A1(G57gat), .A2(G64gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(G57gat), .A2(G64gat), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n541), .A2(KEYINPUT96), .A3(new_n542), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n548), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n548), .A2(new_n552), .A3(new_n553), .A4(KEYINPUT97), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n544), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n239), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n557), .ZN(new_n562));
  INV_X1    g361(.A(new_n544), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n566), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n569), .A2(new_n571), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n561), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n569), .A2(new_n571), .ZN(new_n576));
  INV_X1    g375(.A(new_n561), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n560), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n560), .A3(new_n578), .ZN(new_n581));
  XOR2_X1   g380(.A(G183gat), .B(G211gat), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n575), .A2(new_n560), .A3(new_n578), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n582), .B1(new_n585), .B2(new_n579), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT41), .ZN(new_n590));
  NAND3_X1  g389(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(KEYINPUT98), .A2(G99gat), .A3(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT98), .B1(G99gat), .B2(G106gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT8), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  OR2_X1    g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n595), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n600), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n594), .A2(new_n593), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n591), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT8), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n608), .B2(new_n596), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n603), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT99), .B1(new_n602), .B2(new_n610), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n229), .B(new_n615), .C1(new_n241), .C2(new_n242), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n611), .B(new_n612), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n617), .A2(new_n227), .B1(KEYINPUT41), .B2(new_n589), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n616), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n616), .B2(new_n618), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n590), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n616), .A2(new_n618), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n619), .ZN(new_n625));
  INV_X1    g424(.A(new_n590), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n616), .A2(new_n618), .A3(new_n620), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G134gat), .B(G162gat), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n623), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n623), .B2(new_n628), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n601), .A2(new_n636), .A3(new_n600), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n595), .A2(new_n599), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n595), .B2(new_n599), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n558), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n611), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT100), .B1(new_n564), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n558), .A2(new_n644), .A3(new_n611), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n635), .B(new_n641), .C1(new_n643), .C2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n558), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n651), .B(new_n652), .C1(new_n646), .C2(new_n647), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n558), .A2(new_n640), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n564), .A2(KEYINPUT100), .A3(new_n642), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n644), .B1(new_n558), .B2(new_n611), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n658), .A2(new_n649), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n654), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n659), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n588), .A2(new_n634), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n534), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n478), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(G1gat), .Z(G1324gat));
  OAI21_X1  g471(.A(G8gat), .B1(new_n670), .B2(new_n470), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT16), .B(G8gat), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n670), .A2(new_n470), .A3(new_n675), .ZN(new_n676));
  MUX2_X1   g475(.A(new_n674), .B(KEYINPUT42), .S(new_n676), .Z(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n670), .B2(new_n522), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n515), .A2(G15gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n670), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n670), .A2(new_n441), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NOR3_X1   g482(.A1(new_n587), .A2(new_n633), .A3(new_n668), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n534), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(G29gat), .A3(new_n478), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT104), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n686), .B(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT106), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n621), .A2(new_n622), .A3(new_n590), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n626), .B1(new_n625), .B2(new_n627), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n629), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n623), .A2(new_n628), .A3(new_n630), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n519), .A2(new_n522), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n458), .A2(new_n470), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n416), .A2(new_n441), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n470), .A2(new_n530), .ZN(new_n703));
  INV_X1    g502(.A(new_n532), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n478), .A2(new_n479), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n441), .A2(new_n705), .A3(new_n526), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n703), .A2(new_n704), .B1(new_n706), .B2(KEYINPUT35), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n698), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n633), .B1(new_n524), .B2(new_n533), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n664), .A2(new_n667), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n587), .A2(KEYINPUT105), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n584), .A2(new_n586), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AND4_X1   g515(.A1(new_n263), .A2(new_n711), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n332), .B1(new_n338), .B2(new_n409), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n210), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n689), .A2(new_n719), .ZN(G1328gat));
  NOR3_X1   g519(.A1(new_n685), .A2(G36gat), .A3(new_n470), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  INV_X1    g521(.A(new_n470), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(new_n211), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n717), .A2(G43gat), .A3(new_n516), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n214), .B1(new_n685), .B2(new_n515), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT47), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n726), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1330gat));
  NAND3_X1  g531(.A1(new_n717), .A2(G50gat), .A3(new_n525), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n215), .B1(new_n685), .B2(new_n441), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT48), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1331gat));
  NOR2_X1   g538(.A1(new_n480), .A2(new_n516), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n471), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n533), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n587), .A2(new_n264), .A3(new_n633), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n712), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n478), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n539), .ZN(G1332gat));
  XOR2_X1   g546(.A(new_n745), .B(KEYINPUT107), .Z(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n723), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n750), .B2(new_n749), .ZN(G1333gat));
  NAND2_X1  g552(.A1(new_n748), .A2(new_n516), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G71gat), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n742), .A2(new_n545), .A3(new_n521), .A4(new_n744), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(KEYINPUT50), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n748), .A2(new_n525), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n588), .A2(new_n264), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n633), .B(new_n764), .C1(new_n533), .C2(new_n741), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT51), .ZN(new_n766));
  INV_X1    g565(.A(G85gat), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n718), .A4(new_n668), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n764), .A2(new_n712), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n711), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n711), .B2(new_n770), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(new_n478), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n768), .B1(new_n773), .B2(new_n767), .ZN(G1336gat));
  NOR3_X1   g573(.A1(new_n470), .A2(G92gat), .A3(new_n712), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n711), .A2(new_n770), .ZN(new_n778));
  OAI21_X1  g577(.A(G92gat), .B1(new_n778), .B2(new_n470), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n772), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n711), .A2(new_n769), .A3(new_n770), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n723), .A3(new_n782), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n783), .A2(G92gat), .B1(new_n766), .B2(new_n775), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n780), .B1(new_n784), .B2(new_n777), .ZN(G1337gat));
  INV_X1    g584(.A(G99gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n766), .A2(new_n786), .A3(new_n521), .A4(new_n668), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n771), .A2(new_n772), .A3(new_n522), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n786), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT109), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n787), .C1(new_n788), .C2(new_n786), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1338gat));
  NOR3_X1   g592(.A1(new_n441), .A2(G106gat), .A3(new_n712), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n766), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  OAI21_X1  g595(.A(G106gat), .B1(new_n778), .B2(new_n441), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n525), .A3(new_n782), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n799), .A2(G106gat), .B1(new_n766), .B2(new_n794), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n800), .B2(new_n796), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n743), .A2(new_n668), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n558), .A2(KEYINPUT10), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n615), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n658), .B2(new_n635), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n651), .B1(new_n805), .B2(new_n652), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n805), .B2(new_n652), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n648), .A2(KEYINPUT102), .A3(new_n649), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n805), .A2(new_n652), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n663), .B1(new_n811), .B2(new_n807), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n812), .A3(KEYINPUT55), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n664), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n662), .B1(new_n665), .B2(KEYINPUT54), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n654), .B2(new_n808), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT110), .B1(new_n816), .B2(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n810), .A2(new_n812), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n814), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT106), .B1(new_n631), .B2(new_n632), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n694), .A2(new_n691), .A3(new_n695), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n244), .B1(new_n243), .B2(new_n245), .ZN(new_n826));
  OAI22_X1  g625(.A1(new_n826), .A2(KEYINPUT111), .B1(new_n250), .B2(new_n251), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(KEYINPUT111), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n258), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n262), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n822), .A2(new_n825), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n712), .A2(new_n830), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n822), .B2(new_n263), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n834), .B2(new_n825), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n802), .B1(new_n835), .B2(new_n716), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT112), .B1(new_n836), .B2(new_n525), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n813), .A2(new_n664), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n819), .B1(new_n818), .B2(new_n820), .ZN(new_n839));
  AOI211_X1 g638(.A(KEYINPUT110), .B(KEYINPUT55), .C1(new_n810), .C2(new_n812), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n838), .B(new_n263), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n831), .A2(new_n668), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n825), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n838), .B(new_n831), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n697), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n716), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n743), .A2(new_n668), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n441), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n837), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n723), .A2(new_n478), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n521), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n264), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n836), .A2(new_n478), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n525), .A2(new_n527), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n856), .B1(new_n855), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n470), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n263), .A2(new_n278), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(G1340gat));
  OAI21_X1  g661(.A(G120gat), .B1(new_n853), .B2(new_n712), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT114), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n668), .A2(new_n273), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n860), .B2(new_n865), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n853), .B2(new_n716), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n588), .A2(G127gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n860), .B2(new_n868), .ZN(G1342gat));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n723), .A2(G134gat), .A3(new_n633), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n870), .B(new_n871), .C1(new_n858), .C2(new_n859), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT115), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n858), .B2(new_n859), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n853), .B2(new_n633), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n873), .A2(KEYINPUT116), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT116), .B1(new_n873), .B2(new_n877), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1343gat));
  NAND2_X1  g679(.A1(new_n852), .A2(new_n522), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n836), .A2(KEYINPUT57), .A3(new_n441), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n818), .A2(new_n820), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT117), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n884), .A2(new_n263), .A3(new_n838), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n633), .B1(new_n885), .B2(new_n833), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n587), .B1(new_n886), .B2(new_n832), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n525), .B1(new_n887), .B2(new_n802), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n881), .B(new_n882), .C1(new_n888), .C2(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(G141gat), .A3(new_n263), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n855), .A2(new_n525), .A3(new_n522), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n470), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n264), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(G141gat), .B2(new_n894), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g695(.A(G148gat), .ZN(new_n897));
  AOI211_X1 g696(.A(KEYINPUT59), .B(new_n897), .C1(new_n889), .C2(new_n668), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n441), .A2(KEYINPUT57), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n822), .A2(new_n634), .A3(new_n831), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n587), .B1(new_n886), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n902), .B2(new_n802), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n836), .B2(new_n441), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n905), .A2(new_n712), .A3(new_n881), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n899), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n668), .A2(new_n897), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n898), .A2(new_n907), .B1(new_n893), .B2(new_n908), .ZN(G1345gat));
  INV_X1    g708(.A(new_n716), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n290), .B1(new_n889), .B2(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n893), .A2(G155gat), .A3(new_n588), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  NAND4_X1  g712(.A1(new_n892), .A2(new_n291), .A3(new_n470), .A4(new_n634), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT118), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n889), .A2(new_n825), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n291), .ZN(G1347gat));
  AND3_X1   g716(.A1(new_n848), .A2(KEYINPUT119), .A3(new_n478), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT119), .B1(new_n848), .B2(new_n478), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n857), .A2(new_n723), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT120), .Z(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(KEYINPUT121), .A3(new_n922), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n263), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n470), .A2(new_n718), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n849), .B1(new_n848), .B2(new_n441), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT112), .B(new_n525), .C1(new_n846), .C2(new_n847), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n521), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n851), .A2(new_n934), .A3(new_n521), .A4(new_n929), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n264), .A2(new_n256), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n928), .B1(new_n936), .B2(new_n937), .ZN(G1348gat));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n360), .A3(new_n668), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n936), .A2(new_n668), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n360), .B2(new_n940), .ZN(G1349gat));
  AND2_X1   g740(.A1(new_n587), .A2(new_n372), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n920), .A2(new_n922), .A3(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT123), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n933), .A2(new_n935), .A3(new_n910), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G183gat), .ZN(new_n946));
  XNOR2_X1  g745(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT125), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n944), .A2(new_n950), .A3(new_n946), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n944), .A2(new_n946), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT60), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(G1350gat));
  NAND4_X1  g753(.A1(new_n925), .A2(new_n373), .A3(new_n825), .A4(new_n926), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n933), .A2(new_n935), .A3(new_n634), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n955), .B(new_n962), .C1(new_n958), .C2(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1351gat));
  NAND2_X1  g763(.A1(new_n929), .A2(new_n522), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT127), .Z(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n904), .A3(new_n903), .ZN(new_n967));
  INV_X1    g766(.A(G197gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n967), .A2(new_n968), .A3(new_n264), .ZN(new_n969));
  AND4_X1   g768(.A1(new_n525), .A2(new_n920), .A3(new_n723), .A4(new_n522), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n263), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n971), .B2(new_n968), .ZN(G1352gat));
  OAI21_X1  g771(.A(G204gat), .B1(new_n967), .B2(new_n712), .ZN(new_n973));
  INV_X1    g772(.A(G204gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n974), .A3(new_n668), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n970), .A2(new_n347), .A3(new_n587), .ZN(new_n980));
  OR3_X1    g779(.A1(new_n905), .A2(new_n588), .A3(new_n965), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  AOI21_X1  g783(.A(G218gat), .B1(new_n970), .B2(new_n825), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n967), .A2(new_n346), .A3(new_n633), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


