//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G214), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G131), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n190), .A2(KEYINPUT87), .A3(new_n191), .A4(new_n192), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n194));
  AOI21_X1  g008(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n196), .B2(new_n191), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT87), .B1(new_n196), .B2(new_n191), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT17), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT77), .A4(G125), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(G125), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(KEYINPUT16), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n203), .A2(G146), .A3(new_n206), .A4(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n196), .A2(new_n200), .A3(new_n191), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n201), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT18), .A2(G131), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n196), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G125), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G140), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n208), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT86), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n202), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n225), .A3(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n202), .A2(new_n211), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G113), .B(G122), .ZN(new_n230));
  INV_X1    g044(.A(G104), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT90), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n229), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n201), .B2(new_n216), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n236), .B2(new_n232), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT92), .B(G475), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT88), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n222), .B2(KEYINPUT19), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT19), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n202), .A2(KEYINPUT88), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n223), .A2(new_n225), .A3(KEYINPUT19), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n211), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n213), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n199), .B1(new_n249), .B2(KEYINPUT89), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT89), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n251), .A3(new_n213), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n235), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n234), .B1(new_n253), .B2(new_n232), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n255));
  NOR2_X1   g069(.A1(G475), .A2(G902), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n255), .B1(new_n254), .B2(new_n256), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT91), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(KEYINPUT91), .A3(new_n255), .A4(new_n256), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n241), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g076(.A(KEYINPUT72), .B(G902), .Z(new_n263));
  NAND2_X1  g077(.A1(new_n189), .A2(G128), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT13), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT95), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G128), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n270), .A3(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n264), .A2(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT95), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n273), .A2(new_n189), .A3(KEYINPUT13), .A4(G128), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n266), .A2(new_n271), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G134), .ZN(new_n276));
  AND2_X1   g090(.A1(KEYINPUT64), .A2(G134), .ZN(new_n277));
  NOR2_X1   g091(.A1(KEYINPUT64), .A2(G134), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n271), .A2(KEYINPUT96), .A3(new_n279), .A4(new_n264), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n271), .A2(new_n279), .A3(new_n264), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT96), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n276), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G107), .ZN(new_n285));
  INV_X1    g099(.A(G116), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G122), .ZN(new_n287));
  INV_X1    g101(.A(G122), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G116), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT93), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n287), .B2(new_n289), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n289), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT93), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(G107), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT94), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n297), .A3(KEYINPUT94), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n284), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  INV_X1    g117(.A(G217), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(new_n304), .A3(G953), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n286), .A2(KEYINPUT14), .A3(G122), .ZN(new_n307));
  OAI211_X1 g121(.A(G107), .B(new_n307), .C1(new_n294), .C2(KEYINPUT14), .ZN(new_n308));
  INV_X1    g122(.A(new_n281), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n279), .B1(new_n271), .B2(new_n264), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n293), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n302), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n275), .A2(G134), .B1(new_n281), .B2(new_n282), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n293), .A2(new_n297), .A3(KEYINPUT94), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT94), .B1(new_n293), .B2(new_n297), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n280), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n305), .B1(new_n317), .B2(new_n311), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n263), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G478), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(KEYINPUT15), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n319), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n262), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(G953), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G952), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(G234), .B2(G237), .ZN(new_n328));
  AOI211_X1 g142(.A(new_n326), .B(new_n263), .C1(G234), .C2(G237), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT21), .B(G898), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT6), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n286), .A2(G119), .ZN(new_n334));
  INV_X1    g148(.A(G119), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT67), .B1(new_n335), .B2(G116), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n286), .A3(G119), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n334), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n334), .ZN(new_n342));
  OAI21_X1  g156(.A(G113), .B1(new_n342), .B2(KEYINPUT5), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT3), .B1(new_n231), .B2(G107), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n285), .A3(G104), .ZN(new_n347));
  INV_X1    g161(.A(G101), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n231), .A2(G107), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n345), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n231), .A2(G107), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n285), .A2(G104), .ZN(new_n352));
  OAI21_X1  g166(.A(G101), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(KEYINPUT2), .A2(G113), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT66), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n358));
  INV_X1    g172(.A(G113), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n339), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n344), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n366), .A2(KEYINPUT79), .A3(G101), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT79), .B1(new_n366), .B2(G101), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(G101), .A3(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n339), .A2(new_n362), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n339), .A2(new_n362), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT81), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n366), .A2(G101), .A3(new_n371), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n339), .A2(new_n362), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n377), .B1(new_n378), .B2(new_n363), .ZN(new_n379));
  INV_X1    g193(.A(new_n369), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n366), .A2(G101), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n366), .A2(KEYINPUT79), .A3(G101), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n379), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n365), .B1(new_n376), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G110), .B(G122), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n333), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n370), .A2(new_n375), .A3(KEYINPUT81), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n386), .B1(new_n379), .B2(new_n385), .ZN(new_n392));
  OAI22_X1  g206(.A1(new_n391), .A2(new_n392), .B1(new_n344), .B2(new_n364), .ZN(new_n393));
  INV_X1    g207(.A(new_n389), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G143), .B(G146), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n211), .A2(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT1), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n268), .A2(new_n270), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT1), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n189), .A2(G146), .ZN(new_n403));
  AND4_X1   g217(.A1(new_n402), .A2(new_n398), .A3(new_n403), .A4(G128), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n220), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n398), .A2(new_n403), .A3(KEYINPUT0), .A4(G128), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT0), .B(G128), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n397), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n326), .A2(G224), .ZN(new_n412));
  XOR2_X1   g226(.A(new_n412), .B(KEYINPUT82), .Z(new_n413));
  XNOR2_X1  g227(.A(new_n411), .B(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n393), .A2(new_n333), .A3(new_n394), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n396), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n389), .B(KEYINPUT8), .ZN(new_n417));
  INV_X1    g231(.A(new_n344), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n355), .B1(new_n418), .B2(new_n363), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n340), .A2(KEYINPUT83), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n343), .B1(new_n340), .B2(KEYINPUT83), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n364), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n417), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n412), .B1(KEYINPUT84), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(KEYINPUT84), .B2(new_n424), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n426), .B1(new_n406), .B2(new_n410), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(G224), .B2(new_n326), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n406), .A2(new_n410), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT85), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n406), .A2(new_n431), .A3(new_n410), .A4(new_n428), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n427), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n423), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n388), .A2(new_n389), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G210), .B1(G237), .B2(G902), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n416), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n437), .B1(new_n416), .B2(new_n436), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n325), .B(new_n332), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n324), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n409), .ZN(new_n442));
  OR2_X1    g256(.A1(KEYINPUT64), .A2(G134), .ZN(new_n443));
  INV_X1    g257(.A(G137), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT11), .ZN(new_n445));
  NAND2_X1  g259(.A1(KEYINPUT64), .A2(G134), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(KEYINPUT11), .A3(G134), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT11), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G137), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n447), .A2(new_n191), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n448), .A2(new_n450), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n191), .B1(new_n453), .B2(new_n447), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n442), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n373), .A2(new_n374), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n191), .B1(G134), .B2(G137), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n443), .A2(new_n446), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(G137), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n451), .B(new_n459), .C1(new_n401), .C2(new_n404), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT27), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n187), .A2(new_n462), .A3(G210), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n187), .B2(G210), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT26), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n465), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT26), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n463), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n466), .A2(new_n469), .A3(G101), .ZN(new_n470));
  AOI21_X1  g284(.A(G101), .B1(new_n466), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n461), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT30), .ZN(new_n475));
  INV_X1    g289(.A(new_n460), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n449), .A2(G137), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n477), .A2(new_n277), .A3(new_n278), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n448), .A2(new_n450), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n409), .B1(new_n480), .B2(new_n451), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n475), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n378), .A2(new_n363), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n455), .A2(KEYINPUT30), .A3(new_n460), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT68), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n461), .A2(new_n472), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n474), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT31), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n476), .A2(new_n481), .A3(new_n483), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n456), .B1(new_n455), .B2(new_n460), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT28), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n461), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n472), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n474), .A2(new_n485), .A3(new_n498), .A4(new_n487), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(G472), .A2(G902), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT69), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(KEYINPUT69), .A3(new_n501), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n501), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n485), .A2(new_n461), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n496), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n480), .A2(new_n451), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n398), .A2(new_n403), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT65), .B(G128), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n402), .B1(G143), .B2(new_n211), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n397), .A2(new_n402), .A3(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n279), .A2(new_n444), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n457), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n442), .A2(new_n513), .B1(new_n520), .B2(new_n451), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT28), .B1(new_n521), .B2(new_n456), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n483), .B1(new_n476), .B2(new_n481), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n461), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n524), .B2(KEYINPUT28), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT29), .B1(new_n525), .B2(new_n472), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n509), .A2(KEYINPUT70), .A3(new_n496), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n512), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n492), .A2(KEYINPUT29), .A3(new_n494), .A4(new_n472), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT71), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT71), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n525), .A2(new_n531), .A3(KEYINPUT29), .A4(new_n472), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(new_n263), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n534), .A2(KEYINPUT73), .A3(G472), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT73), .B1(new_n534), .B2(G472), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n507), .B(new_n508), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n515), .A2(G119), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n335), .A2(G128), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT74), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT74), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n542), .A3(new_n539), .ZN(new_n543));
  XOR2_X1   g357(.A(KEYINPUT24), .B(G110), .Z(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n515), .A2(KEYINPUT23), .A3(G119), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n539), .A2(KEYINPUT75), .A3(KEYINPUT23), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n267), .A2(G119), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT75), .B1(new_n539), .B2(KEYINPUT23), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n551), .A2(KEYINPUT76), .A3(G110), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT76), .B1(new_n551), .B2(G110), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n214), .B(new_n545), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n544), .B1(new_n541), .B2(new_n543), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n546), .B(new_n556), .C1(new_n549), .C2(new_n550), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n227), .B(new_n213), .C1(new_n555), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n326), .A2(G221), .A3(G234), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT22), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(G137), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n554), .A2(new_n559), .A3(new_n563), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n263), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n304), .B1(new_n263), .B2(G234), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT25), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n565), .A2(new_n570), .A3(new_n263), .A4(new_n566), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n565), .A2(new_n566), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n569), .A2(G902), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G469), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n397), .B1(G128), .B2(new_n399), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n355), .B1(new_n404), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n517), .B2(new_n518), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n580), .A2(new_n581), .B1(new_n355), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n513), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n385), .A2(new_n442), .A3(new_n372), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n326), .A2(G227), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G140), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT78), .B(G110), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n405), .A2(new_n354), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n580), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n592), .A2(KEYINPUT12), .A3(new_n513), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT12), .B1(new_n592), .B2(new_n513), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n586), .B(new_n590), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n583), .A2(new_n585), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n513), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n590), .B1(new_n598), .B2(new_n586), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n578), .B(new_n263), .C1(new_n596), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(G469), .A2(G902), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n602));
  INV_X1    g416(.A(new_n590), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n598), .A2(new_n586), .A3(new_n590), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(G469), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n441), .A2(new_n537), .A3(new_n577), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  NAND4_X1  g426(.A1(new_n607), .A2(new_n575), .A3(new_n572), .A4(new_n608), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n504), .A2(new_n506), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n616));
  INV_X1    g430(.A(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n500), .B2(new_n263), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n614), .A2(new_n615), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n504), .A3(new_n506), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT97), .B1(new_n621), .B2(new_n613), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n260), .A2(new_n261), .ZN(new_n624));
  INV_X1    g438(.A(new_n241), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n313), .B2(new_n318), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n306), .B1(new_n302), .B2(new_n312), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n317), .A2(new_n305), .A3(new_n311), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(KEYINPUT33), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n263), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n320), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n629), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n319), .A2(new_n320), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n627), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n635), .A2(new_n627), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n626), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n440), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n623), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND2_X1  g459(.A1(new_n257), .A2(KEYINPUT99), .ZN(new_n646));
  INV_X1    g460(.A(new_n258), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n254), .A2(new_n648), .A3(new_n255), .A4(new_n256), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n322), .A3(new_n625), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n440), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n623), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n554), .A2(new_n559), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n656), .B1(new_n554), .B2(new_n559), .ZN(new_n658));
  OAI22_X1  g472(.A1(new_n657), .A2(new_n658), .B1(KEYINPUT36), .B2(new_n564), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n560), .A2(KEYINPUT100), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n564), .A2(KEYINPUT36), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n554), .A2(new_n559), .A3(new_n656), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n574), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n572), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n608), .A3(new_n607), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n621), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n441), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n328), .B1(new_n329), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n651), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n325), .B1(new_n438), .B2(new_n439), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n667), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n535), .A2(new_n536), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n507), .A2(new_n508), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n674), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  NAND2_X1  g494(.A1(new_n416), .A2(new_n436), .ZN(new_n681));
  INV_X1    g495(.A(new_n437), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n416), .A2(new_n436), .A3(new_n437), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT101), .Z(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT38), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(KEYINPUT38), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n617), .B1(new_n524), .B2(new_n496), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n488), .A2(new_n690), .B1(G472), .B2(G902), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT102), .Z(new_n692));
  NAND3_X1  g506(.A1(new_n507), .A2(new_n508), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n507), .A2(new_n695), .A3(new_n508), .A4(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n673), .B(KEYINPUT39), .Z(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n609), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT40), .ZN(new_n701));
  INV_X1    g515(.A(new_n666), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n262), .A2(new_n323), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n325), .A2(new_n701), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n689), .A2(new_n697), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  AND3_X1   g520(.A1(new_n635), .A2(new_n627), .A3(new_n636), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n637), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n262), .A2(new_n708), .A3(new_n673), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n537), .A2(new_n676), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  AND2_X1   g525(.A1(new_n507), .A2(new_n508), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n534), .A2(G472), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT73), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n534), .A2(KEYINPUT73), .A3(G472), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n576), .B1(new_n712), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n603), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n633), .B1(new_n721), .B2(new_n595), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G469), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n608), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n718), .A2(new_n642), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n718), .A2(KEYINPUT104), .A3(new_n642), .A4(new_n726), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT41), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G113), .ZN(G15));
  NAND4_X1  g547(.A1(new_n537), .A2(new_n652), .A3(new_n577), .A4(new_n726), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  AOI211_X1 g549(.A(new_n322), .B(new_n241), .C1(new_n260), .C2(new_n261), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n723), .A2(new_n666), .A3(new_n608), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n675), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n537), .A2(new_n332), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT105), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n335), .ZN(G21));
  INV_X1    g555(.A(new_n501), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT106), .B1(new_n489), .B2(new_n497), .ZN(new_n743));
  INV_X1    g557(.A(new_n499), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n489), .A2(new_n497), .A3(KEYINPUT106), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n722), .A2(new_n578), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n332), .A3(new_n608), .A4(new_n600), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n747), .A2(new_n749), .A3(new_n576), .A4(new_n618), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n675), .A2(new_n262), .A3(new_n323), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NOR2_X1   g567(.A1(new_n747), .A2(new_n618), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n738), .A2(new_n709), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  NOR3_X1   g570(.A1(new_n641), .A2(KEYINPUT42), .A3(new_n673), .ZN(new_n757));
  INV_X1    g571(.A(new_n325), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n685), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n718), .A2(new_n757), .A3(new_n610), .A4(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n508), .A2(KEYINPUT107), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n502), .A2(new_n505), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n508), .A2(KEYINPUT107), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n577), .B1(new_n677), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n709), .A2(new_n610), .A3(new_n759), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT42), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT108), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND4_X1  g584(.A1(new_n718), .A2(new_n610), .A3(new_n674), .A4(new_n759), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  XNOR2_X1  g586(.A(new_n262), .B(KEYINPUT110), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n708), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(KEYINPUT111), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n626), .A2(KEYINPUT110), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n262), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n779), .A3(new_n775), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n708), .B(KEYINPUT109), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT43), .B1(new_n784), .B2(new_n262), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n702), .B1(new_n615), .B2(new_n619), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(KEYINPUT112), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n604), .A2(new_n605), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n604), .A2(KEYINPUT45), .A3(new_n605), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(G469), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n601), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT46), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n600), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n608), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n699), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n791), .A2(new_n759), .A3(new_n792), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT112), .B1(new_n789), .B2(new_n790), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  NAND2_X1  g622(.A1(new_n803), .A2(KEYINPUT47), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n810), .B(new_n608), .C1(new_n801), .C2(new_n802), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n759), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n537), .A2(new_n814), .A3(new_n577), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(new_n709), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n819));
  INV_X1    g633(.A(new_n765), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n759), .A2(new_n726), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n787), .A2(new_n328), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT48), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n785), .B1(new_n776), .B2(new_n782), .ZN(new_n825));
  INV_X1    g639(.A(new_n328), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT48), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n820), .A4(new_n822), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n577), .A2(new_n328), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n697), .A2(new_n821), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n626), .A3(new_n640), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n327), .B(KEYINPUT118), .Z(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n726), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n754), .A2(new_n577), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n825), .A2(new_n826), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n758), .B1(new_n683), .B2(new_n684), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n830), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n830), .B2(new_n840), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT50), .ZN(new_n844));
  INV_X1    g658(.A(new_n837), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n787), .A2(new_n328), .A3(new_n726), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n687), .A2(new_n758), .A3(new_n688), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n847), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n838), .A2(KEYINPUT50), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n825), .A2(new_n826), .A3(new_n837), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n723), .A2(new_n725), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n814), .B1(new_n812), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n626), .A2(new_n640), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n852), .A2(new_n854), .B1(new_n832), .B2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n747), .A2(new_n702), .A3(new_n618), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n827), .A2(KEYINPUT117), .A3(new_n822), .A4(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n787), .A2(new_n328), .A3(new_n822), .A4(new_n857), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n856), .A2(KEYINPUT51), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n842), .A2(new_n843), .B1(new_n851), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n856), .A2(new_n858), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n848), .A2(new_n850), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n865), .B1(KEYINPUT116), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n851), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n863), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n679), .A2(new_n873), .A3(new_n755), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n679), .B2(new_n755), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n609), .A2(new_n666), .A3(new_n673), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n697), .A2(new_n751), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(KEYINPUT52), .A3(new_n710), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n872), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n703), .A3(new_n839), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n694), .B2(new_n696), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n537), .A2(new_n676), .A3(new_n709), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n885), .B(KEYINPUT115), .C1(new_n874), .C2(new_n875), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n882), .A2(new_n883), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n679), .A2(new_n755), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n884), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n880), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n262), .A2(new_n640), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n736), .ZN(new_n893));
  INV_X1    g707(.A(new_n440), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n620), .A3(new_n894), .A4(new_n622), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n669), .A3(new_n739), .A4(new_n752), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n611), .A2(new_n734), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n760), .A2(new_n771), .A3(new_n767), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n709), .A2(new_n754), .ZN(new_n900));
  INV_X1    g714(.A(new_n673), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n650), .A2(new_n625), .A3(new_n323), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT113), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n537), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n902), .A2(KEYINPUT113), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n906), .A2(new_n610), .A3(new_n666), .A4(new_n759), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n731), .A2(new_n898), .A3(new_n899), .A4(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT53), .B1(new_n891), .B2(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n887), .A2(KEYINPUT52), .A3(new_n888), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT52), .B1(new_n887), .B2(new_n888), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n898), .A2(new_n899), .A3(new_n731), .A4(new_n907), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT53), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT54), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n891), .A2(new_n908), .A3(KEYINPUT53), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(G952), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n871), .A2(new_n922), .B1(new_n923), .B2(new_n326), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n723), .B(KEYINPUT49), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n576), .A2(new_n758), .A3(new_n725), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n640), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n773), .ZN(new_n928));
  NOR4_X1   g742(.A1(new_n689), .A2(new_n927), .A3(new_n697), .A4(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n819), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n923), .A2(new_n326), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n870), .A2(new_n864), .ZN(new_n932));
  INV_X1    g746(.A(new_n863), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n934), .B2(new_n921), .ZN(new_n935));
  INV_X1    g749(.A(new_n929), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(KEYINPUT120), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n930), .A2(new_n937), .ZN(G75));
  NOR2_X1   g752(.A1(new_n326), .A2(G952), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n263), .B1(new_n917), .B2(new_n919), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT56), .B1(new_n941), .B2(new_n682), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n396), .A2(new_n415), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n414), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT55), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n940), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n941), .A2(KEYINPUT121), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n941), .A2(KEYINPUT121), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n682), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT56), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n946), .B1(new_n950), .B2(new_n952), .ZN(G51));
  INV_X1    g767(.A(new_n797), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n917), .A2(new_n919), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT54), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n920), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n601), .B(KEYINPUT57), .ZN(new_n960));
  OAI22_X1  g774(.A1(new_n959), .A2(new_n960), .B1(new_n599), .B2(new_n596), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n939), .B1(new_n955), .B2(new_n961), .ZN(G54));
  AND2_X1   g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n949), .A2(new_n254), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n947), .B2(new_n948), .ZN(new_n965));
  INV_X1    g779(.A(new_n254), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n939), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n964), .A2(new_n967), .ZN(G60));
  INV_X1    g782(.A(KEYINPUT122), .ZN(new_n969));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT59), .Z(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n916), .B2(new_n920), .ZN(new_n972));
  INV_X1    g786(.A(new_n629), .ZN(new_n973));
  INV_X1    g787(.A(new_n632), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n969), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n975), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n977), .A2(new_n971), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n939), .B1(new_n958), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n972), .A2(new_n969), .A3(new_n975), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT123), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(KEYINPUT122), .B(new_n977), .C1(new_n922), .C2(new_n971), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT123), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n983), .A2(new_n984), .A3(new_n976), .A4(new_n979), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n985), .ZN(G63));
  XNOR2_X1  g800(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n304), .A2(new_n238), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n987), .B(new_n988), .Z(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n917), .B2(new_n919), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n940), .B1(new_n990), .B2(new_n573), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n664), .B2(new_n990), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g807(.A(G224), .ZN(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n330), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n898), .A2(new_n731), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT125), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n997), .A2(KEYINPUT126), .A3(new_n326), .ZN(new_n998));
  AOI21_X1  g812(.A(KEYINPUT126), .B1(new_n997), .B2(new_n326), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n943), .B1(G898), .B2(new_n326), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(G69));
  NAND2_X1  g816(.A1(new_n482), .A2(new_n484), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n246), .A2(new_n247), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G900), .A2(G953), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n876), .A2(new_n883), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n804), .A2(new_n751), .A3(new_n820), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n817), .A2(new_n899), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n807), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n1005), .B(new_n1006), .C1(new_n1010), .C2(G953), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1007), .A2(new_n705), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n718), .A2(new_n610), .A3(new_n759), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n892), .A2(new_n736), .A3(new_n699), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n817), .A2(new_n1013), .A3(new_n1014), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(G953), .B1(new_n1019), .B2(new_n807), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1011), .B1(new_n1020), .B2(new_n1005), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n326), .B1(G227), .B2(G900), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(G72));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n1019), .A2(new_n807), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n1026), .B2(new_n997), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1027), .A2(new_n472), .A3(new_n509), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1025), .B1(new_n1010), .B2(new_n997), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1029), .A2(new_n461), .A3(new_n496), .A4(new_n485), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n909), .A2(new_n915), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1025), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n512), .A2(new_n527), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1032), .B1(new_n1033), .B2(new_n488), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT127), .Z(new_n1035));
  AOI21_X1  g849(.A(new_n939), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  AND3_X1   g850(.A1(new_n1028), .A2(new_n1030), .A3(new_n1036), .ZN(G57));
endmodule


