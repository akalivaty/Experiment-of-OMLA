//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n211), .B(new_n217), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n225), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n205), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT64), .ZN(new_n242));
  INV_X1    g0042(.A(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G222), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G223), .A2(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n257), .B(new_n260), .C1(G77), .C2(new_n253), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n269), .A2(new_n259), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT65), .B(G226), .Z(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  INV_X1    g0073(.A(new_n214), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n258), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n261), .A2(new_n272), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G200), .ZN(new_n279));
  INV_X1    g0079(.A(G190), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT67), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT67), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n285), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n214), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G150), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n215), .A2(G33), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n201), .A2(new_n215), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n287), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT66), .B(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(G50), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n266), .A2(new_n268), .A3(G13), .A4(G20), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G50), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n294), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT70), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n289), .B1(new_n201), .B2(new_n215), .C1(new_n290), .C2(new_n291), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n300), .B1(new_n304), .B2(new_n287), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(new_n298), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n303), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n308), .B1(new_n303), .B2(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n282), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT72), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT10), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n302), .A2(KEYINPUT70), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n306), .B1(new_n305), .B2(new_n298), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT9), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n281), .B1(new_n317), .B2(new_n309), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT72), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n282), .B(new_n319), .C1(new_n310), .C2(new_n311), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(KEYINPUT71), .A3(new_n319), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n278), .A2(G179), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT68), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(KEYINPUT68), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n278), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n333), .A4(new_n302), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT76), .ZN(new_n335));
  INV_X1    g0135(.A(G226), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n254), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n225), .A2(G1698), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n260), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n269), .A2(G238), .A3(new_n259), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .A4(new_n277), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n277), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n259), .B1(new_n341), .B2(new_n342), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT13), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT73), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(KEYINPUT73), .B(KEYINPUT13), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(G169), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(KEYINPUT75), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n356), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n352), .A2(G169), .A3(new_n353), .A4(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n347), .A2(new_n350), .A3(G179), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n299), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(KEYINPUT12), .A3(new_n226), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n226), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n202), .B2(new_n291), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(KEYINPUT11), .A3(new_n287), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n363), .B(new_n366), .C1(KEYINPUT12), .C2(new_n362), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n295), .A2(new_n297), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n226), .B1(new_n368), .B2(KEYINPUT12), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT11), .B1(new_n365), .B2(new_n287), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n361), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n352), .A2(G200), .A3(new_n353), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT74), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n352), .A2(new_n376), .A3(G200), .A4(new_n353), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n347), .A2(new_n350), .A3(G190), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n373), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n327), .B(new_n334), .C1(new_n335), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n335), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n295), .A2(G77), .A3(new_n297), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n362), .A2(new_n202), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G20), .A2(G77), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT15), .B(G87), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n291), .ZN(new_n390));
  INV_X1    g0190(.A(new_n290), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n288), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n386), .B(new_n387), .C1(new_n392), .C2(new_n295), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT69), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n394), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G238), .A2(G1698), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n253), .B(new_n398), .C1(new_n225), .C2(G1698), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n260), .C1(G107), .C2(new_n253), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n270), .A2(G244), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n277), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(G179), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n332), .B2(new_n402), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n402), .A2(new_n280), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(G200), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n395), .A2(new_n396), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n362), .A2(new_n290), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n368), .B2(new_n290), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n251), .A2(new_n215), .A3(new_n252), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n252), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n226), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n224), .A2(new_n226), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G58), .A2(G68), .ZN(new_n420));
  OAI21_X1  g0220(.A(G20), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n288), .A2(G159), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n413), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n287), .ZN(new_n425));
  NOR4_X1   g0225(.A1(new_n339), .A2(new_n340), .A3(new_n415), .A4(G20), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT77), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n226), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n416), .A2(KEYINPUT77), .A3(new_n417), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n413), .B(new_n423), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n412), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n269), .A2(G232), .A3(new_n259), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n269), .A2(KEYINPUT78), .A3(G232), .A4(new_n259), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n276), .A2(new_n259), .A3(G274), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n336), .A2(G1698), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(G223), .B2(G1698), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n339), .A2(new_n340), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n439), .A2(new_n440), .B1(new_n250), .B2(new_n220), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n437), .B1(new_n441), .B2(new_n260), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n436), .A2(new_n280), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(G200), .B1(new_n436), .B2(new_n442), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT17), .B1(new_n431), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT7), .B1(new_n440), .B2(new_n215), .ZN(new_n447));
  OAI21_X1  g0247(.A(G68), .B1(new_n447), .B2(new_n426), .ZN(new_n448));
  INV_X1    g0248(.A(new_n423), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n295), .B1(new_n450), .B2(new_n413), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT16), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n411), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT17), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n436), .A2(new_n442), .ZN(new_n456));
  INV_X1    g0256(.A(G200), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n436), .A2(new_n280), .A3(new_n442), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n454), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n446), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n436), .A2(G179), .A3(new_n442), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n332), .B1(new_n436), .B2(new_n442), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n454), .A2(new_n465), .A3(KEYINPUT18), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT18), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n456), .A2(G169), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n436), .A2(G179), .A3(new_n442), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n467), .B1(new_n431), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n385), .A2(new_n409), .A3(new_n462), .A4(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n384), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n219), .A2(G1698), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(G238), .B2(G1698), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n478), .B2(new_n440), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n260), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n266), .A2(new_n268), .A3(G45), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n221), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n266), .A2(new_n268), .A3(G45), .A4(new_n273), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n259), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n475), .B1(new_n485), .B2(new_n280), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n480), .A2(new_n484), .A3(KEYINPUT87), .A4(G190), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n220), .A2(new_n204), .A3(new_n205), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n342), .A2(new_n215), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT19), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n215), .B(G68), .C1(new_n339), .C2(new_n340), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n291), .A2(new_n204), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n491), .B(new_n492), .C1(KEYINPUT19), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n287), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n362), .A2(new_n389), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n266), .A2(new_n268), .A3(G33), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n295), .A2(G87), .A3(new_n299), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n457), .B1(new_n480), .B2(new_n484), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G179), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n480), .A2(new_n484), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(G169), .B1(new_n480), .B2(new_n484), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n283), .A2(KEYINPUT67), .B1(G1), .B2(G13), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n299), .A2(new_n497), .A3(new_n506), .A4(new_n286), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n495), .B(new_n496), .C1(new_n389), .C2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n488), .A2(new_n501), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(G250), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n440), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n514), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n253), .A2(new_n516), .A3(KEYINPUT82), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n512), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n219), .A2(G1698), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n339), .B2(new_n340), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n519), .B(KEYINPUT81), .C1(new_n340), .C2(new_n339), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n259), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT85), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT5), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n263), .B1(new_n528), .B2(G41), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n296), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G257), .A3(new_n259), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT83), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n528), .B2(G41), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n262), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(new_n296), .A3(new_n275), .A4(new_n529), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n526), .A2(new_n527), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n515), .A2(new_n517), .ZN(new_n540));
  INV_X1    g0340(.A(new_n512), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n525), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n260), .ZN(new_n543));
  INV_X1    g0343(.A(new_n538), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT85), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(G190), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n532), .A2(new_n537), .A3(KEYINPUT84), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT84), .B1(new_n532), .B2(new_n537), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n543), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n288), .A2(G77), .ZN(new_n553));
  XNOR2_X1  g0353(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n206), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT79), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n557), .A2(KEYINPUT6), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(KEYINPUT6), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(new_n204), .B2(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n556), .A2(new_n560), .A3(G20), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n205), .B1(new_n416), .B2(new_n417), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n553), .B(new_n561), .C1(new_n562), .C2(KEYINPUT80), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(KEYINPUT80), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n287), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n299), .A2(G97), .ZN(new_n566));
  INV_X1    g0366(.A(new_n507), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n546), .A2(new_n552), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT86), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n527), .B1(new_n526), .B2(new_n538), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n543), .A2(KEYINPUT85), .A3(new_n544), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(new_n332), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n548), .A2(new_n543), .A3(new_n550), .A4(new_n502), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n572), .B1(new_n571), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n509), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n531), .A2(G264), .A3(new_n259), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G294), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G257), .A2(G1698), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n440), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT90), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n253), .A2(new_n585), .A3(G250), .A4(new_n254), .ZN(new_n586));
  OAI211_X1 g0386(.A(G250), .B(new_n254), .C1(new_n339), .C2(new_n340), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT90), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n537), .B(new_n581), .C1(new_n589), .C2(new_n259), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n332), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n588), .A2(new_n586), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n260), .B1(new_n592), .B2(new_n584), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n593), .A2(new_n502), .A3(new_n537), .A4(new_n581), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n215), .B(G87), .C1(new_n339), .C2(new_n340), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT22), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT22), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n253), .A2(new_n598), .A3(new_n215), .A4(G87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n476), .A2(G20), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n215), .B2(G107), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n595), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n600), .A2(new_n595), .A3(new_n605), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n295), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT25), .ZN(new_n610));
  OR4_X1    g0410(.A1(KEYINPUT89), .A2(new_n299), .A3(new_n610), .A4(G107), .ZN(new_n611));
  AOI21_X1  g0411(.A(G107), .B1(new_n610), .B2(KEYINPUT89), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n299), .A2(new_n613), .B1(KEYINPUT89), .B2(new_n610), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n611), .A2(new_n614), .B1(new_n567), .B2(G107), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n591), .B(new_n594), .C1(new_n609), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n608), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n287), .B1(new_n618), .B2(new_n606), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n593), .A2(G190), .A3(new_n537), .A4(new_n581), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n590), .A2(G200), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n615), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n531), .A2(G270), .A3(new_n259), .ZN(new_n624));
  INV_X1    g0424(.A(G303), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n251), .A2(new_n625), .A3(new_n252), .ZN(new_n626));
  MUX2_X1   g0426(.A(G257), .B(G264), .S(G1698), .Z(new_n627));
  OAI211_X1 g0427(.A(new_n260), .B(new_n626), .C1(new_n627), .C2(new_n440), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(new_n537), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G200), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n624), .A2(new_n537), .A3(G190), .A4(new_n628), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(G20), .B1(G33), .B2(G283), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n250), .A2(G97), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(new_n634), .B1(G20), .B2(new_n243), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n287), .A2(KEYINPUT20), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT20), .B1(new_n287), .B2(new_n635), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n362), .A2(new_n243), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n507), .B2(new_n243), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT88), .B1(new_n632), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n638), .A2(new_n640), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT88), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n630), .A3(new_n644), .A4(new_n631), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(G169), .B(new_n629), .C1(new_n638), .C2(new_n640), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT21), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(G179), .A2(new_n624), .A3(new_n537), .A4(new_n628), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n647), .A2(new_n648), .B1(new_n641), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n646), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n474), .A2(new_n580), .A3(new_n623), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n472), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT92), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n405), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n397), .A2(new_n404), .A3(KEYINPUT92), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n382), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n373), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n654), .B1(new_n660), .B2(new_n462), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n321), .A2(new_n326), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n334), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n384), .A2(new_n473), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n509), .A2(new_n622), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n617), .A2(new_n649), .A3(new_n651), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n571), .A2(new_n666), .A3(new_n667), .A4(new_n577), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n505), .A2(new_n508), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n509), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n577), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AND4_X1   g0473(.A1(KEYINPUT91), .A2(new_n575), .A3(new_n569), .A4(new_n576), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n526), .A2(new_n547), .A3(new_n549), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n675), .A2(new_n502), .B1(new_n565), .B2(new_n568), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT91), .B1(new_n676), .B2(new_n575), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n509), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n678), .B2(new_n672), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n665), .B1(new_n670), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n664), .A2(new_n680), .ZN(G369));
  AND2_X1   g0481(.A1(new_n215), .A2(G13), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n296), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT27), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n296), .A2(new_n685), .A3(new_n682), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G343), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT93), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n643), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n651), .A2(new_n649), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n652), .B2(new_n692), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n691), .B1(new_n619), .B2(new_n615), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n697), .A2(new_n623), .B1(new_n617), .B2(new_n691), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n690), .B1(new_n651), .B2(new_n649), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(new_n617), .A3(new_n622), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n617), .B2(new_n690), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  NAND3_X1  g0504(.A1(new_n209), .A2(KEYINPUT94), .A3(new_n262), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT94), .B1(new_n209), .B2(new_n262), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR4_X1   g0508(.A1(new_n708), .A2(new_n265), .A3(G116), .A4(new_n489), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n213), .B2(new_n708), .ZN(new_n710));
  XNOR2_X1  g0510(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n485), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G179), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n551), .A2(new_n590), .A3(new_n629), .A4(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n650), .A2(new_n593), .A3(new_n714), .A4(new_n581), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n573), .B2(new_n574), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n718), .B2(KEYINPUT30), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n720), .B(new_n717), .C1(new_n573), .C2(new_n574), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT31), .B(new_n690), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n581), .B1(new_n589), .B2(new_n259), .ZN(new_n724));
  NOR4_X1   g0524(.A1(new_n724), .A2(new_n629), .A3(new_n502), .A4(new_n485), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n545), .B2(new_n539), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n720), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(new_n716), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT31), .B1(new_n729), .B2(new_n690), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n652), .A2(new_n623), .A3(new_n690), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n509), .C1(new_n578), .C2(new_n579), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n713), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n691), .B1(new_n679), .B2(new_n670), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n575), .A2(new_n569), .A3(new_n576), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT26), .B1(new_n738), .B2(new_n509), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT91), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n577), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n676), .A2(KEYINPUT91), .A3(new_n575), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n671), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n743), .B2(KEYINPUT26), .ZN(new_n744));
  OAI211_X1 g0544(.A(KEYINPUT29), .B(new_n691), .C1(new_n744), .C2(new_n670), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n734), .B1(new_n737), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n712), .B1(new_n746), .B2(G1), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT96), .Z(G364));
  AOI21_X1  g0548(.A(new_n265), .B1(new_n682), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n708), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n696), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G330), .B2(new_n695), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n253), .A2(new_n209), .ZN(new_n754));
  INV_X1    g0554(.A(G355), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n755), .B1(G116), .B2(new_n209), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n247), .A2(G45), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n440), .A2(new_n209), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n263), .B2(new_n213), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n756), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n214), .B1(G20), .B2(new_n332), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n751), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n215), .B1(new_n768), .B2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n215), .A2(new_n457), .A3(G179), .A4(G190), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n502), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n625), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n215), .A2(new_n502), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n771), .B(new_n776), .C1(G326), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n280), .A3(G200), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n783), .B2(KEYINPUT98), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(KEYINPUT98), .B2(new_n783), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n215), .A2(new_n502), .A3(new_n280), .A4(G200), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n253), .B1(new_n786), .B2(G322), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n768), .A2(G20), .A3(new_n280), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR4_X1   g0589(.A1(new_n215), .A2(new_n502), .A3(G190), .A4(G200), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G329), .A2(new_n789), .B1(new_n790), .B2(G311), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n780), .A2(new_n785), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n790), .ZN(new_n793));
  INV_X1    g0593(.A(new_n786), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n253), .B1(new_n793), .B2(new_n202), .C1(new_n794), .C2(new_n224), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n775), .A2(new_n220), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n788), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(KEYINPUT32), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n795), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n781), .A2(new_n226), .B1(new_n769), .B2(new_n204), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT97), .ZN(new_n803));
  INV_X1    g0603(.A(G50), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n773), .A2(new_n205), .B1(new_n804), .B2(new_n778), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(KEYINPUT32), .B2(new_n799), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n801), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n792), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n767), .B1(new_n808), .B2(new_n764), .ZN(new_n809));
  INV_X1    g0609(.A(new_n763), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n695), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n753), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  NAND2_X1  g0613(.A1(new_n397), .A2(new_n690), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n405), .A2(new_n814), .A3(new_n408), .ZN(new_n815));
  INV_X1    g0615(.A(new_n814), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n658), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n735), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n815), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n656), .A2(new_n657), .A3(new_n816), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n691), .B(new_n821), .C1(new_n679), .C2(new_n670), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n731), .A2(new_n733), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G330), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT101), .Z(new_n827));
  AOI21_X1  g0627(.A(new_n751), .B1(new_n823), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n751), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n764), .A2(new_n761), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(new_n202), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n764), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n793), .A2(new_n243), .B1(new_n625), .B2(new_n778), .ZN(new_n834));
  INV_X1    g0634(.A(new_n781), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(G283), .B2(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT99), .Z(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n440), .B1(new_n838), .B2(new_n788), .C1(new_n794), .C2(new_n770), .ZN(new_n839));
  INV_X1    g0639(.A(new_n769), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(G97), .B1(new_n772), .B2(G87), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n205), .B2(new_n775), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n837), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n786), .A2(G143), .B1(new_n790), .B2(G159), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n844), .B1(new_n845), .B2(new_n778), .C1(new_n846), .C2(new_n781), .ZN(new_n847));
  XOR2_X1   g0647(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n440), .B1(new_n789), .B2(G132), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n226), .B2(new_n773), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n769), .A2(new_n224), .B1(new_n804), .B2(new_n775), .ZN(new_n853));
  NOR4_X1   g0653(.A1(new_n849), .A2(new_n850), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n843), .A2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n832), .B1(new_n833), .B2(new_n855), .C1(new_n821), .C2(new_n762), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n829), .A2(new_n856), .ZN(G384));
  NAND2_X1  g0657(.A1(new_n556), .A2(new_n560), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT35), .ZN(new_n859));
  OAI211_X1 g0659(.A(G116), .B(new_n216), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT36), .ZN(new_n862));
  OAI21_X1  g0662(.A(G77), .B1(new_n224), .B2(new_n226), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n863), .A2(new_n212), .B1(G50), .B2(new_n226), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n296), .A2(G13), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n373), .A2(new_n690), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT18), .B1(new_n454), .B2(new_n465), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n431), .A2(new_n470), .A3(new_n467), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n431), .A2(new_n445), .A3(KEYINPUT17), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n455), .B1(new_n454), .B2(new_n460), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n452), .A2(KEYINPUT16), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n295), .B1(new_n452), .B2(KEYINPUT16), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n411), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(new_n687), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n463), .A2(new_n464), .A3(new_n688), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n876), .A2(new_n878), .B1(new_n431), .B2(new_n445), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n454), .A2(new_n460), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n431), .A2(new_n470), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n431), .A2(new_n688), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n873), .A2(new_n877), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT102), .B1(new_n886), .B2(KEYINPUT38), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT102), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n880), .A2(new_n885), .ZN(new_n890));
  INV_X1    g0690(.A(new_n877), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n472), .B2(new_n462), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n886), .A2(KEYINPUT38), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n887), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT39), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n890), .A2(new_n892), .A3(new_n889), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n873), .A2(new_n431), .A3(new_n688), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n885), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n868), .B1(new_n896), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n472), .A2(new_n688), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n690), .A2(new_n372), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n373), .A2(new_n382), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n380), .B1(new_n375), .B2(new_n377), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n372), .B(new_n690), .C1(new_n910), .C2(new_n361), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n405), .A2(new_n690), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n822), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n907), .B1(new_n915), .B2(new_n895), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n906), .B1(new_n916), .B2(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n822), .A2(new_n914), .ZN(new_n918));
  INV_X1    g0718(.A(new_n912), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n895), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n907), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT103), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT105), .ZN(new_n926));
  INV_X1    g0726(.A(new_n673), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n743), .B2(KEYINPUT26), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n668), .A2(new_n669), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n690), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n745), .B1(new_n930), .B2(KEYINPUT29), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n926), .B1(new_n931), .B2(new_n474), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n737), .A2(new_n665), .A3(KEYINPUT105), .A4(new_n745), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n664), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n925), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n824), .A2(new_n821), .A3(new_n919), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n887), .A2(new_n893), .A3(new_n894), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT40), .B1(new_n897), .B2(new_n902), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n940), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n665), .A2(new_n824), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(G330), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n936), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n296), .B2(new_n682), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n936), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n866), .B1(new_n948), .B2(new_n949), .ZN(G367));
  AND2_X1   g0750(.A1(new_n571), .A2(new_n577), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n690), .A2(new_n569), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n951), .A2(new_n952), .B1(new_n738), .B2(new_n690), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n699), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n952), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n738), .A2(new_n690), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n701), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n577), .B1(new_n956), .B2(new_n617), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n960), .A2(KEYINPUT42), .B1(new_n961), .B2(new_n691), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(KEYINPUT42), .B2(new_n960), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n690), .A2(new_n499), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n671), .B(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n963), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n968), .B1(new_n963), .B2(new_n969), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n955), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n963), .A2(KEYINPUT43), .A3(new_n966), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(new_n954), .A3(new_n970), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT44), .B1(new_n958), .B2(new_n703), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n953), .A2(new_n978), .A3(new_n702), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n958), .A2(KEYINPUT45), .A3(new_n703), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT45), .B1(new_n958), .B2(new_n703), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n977), .B(new_n979), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT106), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n699), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n701), .B1(new_n698), .B2(new_n700), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n696), .B(new_n985), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n746), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n699), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n982), .A2(KEYINPUT106), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n746), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n708), .B(KEYINPUT41), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n976), .B1(new_n994), .B2(new_n749), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n794), .A2(new_n846), .B1(new_n788), .B2(new_n845), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n440), .B(new_n996), .C1(G50), .C2(new_n790), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n224), .B2(new_n775), .C1(new_n226), .C2(new_n769), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n773), .A2(new_n202), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G143), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n778), .C1(new_n797), .C2(new_n781), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n253), .B1(new_n786), .B2(G303), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n775), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT46), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n775), .B2(new_n243), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n789), .A2(G317), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(new_n1005), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n773), .A2(new_n204), .B1(new_n838), .B2(new_n778), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G294), .B2(new_n835), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n793), .A2(new_n774), .B1(new_n769), .B2(new_n205), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT108), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n998), .A2(new_n1002), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT47), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n833), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n758), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n238), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1022), .B(new_n765), .C1(new_n209), .C2(new_n389), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n751), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT107), .Z(new_n1025));
  OAI211_X1 g0825(.A(new_n1020), .B(new_n1025), .C1(new_n966), .C2(new_n810), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT109), .B1(new_n995), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n992), .B1(new_n990), .B2(new_n746), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n975), .B(new_n973), .C1(new_n1029), .C2(new_n750), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT109), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n1026), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(G387));
  NAND2_X1  g0834(.A1(new_n235), .A2(G45), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n391), .A2(new_n804), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n489), .A2(G116), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n263), .C1(new_n226), .C2(new_n202), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1035), .B(new_n1021), .C1(new_n1037), .C2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(G107), .B2(new_n209), .C1(new_n1038), .C2(new_n754), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n830), .B1(new_n1041), .B2(new_n765), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n698), .B2(new_n810), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n794), .A2(new_n804), .B1(new_n793), .B2(new_n226), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n440), .B(new_n1044), .C1(G150), .C2(new_n789), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n389), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n840), .A2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G159), .A2(new_n779), .B1(new_n835), .B2(new_n391), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n772), .A2(G97), .B1(new_n1004), .B2(G77), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n786), .A2(G317), .B1(new_n790), .B2(G303), .ZN(new_n1051));
  INV_X1    g0851(.A(G322), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1051), .B1(new_n838), .B2(new_n781), .C1(new_n1052), .C2(new_n778), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n769), .A2(new_n774), .B1(new_n770), .B2(new_n775), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT110), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT111), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT49), .Z(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT112), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n253), .B1(new_n789), .B2(G326), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n243), .C2(new_n773), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1061), .A2(KEYINPUT112), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1050), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1043), .B1(new_n1066), .B2(new_n764), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n750), .B2(new_n986), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n746), .A2(new_n986), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n708), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n746), .A2(new_n986), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(G393));
  XNOR2_X1  g0872(.A(new_n982), .B(new_n988), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1073), .A2(new_n749), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n953), .A2(new_n763), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n244), .A2(new_n1021), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n765), .C1(new_n204), .C2(new_n209), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(KEYINPUT113), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n751), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n779), .A2(G317), .B1(new_n786), .B2(G311), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n440), .B1(new_n1052), .B2(new_n788), .C1(new_n793), .C2(new_n770), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n773), .A2(new_n205), .B1(new_n775), .B2(new_n774), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n781), .A2(new_n625), .B1(new_n769), .B2(new_n243), .ZN(new_n1086));
  NOR4_X1   g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT115), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n769), .A2(new_n202), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n773), .A2(new_n220), .B1(new_n804), .B2(new_n781), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(G68), .C2(new_n1004), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n794), .A2(new_n797), .B1(new_n778), .B2(new_n846), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n253), .B1(new_n1001), .B2(new_n788), .C1(new_n793), .C2(new_n290), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1088), .A2(KEYINPUT115), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1089), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1078), .B(new_n1080), .C1(new_n764), .C2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1074), .B1(new_n1075), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1073), .A2(new_n1069), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n708), .A3(new_n990), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1101), .B1(new_n1104), .B2(new_n1105), .ZN(G390));
  INV_X1    g0906(.A(new_n708), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n474), .A2(new_n825), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n663), .B(new_n1108), .C1(new_n932), .C2(new_n933), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n733), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n729), .A2(new_n690), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT31), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n722), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n821), .C1(new_n1110), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n912), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n734), .A2(new_n821), .A3(new_n919), .ZN(new_n1117));
  OAI211_X1 g0917(.A(KEYINPUT26), .B(new_n509), .C1(new_n674), .C2(new_n677), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n672), .B1(new_n577), .B2(new_n671), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n690), .B1(new_n929), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n913), .B1(new_n1121), .B2(new_n821), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1116), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n918), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT117), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AND4_X1   g0927(.A1(G330), .A2(new_n824), .A3(new_n821), .A4(new_n919), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n919), .B1(new_n734), .B2(new_n821), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1126), .B(new_n918), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1109), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n903), .A2(new_n867), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1122), .B2(new_n912), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n867), .B1(new_n918), .B2(new_n919), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n896), .A2(new_n905), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1128), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1134), .B(new_n1117), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1107), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n918), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT117), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n1130), .A3(new_n1123), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(new_n1138), .A3(new_n1139), .A4(new_n1109), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1138), .A2(new_n750), .A3(new_n1139), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT118), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n896), .A2(new_n905), .A3(new_n761), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n831), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1150), .A2(new_n391), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n440), .B1(new_n793), .B2(new_n204), .C1(new_n794), .C2(new_n243), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n781), .A2(new_n205), .B1(new_n778), .B2(new_n774), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n796), .A4(new_n1090), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n773), .A2(new_n226), .B1(new_n770), .B2(new_n788), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT120), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n253), .B1(new_n1158), .B2(new_n788), .C1(new_n773), .C2(new_n804), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT119), .Z(new_n1160));
  NOR2_X1   g0960(.A1(new_n775), .A2(new_n846), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n835), .A2(G137), .B1(new_n840), .B2(G159), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n779), .A2(G128), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G132), .A2(new_n786), .B1(new_n1166), .B2(new_n790), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1155), .A2(new_n1157), .B1(new_n1160), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n830), .B(new_n1151), .C1(new_n1169), .C2(new_n764), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1149), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1146), .A2(new_n1148), .A3(new_n1171), .ZN(G378));
  INV_X1    g0972(.A(KEYINPUT122), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n817), .B(new_n912), .C1(new_n731), .C2(new_n733), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT40), .B1(new_n1174), .B2(new_n895), .ZN(new_n1175));
  OAI21_X1  g0975(.A(G330), .B1(new_n938), .B2(new_n941), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n941), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n713), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n940), .A3(KEYINPUT122), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n334), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n662), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1181), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n327), .A2(new_n334), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n687), .B1(new_n303), .B2(new_n307), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1177), .A2(new_n1180), .A3(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1188), .A2(KEYINPUT122), .A3(new_n940), .A4(new_n1179), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1190), .A2(new_n925), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n925), .B1(new_n1191), .B2(new_n1190), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n750), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(new_n761), .ZN(new_n1195));
  INV_X1    g0995(.A(G128), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n794), .A2(new_n1196), .B1(new_n793), .B2(new_n845), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n835), .A2(G132), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n1158), .B2(new_n778), .C1(new_n775), .C2(new_n1165), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(G150), .C2(new_n840), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT59), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n789), .A2(G124), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G33), .A2(G41), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n773), .C2(new_n797), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT121), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1202), .A2(new_n1203), .A3(new_n1207), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G50), .B(new_n1205), .C1(new_n440), .C2(new_n262), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n773), .A2(new_n224), .B1(new_n243), .B2(new_n778), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G97), .B2(new_n835), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G41), .B(new_n253), .C1(new_n789), .C2(G283), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G107), .A2(new_n786), .B1(new_n1046), .B2(new_n790), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n840), .A2(G68), .B1(G77), .B2(new_n1004), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1209), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1208), .B(new_n1217), .C1(new_n1216), .C2(new_n1215), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n764), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n831), .A2(new_n804), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1195), .A2(new_n751), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1194), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1109), .B1(new_n1223), .B2(new_n1140), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1107), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n925), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1190), .A2(new_n925), .A3(new_n1191), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(KEYINPUT123), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1226), .B1(new_n1145), .B2(new_n1109), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT123), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1193), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1222), .B1(new_n1227), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(G375));
  OAI211_X1 g1038(.A(new_n934), .B(new_n664), .C1(new_n474), .C2(new_n825), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1142), .A2(KEYINPUT117), .B1(new_n1240), .B2(new_n1122), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1130), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n993), .A3(new_n1132), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n912), .A2(new_n761), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n751), .B1(G68), .B2(new_n1150), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n794), .A2(new_n774), .B1(new_n793), .B2(new_n205), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n253), .B(new_n1246), .C1(G303), .C2(new_n789), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n781), .A2(new_n243), .B1(new_n204), .B2(new_n775), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G294), .B2(new_n779), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1247), .A2(new_n1000), .A3(new_n1047), .A4(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n840), .A2(G50), .B1(new_n790), .B2(G150), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT124), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G132), .A2(new_n779), .B1(new_n835), .B2(new_n1166), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n253), .B1(new_n788), .B2(new_n1196), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G137), .B2(new_n786), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n772), .A2(G58), .B1(new_n1004), .B2(G159), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1250), .B1(new_n1252), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1245), .B1(new_n1258), .B2(new_n764), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1144), .A2(new_n750), .B1(new_n1244), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1243), .A2(new_n1260), .ZN(G381));
  INV_X1    g1061(.A(G378), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G390), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1237), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT125), .ZN(G407));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1237), .A2(new_n1262), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(G407), .A2(G213), .A3(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(new_n1268), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n708), .B(new_n1132), .C1(new_n1242), .C2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT60), .B1(new_n1223), .B2(new_n1239), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1260), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G384), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1242), .A2(new_n1272), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1223), .A2(KEYINPUT60), .A3(new_n1239), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n708), .A4(new_n1132), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(G384), .A3(new_n1260), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1171), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1285));
  AOI221_X4 g1085(.A(new_n1222), .B1(new_n1148), .B2(new_n1285), .C1(new_n1227), .C2(new_n1236), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1221), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1230), .A2(new_n1231), .B1(new_n1145), .B2(new_n1109), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(new_n993), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1232), .A2(new_n750), .A3(new_n1235), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G378), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1271), .B(new_n1283), .C1(new_n1286), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1222), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n708), .B1(new_n1288), .B2(KEYINPUT57), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G378), .B(new_n1295), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1221), .B1(new_n1225), .B2(new_n992), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1232), .A2(new_n750), .A3(new_n1235), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1262), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1268), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1283), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1268), .A2(G2897), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1277), .A2(new_n1281), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1291), .B1(G378), .B2(new_n1237), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1309), .B2(new_n1268), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1293), .A2(new_n1294), .A3(new_n1304), .A4(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(new_n812), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1030), .A2(new_n1026), .ZN(new_n1314));
  AND2_X1   g1114(.A1(G390), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1263), .B2(new_n1315), .ZN(new_n1316));
  OR2_X1    g1116(.A1(G390), .A2(new_n1314), .ZN(new_n1317));
  OAI21_X1  g1117(.A(G390), .B1(new_n995), .B2(new_n1027), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(new_n1312), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1311), .A2(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1280), .A2(G384), .A3(new_n1260), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G384), .B1(new_n1280), .B2(new_n1260), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G2897), .B(new_n1268), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1277), .A2(new_n1281), .A3(new_n1305), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1320), .B(new_n1294), .C1(new_n1302), .C2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  AOI211_X1 g1129(.A(new_n1268), .B(new_n1282), .C1(new_n1298), .C2(new_n1301), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT126), .B1(new_n1330), .B2(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(KEYINPUT63), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1292), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1329), .A2(new_n1331), .A3(new_n1332), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1322), .A2(new_n1336), .ZN(G405));
  NOR2_X1   g1137(.A1(new_n1283), .A2(KEYINPUT127), .ZN(new_n1338));
  AND2_X1   g1138(.A1(new_n1320), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT127), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1298), .B1(new_n1340), .B2(new_n1282), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1237), .A2(G378), .ZN(new_n1342));
  OR2_X1    g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1320), .A2(new_n1338), .ZN(new_n1344));
  OR3_X1    g1144(.A1(new_n1339), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1343), .B1(new_n1339), .B2(new_n1344), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(G402));
endmodule


