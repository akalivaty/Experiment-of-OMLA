//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139, new_n1140, new_n1141;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n464), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n467), .A2(KEYINPUT68), .A3(G137), .A4(new_n463), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n463), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  MUX2_X1   g058(.A(G100), .B(G112), .S(G2105), .Z(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(G114), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G102), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n467), .A2(new_n498), .A3(G138), .A4(new_n463), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT69), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n495), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(new_n506), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n514), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n508), .A2(G51), .B1(new_n520), .B2(KEYINPUT70), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n521), .B1(KEYINPUT70), .B2(new_n520), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT5), .B(G543), .Z(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n506), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n527), .A2(G89), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n524), .A2(new_n525), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(new_n508), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n513), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n516), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n527), .A2(G81), .B1(new_n508), .B2(G43), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n526), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n562), .A2(new_n563), .B1(G91), .B2(new_n527), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  NAND2_X1  g141(.A1(new_n527), .A2(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n508), .A2(G49), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT74), .B1(new_n513), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n527), .A2(new_n573), .A3(G86), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n526), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n508), .B2(G48), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(G305));
  XNOR2_X1  g155(.A(KEYINPUT75), .B(G85), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n527), .A2(new_n581), .B1(new_n508), .B2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n516), .B2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n527), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  NAND2_X1  g162(.A1(new_n512), .A2(G66), .ZN(new_n588));
  INV_X1    g163(.A(G79), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT76), .B1(new_n589), .B2(new_n507), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n589), .A2(new_n507), .A3(KEYINPUT76), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n508), .B2(G54), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT77), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n585), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n585), .B1(new_n595), .B2(G868), .ZN(G321));
  NAND2_X1  g172(.A1(G168), .A2(G868), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G868), .B2(G299), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT78), .ZN(G297));
  XNOR2_X1  g175(.A(new_n599), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NOR2_X1   g178(.A1(new_n545), .A2(G868), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n595), .A2(new_n602), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n480), .A2(G2104), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  OAI22_X1  g187(.A1(new_n609), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n610), .B2(new_n609), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT80), .B2(G2100), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(new_n611), .A3(new_n612), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n480), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n482), .A2(G123), .ZN(new_n619));
  MUX2_X1   g194(.A(G99), .B(G111), .S(G2105), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G2104), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n616), .A2(new_n617), .A3(new_n624), .ZN(G156));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2427), .ZN(new_n629));
  INV_X1    g204(.A(G2430), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n632), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT17), .Z(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT81), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n644), .A2(new_n647), .ZN(new_n650));
  INV_X1    g225(.A(new_n643), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n650), .B(new_n646), .C1(new_n651), .C2(new_n647), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n645), .A3(new_n647), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n623), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n612), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  AOI211_X1 g242(.A(new_n665), .B(new_n667), .C1(new_n660), .C2(new_n664), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  MUX2_X1   g250(.A(G6), .B(G305), .S(G16), .Z(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT32), .B(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(G16), .A2(G22), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(G166), .B2(G16), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(G1971), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(G288), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT33), .B(G1976), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n686), .B(new_n687), .Z(new_n688));
  NOR3_X1   g263(.A1(new_n678), .A2(new_n682), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n683), .A2(G24), .ZN(new_n693));
  XNOR2_X1  g268(.A(G290), .B(KEYINPUT82), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n683), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT83), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G95), .B(G107), .S(G2105), .Z(new_n698));
  AOI22_X1  g273(.A1(G119), .A2(new_n482), .B1(new_n698), .B2(G2104), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n480), .A2(G131), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  NOR4_X1   g280(.A1(new_n691), .A2(new_n692), .A3(new_n697), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(KEYINPUT85), .A2(KEYINPUT36), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n683), .A2(G4), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n595), .B2(new_n683), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT86), .B(G1348), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G26), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n482), .A2(G128), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT90), .Z(new_n717));
  MUX2_X1   g292(.A(G104), .B(G116), .S(G2105), .Z(new_n718));
  AOI22_X1  g293(.A1(G140), .A2(new_n480), .B1(new_n718), .B2(G2104), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n715), .B1(new_n720), .B2(G29), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2067), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n683), .A2(G19), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT87), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n546), .B2(new_n683), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT88), .B(G1341), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT89), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n712), .A2(new_n722), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  NOR2_X1   g305(.A1(G168), .A2(new_n683), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n683), .B2(G21), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  AND2_X1   g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NOR2_X1   g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n713), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G160), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n713), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT92), .Z(new_n744));
  AND2_X1   g319(.A1(new_n713), .A2(G33), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n748), .A2(new_n749), .B1(new_n480), .B2(G139), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n463), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n745), .B1(new_n752), .B2(G29), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(G2072), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(G2072), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT30), .A2(G28), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT30), .A2(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n622), .B2(new_n713), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n755), .A2(new_n756), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n683), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n683), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1961), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n742), .B2(new_n741), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n744), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G29), .A2(G32), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT26), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n463), .A2(G2104), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(G105), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n480), .A2(G141), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n482), .A2(G129), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n769), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT93), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT27), .B(G1996), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G27), .A2(G29), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G164), .B2(G29), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G162), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G29), .B2(G35), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT29), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n683), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT23), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT96), .B(G1956), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n789), .A2(G2090), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n794), .ZN(new_n798));
  INV_X1    g373(.A(G2090), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n798), .A2(new_n795), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n781), .A2(new_n785), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n735), .A2(new_n736), .A3(new_n768), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n708), .A2(new_n730), .A3(new_n802), .ZN(G150));
  INV_X1    g378(.A(G150), .ZN(G311));
  NAND2_X1  g379(.A1(new_n508), .A2(G55), .ZN(new_n805));
  INV_X1    g380(.A(G93), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n513), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n516), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G860), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n595), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  INV_X1    g390(.A(new_n810), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(KEYINPUT97), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n810), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(new_n820), .B(new_n819), .S(new_n545), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n815), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT98), .Z(new_n825));
  OAI21_X1  g400(.A(new_n811), .B1(new_n823), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n813), .B1(new_n825), .B2(new_n826), .ZN(G145));
  AOI22_X1  g402(.A1(G130), .A2(new_n482), .B1(new_n480), .B2(G142), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n829), .A2(new_n463), .A3(G118), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n463), .B2(G118), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n828), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n609), .B(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n701), .B(KEYINPUT100), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n491), .A2(new_n492), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n498), .B1(new_n480), .B2(G138), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n776), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n836), .B(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n720), .B(new_n752), .Z(new_n843));
  AOI21_X1  g418(.A(KEYINPUT101), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n842), .B2(new_n843), .ZN(new_n845));
  XNOR2_X1  g420(.A(G160), .B(G162), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n622), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n845), .A2(new_n847), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g427(.A1(new_n816), .A2(G868), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n594), .B(G299), .Z(new_n854));
  INV_X1    g429(.A(KEYINPUT41), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(KEYINPUT102), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(KEYINPUT102), .B2(new_n857), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n605), .B(new_n821), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n854), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n861), .A2(KEYINPUT103), .B1(new_n862), .B2(new_n860), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(KEYINPUT103), .B2(new_n861), .ZN(new_n864));
  XNOR2_X1  g439(.A(G288), .B(KEYINPUT104), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G290), .ZN(new_n866));
  XOR2_X1   g441(.A(G303), .B(G305), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(KEYINPUT105), .ZN(new_n870));
  MUX2_X1   g445(.A(new_n869), .B(new_n870), .S(KEYINPUT42), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n864), .B(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n853), .B1(new_n872), .B2(G868), .ZN(G295));
  AOI21_X1  g448(.A(new_n853), .B1(new_n872), .B2(G868), .ZN(G331));
  XNOR2_X1  g449(.A(G286), .B(G301), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n821), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n859), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n862), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT106), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n876), .B2(new_n862), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(new_n870), .ZN(new_n883));
  INV_X1    g458(.A(new_n876), .ZN(new_n884));
  INV_X1    g459(.A(new_n856), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n857), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n870), .B1(new_n886), .B2(new_n878), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n849), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n882), .A2(new_n870), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n883), .A2(KEYINPUT43), .A3(new_n849), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT44), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(KEYINPUT43), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n883), .A2(new_n849), .A3(new_n891), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(KEYINPUT43), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n893), .B1(KEYINPUT44), .B2(new_n896), .ZN(G397));
  AOI21_X1  g472(.A(G1384), .B1(new_n500), .B2(new_n837), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(KEYINPUT45), .ZN(new_n899));
  INV_X1    g474(.A(G40), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n469), .A2(new_n476), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G2067), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n720), .B(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n776), .B(G1996), .Z(new_n906));
  AND2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n701), .B(new_n703), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(G290), .B(G1986), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n903), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g487(.A1(G303), .A2(G8), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT55), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n464), .ZN(new_n916));
  OAI21_X1  g491(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n465), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n918), .B2(G2105), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n919), .A2(G40), .A3(new_n474), .A4(new_n475), .ZN(new_n920));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n502), .A2(KEYINPUT50), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT50), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(G1384), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n799), .ZN(new_n928));
  INV_X1    g503(.A(G1971), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n840), .A2(KEYINPUT45), .A3(new_n921), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n901), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT45), .B1(new_n502), .B2(new_n921), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n927), .B1(new_n926), .B2(new_n799), .ZN(new_n935));
  OAI211_X1 g510(.A(G8), .B(new_n915), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n578), .A2(G651), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n508), .A2(G48), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n513), .A2(new_n571), .ZN(new_n941));
  OAI21_X1  g516(.A(G1981), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(G305), .B2(G1981), .ZN(new_n943));
  NOR2_X1   g518(.A1(KEYINPUT108), .A2(KEYINPUT49), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI221_X1 g520(.A(new_n942), .B1(KEYINPUT108), .B2(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n840), .A2(new_n921), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n920), .ZN(new_n948));
  INV_X1    g523(.A(G8), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1976), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT52), .B1(G288), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n950), .B(new_n953), .C1(new_n952), .C2(G288), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n901), .A2(new_n898), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n955), .B(G8), .C1(new_n952), .C2(G288), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT52), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n951), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n937), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n951), .A2(new_n952), .A3(new_n685), .ZN(new_n960));
  NOR2_X1   g535(.A1(G305), .A2(G1981), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n950), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n934), .A2(new_n935), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(new_n949), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n958), .B1(new_n965), .B2(new_n915), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT111), .B(new_n958), .C1(new_n965), .C2(new_n915), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n502), .A2(new_n921), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n502), .A2(KEYINPUT109), .A3(KEYINPUT45), .A4(new_n921), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n920), .B1(new_n947), .B2(new_n972), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n733), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n926), .A2(new_n742), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n979), .A2(G8), .A3(G168), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT63), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n937), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n968), .A2(new_n969), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT110), .B(KEYINPUT63), .Z(new_n984));
  NOR2_X1   g559(.A1(new_n947), .A2(new_n923), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT50), .B1(new_n502), .B2(new_n921), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n901), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n933), .B1(new_n987), .B2(G2090), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G8), .ZN(new_n989));
  INV_X1    g564(.A(new_n915), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n958), .A2(new_n991), .A3(new_n936), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n984), .B1(new_n992), .B2(new_n980), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n963), .B1(new_n983), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n926), .A2(KEYINPUT115), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n996), .B(new_n920), .C1(new_n922), .C2(new_n925), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n995), .A2(new_n997), .A3(G1961), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2078), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n931), .A2(new_n932), .A3(G2078), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(KEYINPUT53), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G171), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT119), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1006), .B(G171), .C1(new_n998), .C2(new_n1003), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n926), .A2(KEYINPUT115), .ZN(new_n1008));
  INV_X1    g583(.A(new_n997), .ZN(new_n1009));
  INV_X1    g584(.A(G1961), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1002), .A2(KEYINPUT53), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT120), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT53), .B1(new_n1013), .B2(G2078), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n1013), .B2(G2078), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n975), .A2(new_n930), .A3(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1011), .A2(G301), .A3(new_n1012), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1005), .A2(new_n1007), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n998), .A2(new_n1003), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n1022), .B2(G301), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1016), .B1(new_n1002), .B2(KEYINPUT53), .ZN(new_n1024));
  OAI21_X1  g599(.A(G171), .B1(new_n998), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n992), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT118), .B(G8), .C1(new_n979), .C2(G286), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT51), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT118), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n976), .A2(new_n733), .B1(new_n742), .B2(new_n926), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(G168), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(G168), .ZN(new_n1033));
  OAI21_X1  g608(.A(G8), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1028), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1020), .A2(new_n1021), .A3(new_n1026), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n560), .A2(new_n564), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n564), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT57), .B1(new_n559), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT112), .B(G1956), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n987), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n931), .A2(new_n932), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT56), .B(G2072), .Z(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT113), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT114), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n920), .B1(KEYINPUT45), .B2(new_n898), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n971), .A2(new_n972), .ZN(new_n1050));
  AND4_X1   g625(.A1(KEYINPUT114), .A2(new_n1049), .A3(new_n1050), .A4(new_n1047), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1044), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1049), .A2(new_n1050), .A3(KEYINPUT114), .A4(new_n1047), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(KEYINPUT116), .A3(new_n1044), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1042), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n955), .A2(G2067), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n995), .A2(new_n997), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(new_n711), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(new_n594), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  AOI221_X4 g643(.A(new_n1041), .B1(new_n987), .B2(new_n1043), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1042), .B1(new_n1059), .B2(new_n1044), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n594), .A2(KEYINPUT60), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n931), .A2(new_n932), .A3(G1996), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT58), .B(G1341), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n948), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n546), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n1077));
  NAND2_X1  g652(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n546), .B(new_n1078), .C1(new_n1073), .C2(new_n1075), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1064), .A2(new_n1072), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1066), .A2(KEYINPUT61), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1071), .B(new_n1080), .C1(new_n1061), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1064), .A2(new_n594), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1064), .A2(new_n594), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1067), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1036), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1011), .A2(new_n1001), .A3(new_n1012), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1025), .B(KEYINPUT54), .C1(new_n1089), .C2(G171), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n958), .A2(new_n991), .A3(new_n936), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n979), .A2(G286), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n977), .A2(G168), .A3(new_n978), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1030), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1095), .A2(G8), .B1(KEYINPUT51), .B2(new_n1027), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1021), .B1(new_n1097), .B2(new_n1020), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n912), .B(new_n994), .C1(new_n1088), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1035), .A2(KEYINPUT62), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1091), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1096), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1106), .A2(KEYINPUT123), .A3(new_n1102), .A4(new_n1091), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1104), .B(new_n1107), .C1(new_n1105), .C2(new_n1096), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1099), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1020), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1035), .A2(new_n1091), .A3(new_n1090), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT121), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n1036), .A3(new_n1087), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n912), .B1(new_n1113), .B2(new_n994), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n911), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n907), .A2(new_n700), .A3(new_n699), .A4(new_n703), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n717), .A2(new_n904), .A3(new_n719), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n902), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT124), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n902), .B1(new_n905), .B2(new_n777), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT46), .B1(new_n902), .B2(G1996), .ZN(new_n1121));
  OR3_X1    g696(.A1(new_n902), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1124));
  XNOR2_X1  g699(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  OR3_X1    g700(.A1(new_n902), .A2(G1986), .A3(G290), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT48), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1128), .B(new_n1129), .C1(new_n909), .C2(new_n903), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1119), .A2(new_n1125), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1115), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT126), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1115), .A2(new_n1134), .A3(new_n1131), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g711(.A1(new_n890), .A2(new_n892), .ZN(new_n1138));
  NAND4_X1  g712(.A1(new_n674), .A2(G319), .A3(new_n641), .A4(new_n657), .ZN(new_n1139));
  XNOR2_X1  g713(.A(new_n1139), .B(KEYINPUT127), .ZN(new_n1140));
  AND2_X1   g714(.A1(new_n1140), .A2(new_n851), .ZN(new_n1141));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1141), .ZN(G225));
  INV_X1    g716(.A(G225), .ZN(G308));
endmodule


