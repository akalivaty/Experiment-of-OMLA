//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(G8gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT17), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT90), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT89), .B(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT14), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n210), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n207), .A2(KEYINPUT90), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n217), .ZN(new_n221));
  AND4_X1   g020(.A1(new_n208), .A2(new_n218), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n218), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n206), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n206), .A2(KEYINPUT91), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n205), .B(G8gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT91), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n218), .A2(new_n221), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n224), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n232), .B(KEYINPUT13), .Z(new_n236));
  INV_X1    g035(.A(new_n231), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n229), .A2(new_n230), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n224), .A2(new_n231), .A3(KEYINPUT18), .A4(new_n232), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT11), .B(G169gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G197gat), .ZN(new_n243));
  XOR2_X1   g042(.A(G113gat), .B(G141gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n235), .A2(new_n239), .A3(new_n246), .A4(new_n240), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n248), .A2(KEYINPUT92), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT92), .B1(new_n248), .B2(new_n249), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(G155gat), .A2(G162gat), .ZN(new_n258));
  OR2_X1    g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(KEYINPUT2), .ZN(new_n260));
  INV_X1    g059(.A(G141gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(G148gat), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n262), .A2(KEYINPUT79), .ZN(new_n263));
  INV_X1    g062(.A(G148gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n254), .B2(new_n255), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n257), .B(new_n260), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G141gat), .B(G148gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n258), .B(new_n259), .C1(new_n267), .C2(KEYINPUT2), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT77), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n264), .A2(G141gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n262), .B2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(KEYINPUT77), .A3(new_n258), .A4(new_n259), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n266), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT66), .B(G120gat), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n283), .A2(G120gat), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n280), .B(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(G127gat), .A2(G134gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT65), .B(G127gat), .Z(new_n289));
  INV_X1    g088(.A(G134gat), .ZN(new_n290));
  OAI221_X1 g089(.A(new_n287), .B1(new_n288), .B2(KEYINPUT1), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n275), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n278), .A2(new_n279), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n275), .A2(KEYINPUT81), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n266), .A2(new_n270), .A3(new_n296), .A4(new_n274), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n286), .A2(new_n291), .A3(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n302), .A3(KEYINPUT4), .ZN(new_n303));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n275), .A2(new_n292), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n294), .A2(new_n303), .A3(new_n304), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT5), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n275), .B(new_n292), .ZN(new_n310));
  INV_X1    g109(.A(new_n304), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n298), .ZN(new_n314));
  INV_X1    g113(.A(new_n302), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n306), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n305), .A2(new_n306), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n311), .A2(KEYINPUT5), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n316), .A2(new_n294), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT0), .B(G57gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(G85gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n322), .B(new_n323), .Z(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n313), .A2(new_n319), .A3(new_n324), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n320), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT87), .ZN(new_n333));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT24), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(G183gat), .A3(G190gat), .ZN(new_n338));
  OR2_X1    g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(KEYINPUT24), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n336), .A2(new_n338), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n341), .A2(new_n342), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n346), .A2(KEYINPUT25), .A3(new_n338), .A4(new_n336), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT27), .B(G183gat), .ZN(new_n349));
  INV_X1    g148(.A(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n351), .A2(KEYINPUT28), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n351), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT64), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT26), .B1(new_n334), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n342), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n334), .A2(new_n354), .A3(KEYINPUT26), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n352), .A2(new_n353), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT29), .B1(new_n348), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT72), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363));
  INV_X1    g162(.A(G211gat), .ZN(new_n364));
  INV_X1    g163(.A(G218gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n363), .B1(KEYINPUT22), .B2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G211gat), .B(G218gat), .Z(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n358), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n361), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n362), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n369), .B(KEYINPUT71), .ZN(new_n373));
  INV_X1    g172(.A(new_n371), .ZN(new_n374));
  XOR2_X1   g173(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n361), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n373), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G8gat), .B(G36gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(G64gat), .ZN(new_n380));
  INV_X1    g179(.A(G92gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n372), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n369), .B1(new_n362), .B2(new_n371), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n374), .A2(new_n377), .A3(new_n373), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT37), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT37), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n388), .A3(new_n378), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n387), .A2(new_n382), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n332), .A2(new_n333), .A3(new_n384), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n378), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n372), .A2(new_n396), .A3(new_n378), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n388), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n389), .A2(new_n382), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n390), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n329), .A2(new_n392), .A3(new_n331), .A4(new_n384), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT87), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n404), .B(KEYINPUT83), .Z(new_n405));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n406));
  INV_X1    g205(.A(new_n369), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(new_n375), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n314), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n279), .A2(new_n376), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n407), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n405), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n373), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n369), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n406), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n369), .B2(new_n415), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n404), .B1(new_n419), .B2(new_n275), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n412), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n424), .B(G22gat), .Z(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n422), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n421), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n425), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n316), .A2(new_n294), .A3(new_n317), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n311), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT85), .B1(new_n310), .B2(new_n311), .ZN(new_n434));
  OR3_X1    g233(.A1(new_n310), .A2(KEYINPUT85), .A3(new_n311), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n433), .A2(KEYINPUT39), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT39), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n437), .A3(new_n311), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n324), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n383), .B1(new_n395), .B2(new_n397), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n384), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n384), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n440), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n441), .A2(new_n326), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n403), .A2(new_n431), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT68), .B1(new_n348), .B2(new_n358), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n315), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n348), .A2(KEYINPUT68), .A3(new_n358), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n315), .B1(new_n454), .B2(new_n452), .ZN(new_n455));
  INV_X1    g254(.A(G227gat), .ZN(new_n456));
  INV_X1    g255(.A(G233gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n453), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G43gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G71gat), .B(G99gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n464), .B(new_n465), .Z(new_n466));
  AOI21_X1  g265(.A(new_n459), .B1(new_n453), .B2(new_n455), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(KEYINPUT33), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n455), .ZN(new_n472));
  AOI221_X4 g271(.A(new_n469), .B1(KEYINPUT33), .B2(new_n466), .C1(new_n472), .C2(new_n458), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n463), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n458), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n478), .A3(new_n466), .ZN(new_n479));
  INV_X1    g278(.A(new_n473), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n462), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n474), .A2(new_n481), .A3(KEYINPUT69), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(new_n463), .C1(new_n471), .C2(new_n473), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT36), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n474), .A2(new_n481), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT70), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(new_n491), .A3(new_n488), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n486), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  OR3_X1    g292(.A1(new_n442), .A2(KEYINPUT75), .A3(new_n444), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT75), .B1(new_n442), .B2(new_n444), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n332), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n447), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n426), .A2(new_n430), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n451), .A2(new_n493), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n332), .A2(new_n448), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT88), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n487), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT88), .B1(new_n474), .B2(new_n481), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n431), .B(new_n503), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AND4_X1   g306(.A1(KEYINPUT35), .A2(new_n496), .A3(new_n497), .A4(new_n447), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n499), .B1(new_n484), .B2(new_n482), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n502), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n253), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G127gat), .B(G155gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n512), .B(KEYINPUT20), .Z(new_n513));
  XNOR2_X1  g312(.A(G57gat), .B(G64gat), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G71gat), .ZN(new_n516));
  INV_X1    g315(.A(G78gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G71gat), .A2(G78gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT9), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n519), .B(new_n518), .C1(new_n514), .C2(new_n521), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT21), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n225), .A2(new_n228), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(G211gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n525), .A2(KEYINPUT21), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(G211gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n513), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  INV_X1    g334(.A(new_n513), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G231gat), .A2(G233gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT19), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT93), .B(G183gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n534), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n222), .A2(new_n223), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT94), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n550), .B2(KEYINPUT7), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(KEYINPUT95), .A3(G85gat), .A4(G92gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n557), .A3(KEYINPUT7), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n552), .A2(new_n554), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(G99gat), .B2(G106gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n381), .A2(KEYINPUT96), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G99gat), .B(G106gat), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n569), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n559), .A2(new_n571), .A3(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n548), .B1(new_n549), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G134gat), .B(G162gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n230), .A2(new_n572), .A3(new_n570), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n574), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n546), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n545), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n541), .B1(new_n534), .B2(new_n537), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n542), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G204gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT99), .ZN(new_n590));
  INV_X1    g389(.A(G176gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT100), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n523), .A2(new_n524), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n559), .A2(new_n571), .A3(new_n567), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n571), .B1(new_n559), .B2(new_n567), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n570), .A2(new_n525), .A3(new_n572), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT97), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n570), .A2(new_n525), .A3(new_n603), .A4(new_n572), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n596), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI211_X1 g406(.A(KEYINPUT98), .B(KEYINPUT10), .C1(new_n602), .C2(new_n604), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n601), .A2(new_n606), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n595), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n605), .A2(new_n593), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n592), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  INV_X1    g414(.A(new_n592), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n617));
  INV_X1    g416(.A(new_n593), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n587), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n511), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n332), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g424(.A(KEYINPUT16), .B(G8gat), .Z(new_n626));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT102), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n626), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n448), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n631), .B2(new_n627), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n630), .B(KEYINPUT101), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n627), .A2(G8gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(G1325gat));
  INV_X1    g434(.A(G15gat), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n622), .A2(new_n636), .A3(new_n493), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n505), .A2(new_n506), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n636), .B2(new_n640), .ZN(G1326gat));
  NOR2_X1   g440(.A1(new_n622), .A2(new_n431), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT43), .B(G22gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1327gat));
  INV_X1    g443(.A(new_n584), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n501), .B2(new_n510), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n542), .A2(new_n585), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n620), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n646), .A2(new_n648), .A3(new_n649), .A4(new_n252), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n332), .A3(new_n211), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT45), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n645), .A2(KEYINPUT44), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n501), .A2(new_n510), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n501), .B2(new_n510), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n501), .A2(new_n510), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n584), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT44), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n620), .B(KEYINPUT103), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n248), .A2(new_n249), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n648), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT104), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n662), .A2(KEYINPUT106), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT106), .B1(new_n662), .B2(new_n667), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n497), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n653), .B1(new_n671), .B2(new_n211), .ZN(G1328gat));
  INV_X1    g471(.A(new_n448), .ZN(new_n673));
  OAI21_X1  g472(.A(G36gat), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n650), .A2(G36gat), .A3(new_n673), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(KEYINPUT107), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n674), .B(new_n677), .C1(new_n678), .C2(new_n675), .ZN(G1329gat));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n667), .ZN(new_n680));
  OAI21_X1  g479(.A(G43gat), .B1(new_n680), .B2(new_n493), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n650), .A2(G43gat), .A3(new_n638), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(KEYINPUT47), .A3(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(KEYINPUT108), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(KEYINPUT108), .ZN(new_n686));
  INV_X1    g485(.A(new_n493), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n668), .B2(new_n669), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n682), .B1(new_n688), .B2(G43gat), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n685), .B(new_n686), .C1(KEYINPUT47), .C2(new_n689), .ZN(G1330gat));
  OAI21_X1  g489(.A(G50gat), .B1(new_n680), .B2(new_n431), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n650), .A2(G50gat), .A3(new_n431), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(KEYINPUT48), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n499), .B1(new_n668), .B2(new_n669), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n692), .B1(new_n695), .B2(G50gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g496(.A1(new_n656), .A2(new_n657), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n587), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n663), .A2(new_n664), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n497), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT109), .B(G57gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1332gat));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n673), .ZN(new_n705));
  NOR2_X1   g504(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n706));
  AND2_X1   g505(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n705), .B2(new_n706), .ZN(G1333gat));
  OAI21_X1  g508(.A(new_n516), .B1(new_n701), .B2(new_n638), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n699), .A2(G71gat), .A3(new_n700), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n493), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g512(.A1(new_n701), .A2(new_n431), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(new_n517), .ZN(G1335gat));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n647), .A2(new_n664), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n646), .B2(KEYINPUT110), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n719), .B(new_n645), .C1(new_n501), .C2(new_n510), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n660), .A2(new_n719), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n646), .A2(KEYINPUT110), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n722), .A2(KEYINPUT51), .A3(new_n717), .A4(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n649), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n566), .A3(new_n332), .ZN(new_n726));
  INV_X1    g525(.A(new_n717), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n649), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n658), .B2(new_n661), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731), .B2(new_n497), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n726), .A2(new_n732), .ZN(G1336gat));
  INV_X1    g532(.A(new_n663), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n673), .A2(G92gat), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n727), .B1(new_n660), .B2(new_n719), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT51), .B1(new_n736), .B2(new_n723), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n718), .A2(new_n716), .A3(new_n720), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n734), .B(new_n735), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n662), .A2(new_n448), .A3(new_n728), .ZN(new_n740));
  INV_X1    g539(.A(new_n565), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n739), .B2(new_n742), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n565), .B1(new_n730), .B2(new_n448), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT52), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n742), .B2(KEYINPUT111), .ZN(new_n751));
  INV_X1    g550(.A(new_n735), .ZN(new_n752));
  AOI211_X1 g551(.A(new_n663), .B(new_n752), .C1(new_n721), .C2(new_n724), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT112), .B1(new_n753), .B2(new_n746), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n749), .A2(new_n756), .ZN(G1337gat));
  INV_X1    g556(.A(G99gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n725), .A2(new_n758), .A3(new_n639), .ZN(new_n759));
  OAI21_X1  g558(.A(G99gat), .B1(new_n731), .B2(new_n493), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1338gat));
  OAI21_X1  g560(.A(G106gat), .B1(new_n731), .B2(new_n431), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n431), .A2(G106gat), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n734), .B(new_n763), .C1(new_n737), .C2(new_n738), .ZN(new_n764));
  NAND2_X1  g563(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n766), .B(new_n767), .Z(G1339gat));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n605), .A2(new_n606), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT98), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n605), .A2(new_n596), .A3(new_n606), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n771), .A2(new_n595), .A3(new_n611), .A4(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(KEYINPUT54), .C1(new_n617), .C2(new_n618), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n611), .A3(new_n772), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n776), .A3(new_n594), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n774), .A2(KEYINPUT55), .A3(new_n592), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n619), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n616), .B1(new_n612), .B2(new_n776), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT55), .B1(new_n780), .B2(new_n774), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n769), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  INV_X1    g582(.A(new_n774), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n777), .A2(new_n592), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(KEYINPUT114), .A3(new_n619), .A4(new_n778), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(new_n664), .A3(new_n787), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n237), .A2(new_n238), .A3(new_n236), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n232), .B1(new_n224), .B2(new_n231), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n245), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n249), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n620), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n788), .A2(KEYINPUT115), .A3(new_n793), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(new_n645), .A3(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n584), .A2(new_n792), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n782), .A3(new_n787), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n647), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n587), .A2(new_n620), .A3(new_n664), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n497), .A2(new_n448), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n509), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n283), .A3(new_n664), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n638), .A2(new_n499), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n253), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(G1340gat));
  OR3_X1    g611(.A1(new_n806), .A2(new_n282), .A3(new_n649), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n805), .A2(new_n809), .A3(new_n734), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(G120gat), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n814), .B2(G120gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(G1341gat));
  NOR3_X1   g618(.A1(new_n810), .A2(new_n289), .A3(new_n648), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n807), .A2(new_n647), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n289), .B2(new_n821), .ZN(G1342gat));
  NOR3_X1   g621(.A1(new_n806), .A2(G134gat), .A3(new_n645), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n810), .B2(new_n645), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(G1343gat));
  OAI21_X1  g627(.A(new_n499), .B1(new_n801), .B2(new_n802), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n493), .A2(new_n804), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n253), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT58), .B1(new_n834), .B2(new_n261), .ZN(new_n835));
  INV_X1    g634(.A(new_n256), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n779), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n780), .B2(new_n774), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n780), .A2(new_n840), .A3(new_n774), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n783), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n252), .B(new_n839), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n584), .B1(new_n844), .B2(new_n793), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n647), .B1(new_n846), .B2(new_n800), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n499), .B1(new_n847), .B2(new_n802), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n831), .B1(new_n848), .B2(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n838), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n836), .B1(new_n850), .B2(new_n253), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n838), .A2(new_n664), .A3(new_n849), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n836), .A2(new_n853), .B1(new_n834), .B2(new_n261), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(G1344gat));
  NOR3_X1   g655(.A1(new_n833), .A2(G148gat), .A3(new_n649), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT118), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n253), .A2(new_n586), .A3(new_n649), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n799), .A2(new_n839), .A3(new_n786), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n648), .B1(new_n845), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g663(.A(KEYINPUT57), .B(new_n431), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n829), .B2(KEYINPUT57), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n620), .A3(new_n832), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n264), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n859), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n850), .A2(new_n649), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(KEYINPUT59), .A3(new_n264), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n858), .B1(new_n871), .B2(new_n873), .ZN(G1345gat));
  INV_X1    g673(.A(G155gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n850), .A2(new_n875), .A3(new_n648), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n833), .A2(new_n648), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT121), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(new_n875), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n850), .B2(new_n645), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n645), .A2(G162gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n833), .B2(new_n881), .ZN(G1347gat));
  AND2_X1   g681(.A1(new_n803), .A2(new_n509), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n673), .A2(new_n332), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(G169gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n664), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n639), .A2(new_n884), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT122), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n803), .A2(new_n431), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891), .B2(new_n253), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n888), .A2(new_n892), .ZN(G1348gat));
  NOR3_X1   g692(.A1(new_n891), .A2(new_n591), .A3(new_n663), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n886), .A2(new_n620), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n591), .ZN(G1349gat));
  NAND4_X1  g695(.A1(new_n883), .A2(new_n647), .A3(new_n349), .A4(new_n884), .ZN(new_n897));
  OAI21_X1  g696(.A(G183gat), .B1(new_n891), .B2(new_n648), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n897), .A2(new_n898), .B1(KEYINPUT123), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(KEYINPUT123), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n900), .B(new_n901), .ZN(G1350gat));
  AND4_X1   g701(.A1(new_n350), .A2(new_n883), .A3(new_n584), .A4(new_n884), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT124), .ZN(new_n904));
  OAI21_X1  g703(.A(G190gat), .B1(new_n891), .B2(new_n645), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1351gat));
  INV_X1    g706(.A(G197gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n493), .A2(new_n884), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n830), .A2(new_n908), .A3(new_n664), .A4(new_n910), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT125), .Z(new_n912));
  NAND2_X1  g711(.A1(new_n866), .A2(new_n910), .ZN(new_n913));
  OAI21_X1  g712(.A(G197gat), .B1(new_n913), .B2(new_n253), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n830), .A2(new_n910), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n916), .A2(G204gat), .A3(new_n649), .ZN(new_n917));
  AND2_X1   g716(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n918));
  NOR2_X1   g717(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G204gat), .B1(new_n913), .B2(new_n663), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n920), .B(new_n921), .C1(new_n918), .C2(new_n917), .ZN(G1353gat));
  NAND2_X1  g721(.A1(new_n829), .A2(KEYINPUT57), .ZN(new_n923));
  INV_X1    g722(.A(new_n865), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n923), .A2(new_n647), .A3(new_n924), .A4(new_n910), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n866), .A2(KEYINPUT127), .A3(new_n647), .A4(new_n910), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(G211gat), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n927), .A2(KEYINPUT63), .A3(new_n928), .A4(G211gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n830), .A2(new_n364), .A3(new_n647), .A4(new_n910), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1354gat));
  OAI21_X1  g734(.A(G218gat), .B1(new_n913), .B2(new_n645), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n584), .A2(new_n365), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n916), .B2(new_n937), .ZN(G1355gat));
endmodule


