//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT64), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT65), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G137), .A3(new_n460), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(new_n460), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(G160));
  NAND2_X1  g044(.A1(new_n464), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(new_n460), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  AOI22_X1  g048(.A1(G124), .A2(new_n471), .B1(new_n473), .B2(G136), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(KEYINPUT66), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(KEYINPUT66), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT67), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OAI21_X1  g056(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(G114), .B2(new_n460), .ZN(new_n484));
  INV_X1    g059(.A(G126), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n470), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT4), .B1(new_n472), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n464), .A2(new_n489), .A3(G138), .A4(new_n460), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(G164));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G651), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(G651), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(G543), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G50), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n505), .A2(new_n495), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n497), .A2(new_n498), .A3(new_n504), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G88), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n501), .A2(new_n506), .A3(new_n509), .ZN(G303));
  INV_X1    g085(.A(G303), .ZN(G166));
  NOR2_X1   g086(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n494), .B2(new_n496), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(G89), .A3(new_n504), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n497), .A2(G51), .A3(G543), .A4(new_n498), .ZN(new_n515));
  AND2_X1   g090(.A1(G63), .A2(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT7), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n519), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n504), .A2(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n514), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(G168));
  INV_X1    g098(.A(G64), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(new_n502), .B2(new_n503), .ZN(new_n525));
  AND2_X1   g100(.A1(G77), .A2(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n497), .A2(G90), .A3(new_n504), .A4(new_n498), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n497), .A2(G52), .A3(G543), .A4(new_n498), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G171));
  INV_X1    g106(.A(G56), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n502), .B2(new_n503), .ZN(new_n533));
  AND2_X1   g108(.A1(G68), .A2(G543), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n497), .A2(G81), .A3(new_n504), .A4(new_n498), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n497), .A2(G43), .A3(G543), .A4(new_n498), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  AND2_X1   g118(.A1(G53), .A2(G543), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n495), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT68), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n498), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(KEYINPUT9), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT9), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n513), .B2(new_n544), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT69), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n497), .A2(G91), .A3(new_n504), .A4(new_n498), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n513), .A2(KEYINPUT70), .A3(G91), .A4(new_n504), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT5), .A2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(KEYINPUT5), .A2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g139(.A(KEYINPUT71), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(G651), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n547), .A2(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n513), .A2(new_n549), .A3(new_n544), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n551), .A2(new_n556), .A3(new_n566), .A4(new_n570), .ZN(G299));
  NAND2_X1  g146(.A1(new_n530), .A2(KEYINPUT72), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT72), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G301));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n522), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT73), .A4(new_n521), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G286));
  NAND2_X1  g156(.A1(new_n500), .A2(G49), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n508), .A2(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND3_X1  g160(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n507), .B2(new_n587), .C1(new_n495), .C2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n495), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT74), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n508), .A2(G85), .B1(new_n500), .B2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n507), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n513), .A2(KEYINPUT10), .A3(G92), .A4(new_n504), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(G66), .B1(new_n558), .B2(new_n559), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n495), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n500), .B2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n575), .ZN(G321));
  XNOR2_X1  g181(.A(G321), .B(KEYINPUT75), .ZN(G284));
  MUX2_X1   g182(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g183(.A(G297), .B(KEYINPUT76), .ZN(G280));
  AOI22_X1  g184(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n495), .A2(new_n610), .B1(new_n499), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n597), .B2(new_n598), .ZN(new_n613));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND3_X1  g190(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n604), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n471), .A2(G123), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT77), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G2105), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(new_n473), .B2(G135), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n462), .A2(new_n464), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n629), .A2(new_n634), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT78), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n650), .B(G14), .C1(new_n648), .C2(new_n647), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(G401));
  NOR2_X1   g227(.A1(G2072), .A2(G2078), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n442), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT17), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT80), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT81), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n654), .ZN(new_n661));
  INV_X1    g236(.A(new_n658), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n662), .C1(new_n655), .C2(new_n657), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n657), .A2(new_n654), .A3(new_n662), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n670), .C2(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT82), .ZN(new_n679));
  XOR2_X1   g254(.A(G1981), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n679), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1971), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(KEYINPUT90), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(KEYINPUT90), .ZN(new_n691));
  NOR2_X1   g266(.A1(G16), .A2(G23), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G288), .B2(new_n686), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT33), .B(G1976), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  MUX2_X1   g271(.A(G6), .B(G305), .S(G16), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT32), .B(G1981), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT88), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT87), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n697), .B(new_n700), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n690), .A2(new_n691), .A3(new_n696), .A4(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n703));
  OR2_X1    g278(.A1(G16), .A2(G24), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G290), .B2(new_n686), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT85), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(G25), .A2(G29), .ZN(new_n711));
  OR2_X1    g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT83), .Z(new_n714));
  INV_X1    g289(.A(G119), .ZN(new_n715));
  INV_X1    g290(.A(G131), .ZN(new_n716));
  OAI22_X1  g291(.A1(new_n715), .A2(new_n470), .B1(new_n472), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n711), .B1(new_n718), .B2(G29), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT84), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n709), .A2(new_n710), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n703), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT36), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n727), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT29), .Z(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n686), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n686), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT94), .B(G1966), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n686), .A2(G5), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G171), .B2(new_n686), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G1961), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(G1961), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n735), .A2(new_n737), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n738), .A2(new_n741), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n732), .A2(new_n733), .A3(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n686), .A2(G20), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G299), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n686), .ZN(new_n750));
  INV_X1    g325(.A(G1956), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT31), .B(G11), .Z(new_n753));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n727), .B1(new_n754), .B2(G28), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT95), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n756), .A2(KEYINPUT95), .B1(new_n754), .B2(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n753), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n628), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n727), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT96), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n473), .A2(G141), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n471), .A2(G129), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n462), .A2(G105), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT26), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(new_n727), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n727), .B2(G32), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  INV_X1    g350(.A(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G160), .B2(new_n727), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G2084), .ZN(new_n780));
  NOR2_X1   g355(.A1(G164), .A2(new_n727), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G27), .B2(new_n727), .ZN(new_n782));
  INV_X1    g357(.A(G2078), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n779), .A2(G2084), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT97), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n774), .A2(new_n780), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n782), .A2(new_n783), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n788), .B1(KEYINPUT97), .B2(new_n785), .C1(new_n772), .C2(new_n773), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n727), .A2(G33), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n473), .A2(G139), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT92), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT25), .Z(new_n794));
  AOI22_X1  g369(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n460), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(new_n727), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2072), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n762), .A2(new_n787), .A3(new_n789), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n686), .A2(G4), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n613), .B2(new_n686), .ZN(new_n802));
  INV_X1    g377(.A(G1348), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n473), .A2(G140), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n471), .A2(G128), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n460), .A2(G116), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n805), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G29), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n727), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G2067), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n686), .A2(G19), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n538), .B2(new_n686), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G1341), .Z(new_n818));
  NAND3_X1  g393(.A1(new_n804), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT91), .Z(new_n820));
  AND4_X1   g395(.A1(new_n745), .A2(new_n752), .A3(new_n800), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n726), .A2(new_n821), .ZN(G150));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n823));
  XNOR2_X1  g398(.A(G150), .B(new_n823), .ZN(G311));
  NAND4_X1  g399(.A1(new_n497), .A2(G55), .A3(G543), .A4(new_n498), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n497), .A2(G93), .A3(new_n504), .A4(new_n498), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT100), .B1(new_n829), .B2(new_n495), .ZN(new_n830));
  OAI21_X1  g405(.A(G67), .B1(new_n558), .B2(new_n559), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n833), .A2(new_n834), .A3(G651), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n827), .A2(new_n828), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT102), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n828), .B1(new_n825), .B2(new_n826), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n836), .A2(new_n837), .A3(new_n538), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n538), .A2(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n616), .A2(KEYINPUT102), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n834), .B1(new_n833), .B2(G651), .ZN(new_n844));
  AOI211_X1 g419(.A(KEYINPUT100), .B(new_n495), .C1(new_n831), .C2(new_n832), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n841), .B(new_n842), .C1(new_n846), .C2(new_n838), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT38), .Z(new_n849));
  NOR2_X1   g424(.A1(new_n604), .A2(new_n614), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n846), .A2(new_n838), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT103), .ZN(G145));
  NAND2_X1  g435(.A1(new_n488), .A2(new_n490), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n486), .A2(KEYINPUT104), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n863), .B(new_n484), .C1(new_n470), .C2(new_n485), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n809), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n770), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n797), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n718), .B(new_n631), .ZN(new_n869));
  OR2_X1    g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n871));
  INV_X1    g446(.A(G130), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n470), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(G142), .B2(new_n473), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n869), .B(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n868), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n876), .B2(new_n868), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n628), .B(G160), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n480), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n881), .B2(new_n879), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n856), .A2(new_n617), .ZN(new_n885));
  XNOR2_X1  g460(.A(G290), .B(G305), .ZN(new_n886));
  XOR2_X1   g461(.A(G303), .B(G288), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT42), .Z(new_n889));
  XOR2_X1   g464(.A(new_n848), .B(new_n619), .Z(new_n890));
  AND3_X1   g465(.A1(G299), .A2(KEYINPUT106), .A3(new_n613), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n565), .A2(G651), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n896), .A2(new_n564), .B1(new_n554), .B2(new_n555), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n897), .A3(new_n604), .ZN(new_n898));
  NAND2_X1  g473(.A1(G299), .A2(new_n613), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n892), .A2(new_n901), .A3(KEYINPUT107), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT107), .B1(new_n892), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n890), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n898), .A2(new_n899), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n749), .A2(KEYINPUT108), .A3(new_n604), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n892), .B2(new_n901), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n904), .B1(new_n912), .B2(new_n890), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n889), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n885), .B1(new_n914), .B2(new_n617), .ZN(G295));
  OAI21_X1  g490(.A(new_n885), .B1(new_n914), .B2(new_n617), .ZN(G331));
  NAND3_X1  g491(.A1(new_n578), .A2(G171), .A3(new_n579), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n572), .A2(G168), .A3(new_n574), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n848), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n840), .A3(new_n847), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n892), .A2(new_n901), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n919), .A2(new_n840), .A3(new_n847), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n919), .B1(new_n840), .B2(new_n847), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n922), .A2(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n925), .B1(new_n911), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n888), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n900), .B1(G299), .B2(new_n613), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n604), .B1(new_n895), .B2(new_n897), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n907), .B1(new_n940), .B2(new_n891), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n906), .A2(new_n908), .A3(KEYINPUT41), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n923), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n941), .A2(new_n923), .A3(KEYINPUT110), .A4(new_n942), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n929), .B(new_n930), .C1(new_n902), .C2(new_n903), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n948), .A2(KEYINPUT111), .A3(new_n888), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT111), .B1(new_n948), .B2(new_n888), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n935), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n937), .B1(new_n951), .B2(KEYINPUT43), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n932), .A2(new_n933), .ZN(new_n956));
  INV_X1    g531(.A(G37), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n948), .A2(new_n888), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n948), .A2(KEYINPUT111), .A3(new_n888), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n955), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n951), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n934), .A2(new_n935), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT44), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT113), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n972), .B(new_n969), .C1(new_n965), .C2(new_n966), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n954), .B1(new_n971), .B2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n865), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT114), .B(G40), .Z(new_n979));
  NOR3_X1   g554(.A1(new_n466), .A2(new_n468), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n770), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(G1996), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n809), .B(new_n814), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n982), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n987), .B1(new_n992), .B2(new_n770), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n718), .B(new_n721), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(new_n983), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(G290), .A2(G1986), .ZN(new_n996));
  NAND2_X1  g571(.A1(G290), .A2(G1986), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n983), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  INV_X1    g575(.A(new_n486), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n861), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n975), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n865), .A2(new_n1005), .A3(new_n975), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(new_n980), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(G2084), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n978), .A2(KEYINPUT120), .A3(new_n980), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n865), .B2(new_n975), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n981), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n861), .B2(new_n1001), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT45), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1008), .B1(new_n1015), .B2(new_n736), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1000), .B1(new_n1016), .B2(G168), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(G168), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT51), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n865), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n980), .B1(new_n1013), .B2(KEYINPUT45), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT116), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n865), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n977), .B1(G164), .B2(G1384), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n980), .A4(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT117), .B(G1971), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1007), .A2(G2090), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XOR2_X1   g610(.A(new_n1035), .B(KEYINPUT55), .Z(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  OR2_X1    g613(.A1(G288), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n980), .A2(new_n975), .A3(new_n865), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1039), .A2(new_n1040), .A3(new_n1043), .A4(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G305), .A2(G1981), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n588), .A2(new_n495), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n508), .A2(G86), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n586), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1047), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1040), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1046), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n1047), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1040), .A2(G8), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(KEYINPUT119), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1045), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n980), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1005), .B1(new_n865), .B2(new_n975), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n1064), .A2(G2090), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1000), .B1(new_n1032), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1037), .B(new_n1063), .C1(new_n1036), .C2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(G2078), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1006), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n980), .B1(new_n1013), .B2(new_n1005), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT122), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1004), .A2(new_n1075), .A3(new_n1006), .A4(new_n980), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT123), .B(G1961), .Z(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n466), .A2(KEYINPUT124), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n466), .A2(KEYINPUT124), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1069), .A2(G2078), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G40), .ZN(new_n1082));
  NOR4_X1   g657(.A1(new_n1079), .A2(new_n1080), .A3(new_n468), .A4(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(new_n1027), .A3(new_n978), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1071), .A2(G301), .A3(new_n1078), .A4(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1009), .A2(new_n1012), .A3(new_n1081), .A4(new_n1014), .ZN(new_n1086));
  AOI21_X1  g661(.A(G2078), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1078), .B(new_n1086), .C1(new_n1087), .C2(KEYINPUT53), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n575), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1068), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n751), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n749), .A2(KEYINPUT57), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n567), .A2(KEYINPUT121), .A3(new_n569), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n548), .B2(new_n550), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n897), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1094), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1027), .A2(new_n980), .A3(new_n1029), .A4(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1093), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1074), .A2(new_n803), .A3(new_n1076), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1040), .A2(G2067), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n604), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1101), .B1(new_n1093), .B2(new_n1103), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1104), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1110), .B1(new_n1111), .B2(new_n1108), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1093), .A2(new_n1103), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n1100), .A3(new_n1094), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1027), .A2(new_n988), .A3(new_n980), .A4(new_n1029), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT58), .B(G1341), .Z(new_n1117));
  NAND2_X1  g692(.A1(new_n1040), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n616), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1105), .A2(KEYINPUT60), .A3(new_n604), .A4(new_n1106), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1112), .A2(new_n1115), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1105), .A2(KEYINPUT60), .A3(new_n1106), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT60), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n604), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1109), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1088), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1091), .B1(new_n1128), .B2(G301), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1078), .B(new_n1084), .C1(new_n1087), .C2(KEYINPUT53), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(G171), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1092), .A2(new_n1127), .A3(new_n1135), .ZN(new_n1136));
  OR3_X1    g711(.A1(new_n1068), .A2(KEYINPUT62), .A3(new_n1089), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1023), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1068), .A2(new_n1089), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1139), .A2(new_n1020), .A3(KEYINPUT62), .A4(new_n1022), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1016), .A2(new_n1000), .A3(G286), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1068), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1037), .A2(new_n1063), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1000), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1146), .A2(new_n1036), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1145), .A2(KEYINPUT63), .A3(new_n1142), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1063), .A2(new_n1036), .A3(new_n1146), .ZN(new_n1150));
  AOI211_X1 g725(.A(G1976), .B(G288), .C1(new_n1057), .C2(new_n1062), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1052), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1061), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1140), .A2(new_n1149), .A3(new_n1150), .A4(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n999), .B1(new_n1138), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n986), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n982), .B1(new_n1156), .B2(new_n984), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n991), .A2(KEYINPUT46), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n991), .A2(KEYINPUT46), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT47), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1163));
  OAI211_X1 g738(.A(KEYINPUT47), .B(new_n1157), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n809), .A2(G2067), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n714), .A2(new_n721), .A3(new_n717), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n993), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n983), .A2(new_n996), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT48), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n1169), .A2(new_n983), .B1(new_n995), .B2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1165), .A2(new_n1166), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1155), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1155), .A2(new_n1173), .A3(KEYINPUT127), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(G319), .ZN(new_n1180));
  NOR4_X1   g754(.A1(G401), .A2(new_n1180), .A3(G227), .A4(G229), .ZN(new_n1181));
  AND3_X1   g755(.A1(new_n1181), .A2(new_n883), .A3(new_n952), .ZN(G308));
  NAND3_X1  g756(.A1(new_n1181), .A2(new_n883), .A3(new_n952), .ZN(G225));
endmodule


