

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578;

  XOR2_X1 U322 ( .A(G78GAT), .B(G148GAT), .Z(n290) );
  NOR2_X1 U323 ( .A1(n573), .A2(n496), .ZN(n497) );
  NOR2_X1 U324 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U325 ( .A(n331), .B(n330), .ZN(n336) );
  XNOR2_X1 U326 ( .A(n336), .B(n335), .ZN(n340) );
  NOR2_X1 U327 ( .A1(n547), .A2(n546), .ZN(n559) );
  XOR2_X1 U328 ( .A(n373), .B(n372), .Z(n547) );
  XOR2_X1 U329 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n292) );
  XNOR2_X1 U330 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n291) );
  XNOR2_X1 U331 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U332 ( .A(G57GAT), .B(G148GAT), .Z(n294) );
  XNOR2_X1 U333 ( .A(G141GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U335 ( .A(n296), .B(n295), .ZN(n311) );
  XOR2_X1 U336 ( .A(G155GAT), .B(KEYINPUT2), .Z(n298) );
  XNOR2_X1 U337 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n297) );
  XNOR2_X1 U338 ( .A(n298), .B(n297), .ZN(n376) );
  XOR2_X1 U339 ( .A(G85GAT), .B(n376), .Z(n300) );
  NAND2_X1 U340 ( .A1(G225GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U341 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U342 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n302) );
  XNOR2_X1 U343 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U345 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U346 ( .A(KEYINPUT85), .B(G134GAT), .Z(n306) );
  XNOR2_X1 U347 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n305) );
  XNOR2_X1 U348 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U349 ( .A(G113GAT), .B(n307), .Z(n372) );
  XNOR2_X1 U350 ( .A(G29GAT), .B(n372), .ZN(n308) );
  XNOR2_X1 U351 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U352 ( .A(n311), .B(n310), .ZN(n542) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G1GAT), .Z(n418) );
  XOR2_X1 U354 ( .A(G169GAT), .B(G8GAT), .Z(n352) );
  XOR2_X1 U355 ( .A(n418), .B(n352), .Z(n313) );
  NAND2_X1 U356 ( .A1(G229GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U358 ( .A(G141GAT), .B(G22GAT), .Z(n377) );
  XOR2_X1 U359 ( .A(n314), .B(n377), .Z(n322) );
  XOR2_X1 U360 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n316) );
  XNOR2_X1 U361 ( .A(G113GAT), .B(G197GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U363 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n318) );
  XNOR2_X1 U364 ( .A(KEYINPUT71), .B(KEYINPUT68), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U367 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U368 ( .A(G29GAT), .B(KEYINPUT8), .Z(n324) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G36GAT), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U371 ( .A(G50GAT), .B(KEYINPUT7), .Z(n325) );
  XNOR2_X1 U372 ( .A(n326), .B(n325), .ZN(n425) );
  XOR2_X1 U373 ( .A(n327), .B(n425), .Z(n527) );
  INV_X1 U374 ( .A(n527), .ZN(n565) );
  XOR2_X1 U375 ( .A(n565), .B(KEYINPUT72), .Z(n502) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n290), .B(n328), .ZN(n380) );
  XNOR2_X1 U378 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n329), .B(KEYINPUT13), .ZN(n417) );
  XNOR2_X1 U380 ( .A(n380), .B(n417), .ZN(n331) );
  XOR2_X1 U381 ( .A(G99GAT), .B(G85GAT), .Z(n430) );
  INV_X1 U382 ( .A(n430), .ZN(n330) );
  XOR2_X1 U383 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n333) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U386 ( .A(n334), .B(KEYINPUT33), .Z(n335) );
  XOR2_X1 U387 ( .A(G120GAT), .B(G71GAT), .Z(n367) );
  XOR2_X1 U388 ( .A(G64GAT), .B(G92GAT), .Z(n338) );
  XNOR2_X1 U389 ( .A(G176GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n348) );
  XNOR2_X1 U391 ( .A(n367), .B(n348), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n569) );
  NOR2_X1 U393 ( .A1(n502), .A2(n569), .ZN(n460) );
  XNOR2_X1 U394 ( .A(KEYINPUT19), .B(KEYINPUT88), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n341), .B(G183GAT), .ZN(n342) );
  XOR2_X1 U396 ( .A(n342), .B(KEYINPUT89), .Z(n344) );
  XNOR2_X1 U397 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n371) );
  XOR2_X1 U399 ( .A(KEYINPUT21), .B(G218GAT), .Z(n346) );
  XNOR2_X1 U400 ( .A(KEYINPUT91), .B(G211GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U402 ( .A(G197GAT), .B(n347), .Z(n386) );
  XNOR2_X1 U403 ( .A(n371), .B(n386), .ZN(n356) );
  XOR2_X1 U404 ( .A(G190GAT), .B(KEYINPUT77), .Z(n429) );
  XOR2_X1 U405 ( .A(n429), .B(n348), .Z(n350) );
  NAND2_X1 U406 ( .A1(G226GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U408 ( .A(n351), .B(KEYINPUT96), .Z(n354) );
  XNOR2_X1 U409 ( .A(G36GAT), .B(n352), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n539) );
  XNOR2_X1 U412 ( .A(n539), .B(KEYINPUT97), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n357), .B(KEYINPUT27), .ZN(n396) );
  INV_X1 U414 ( .A(n542), .ZN(n401) );
  NAND2_X1 U415 ( .A1(n396), .A2(n401), .ZN(n509) );
  XOR2_X1 U416 ( .A(KEYINPUT87), .B(G190GAT), .Z(n359) );
  XNOR2_X1 U417 ( .A(G43GAT), .B(G99GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U419 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n361) );
  XNOR2_X1 U420 ( .A(G169GAT), .B(G15GAT), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U422 ( .A(n363), .B(n362), .Z(n369) );
  XOR2_X1 U423 ( .A(KEYINPUT90), .B(G176GAT), .Z(n365) );
  NAND2_X1 U424 ( .A1(G227GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n373) );
  XNOR2_X1 U429 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n388) );
  XOR2_X1 U430 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n375) );
  XNOR2_X1 U431 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n385) );
  XOR2_X1 U433 ( .A(n377), .B(n376), .Z(n379) );
  NAND2_X1 U434 ( .A1(G228GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U436 ( .A(n381), .B(n380), .Z(n383) );
  XNOR2_X1 U437 ( .A(KEYINPUT92), .B(G204GAT), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U440 ( .A(n387), .B(n386), .Z(n544) );
  XNOR2_X1 U441 ( .A(n388), .B(n544), .ZN(n510) );
  NAND2_X1 U442 ( .A1(n547), .A2(n510), .ZN(n389) );
  NOR2_X1 U443 ( .A1(n509), .A2(n389), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n390), .B(KEYINPUT98), .ZN(n403) );
  XNOR2_X1 U445 ( .A(KEYINPUT25), .B(KEYINPUT100), .ZN(n393) );
  NOR2_X1 U446 ( .A1(n539), .A2(n547), .ZN(n391) );
  NOR2_X1 U447 ( .A1(n544), .A2(n391), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U449 ( .A(KEYINPUT26), .B(KEYINPUT99), .Z(n395) );
  NAND2_X1 U450 ( .A1(n544), .A2(n547), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n564) );
  INV_X1 U452 ( .A(n564), .ZN(n525) );
  NAND2_X1 U453 ( .A1(n396), .A2(n525), .ZN(n397) );
  NAND2_X1 U454 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U455 ( .A(KEYINPUT101), .B(n399), .ZN(n400) );
  NOR2_X1 U456 ( .A1(n401), .A2(n400), .ZN(n402) );
  NOR2_X1 U457 ( .A1(n403), .A2(n402), .ZN(n457) );
  XOR2_X1 U458 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n444) );
  XOR2_X1 U459 ( .A(G78GAT), .B(G211GAT), .Z(n405) );
  XNOR2_X1 U460 ( .A(G22GAT), .B(G127GAT), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U462 ( .A(KEYINPUT82), .B(KEYINPUT78), .Z(n407) );
  XNOR2_X1 U463 ( .A(G155GAT), .B(KEYINPUT81), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U465 ( .A(n409), .B(n408), .Z(n414) );
  XOR2_X1 U466 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n411) );
  NAND2_X1 U467 ( .A1(G231GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(KEYINPUT12), .B(n412), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n424) );
  XOR2_X1 U471 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n416) );
  XNOR2_X1 U472 ( .A(G8GAT), .B(G64GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n422) );
  XOR2_X1 U474 ( .A(n417), .B(G71GAT), .Z(n420) );
  XNOR2_X1 U475 ( .A(n418), .B(G183GAT), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U477 ( .A(n422), .B(n421), .Z(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n573) );
  INV_X1 U479 ( .A(n425), .ZN(n442) );
  XOR2_X1 U480 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n427) );
  NAND2_X1 U481 ( .A1(G232GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT10), .B(n428), .ZN(n440) );
  XOR2_X1 U484 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n432) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U487 ( .A(KEYINPUT75), .B(G92GAT), .Z(n434) );
  XNOR2_X1 U488 ( .A(G134GAT), .B(G106GAT), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(n436), .B(n435), .Z(n438) );
  XNOR2_X1 U491 ( .A(G218GAT), .B(G162GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U494 ( .A(n442), .B(n441), .Z(n558) );
  INV_X1 U495 ( .A(n558), .ZN(n536) );
  NAND2_X1 U496 ( .A1(n573), .A2(n536), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n445), .B(KEYINPUT16), .ZN(n446) );
  NOR2_X1 U499 ( .A1(n457), .A2(n446), .ZN(n472) );
  NAND2_X1 U500 ( .A1(n460), .A2(n472), .ZN(n454) );
  NOR2_X1 U501 ( .A1(n542), .A2(n454), .ZN(n448) );
  XNOR2_X1 U502 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U504 ( .A(G1GAT), .B(n449), .Z(G1324GAT) );
  NOR2_X1 U505 ( .A1(n539), .A2(n454), .ZN(n450) );
  XOR2_X1 U506 ( .A(G8GAT), .B(n450), .Z(G1325GAT) );
  NOR2_X1 U507 ( .A1(n547), .A2(n454), .ZN(n452) );
  XNOR2_X1 U508 ( .A(KEYINPUT35), .B(KEYINPUT103), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U510 ( .A(G15GAT), .B(n453), .Z(G1326GAT) );
  NOR2_X1 U511 ( .A1(n510), .A2(n454), .ZN(n455) );
  XOR2_X1 U512 ( .A(KEYINPUT104), .B(n455), .Z(n456) );
  XNOR2_X1 U513 ( .A(G22GAT), .B(n456), .ZN(G1327GAT) );
  XNOR2_X1 U514 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n464) );
  XOR2_X1 U515 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n462) );
  NOR2_X1 U516 ( .A1(n457), .A2(n573), .ZN(n458) );
  XNOR2_X1 U517 ( .A(KEYINPUT36), .B(n558), .ZN(n576) );
  NAND2_X1 U518 ( .A1(n458), .A2(n576), .ZN(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT37), .B(n459), .ZN(n483) );
  NAND2_X1 U520 ( .A1(n460), .A2(n483), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(n470) );
  NOR2_X1 U522 ( .A1(n542), .A2(n470), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(G1328GAT) );
  NOR2_X1 U524 ( .A1(n539), .A2(n470), .ZN(n465) );
  XOR2_X1 U525 ( .A(KEYINPUT106), .B(n465), .Z(n466) );
  XNOR2_X1 U526 ( .A(G36GAT), .B(n466), .ZN(G1329GAT) );
  NOR2_X1 U527 ( .A1(n470), .A2(n547), .ZN(n468) );
  XNOR2_X1 U528 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n467) );
  XNOR2_X1 U529 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U530 ( .A(G43GAT), .B(n469), .ZN(G1330GAT) );
  NOR2_X1 U531 ( .A1(n470), .A2(n510), .ZN(n471) );
  XOR2_X1 U532 ( .A(G50GAT), .B(n471), .Z(G1331GAT) );
  XNOR2_X1 U533 ( .A(n569), .B(KEYINPUT41), .ZN(n529) );
  XOR2_X1 U534 ( .A(KEYINPUT108), .B(n529), .Z(n554) );
  AND2_X1 U535 ( .A1(n527), .A2(n554), .ZN(n482) );
  NAND2_X1 U536 ( .A1(n482), .A2(n472), .ZN(n478) );
  NOR2_X1 U537 ( .A1(n542), .A2(n478), .ZN(n473) );
  XOR2_X1 U538 ( .A(G57GAT), .B(n473), .Z(n474) );
  XNOR2_X1 U539 ( .A(KEYINPUT42), .B(n474), .ZN(G1332GAT) );
  NOR2_X1 U540 ( .A1(n539), .A2(n478), .ZN(n475) );
  XOR2_X1 U541 ( .A(G64GAT), .B(n475), .Z(G1333GAT) );
  NOR2_X1 U542 ( .A1(n547), .A2(n478), .ZN(n477) );
  XNOR2_X1 U543 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n476) );
  XNOR2_X1 U544 ( .A(n477), .B(n476), .ZN(G1334GAT) );
  NOR2_X1 U545 ( .A1(n510), .A2(n478), .ZN(n480) );
  XNOR2_X1 U546 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n479) );
  XNOR2_X1 U547 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U548 ( .A(G78GAT), .B(n481), .ZN(G1335GAT) );
  NAND2_X1 U549 ( .A1(n483), .A2(n482), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n542), .A2(n492), .ZN(n485) );
  XNOR2_X1 U551 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n484) );
  XNOR2_X1 U552 ( .A(n485), .B(n484), .ZN(G1336GAT) );
  NOR2_X1 U553 ( .A1(n539), .A2(n492), .ZN(n486) );
  XOR2_X1 U554 ( .A(KEYINPUT112), .B(n486), .Z(n487) );
  XNOR2_X1 U555 ( .A(G92GAT), .B(n487), .ZN(G1337GAT) );
  NOR2_X1 U556 ( .A1(n547), .A2(n492), .ZN(n489) );
  XNOR2_X1 U557 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n488) );
  XNOR2_X1 U558 ( .A(n489), .B(n488), .ZN(G1338GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n491) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n490) );
  XNOR2_X1 U561 ( .A(n491), .B(n490), .ZN(n494) );
  NOR2_X1 U562 ( .A1(n510), .A2(n492), .ZN(n493) );
  XOR2_X1 U563 ( .A(n494), .B(n493), .Z(G1339GAT) );
  INV_X1 U564 ( .A(n502), .ZN(n548) );
  NOR2_X1 U565 ( .A1(n527), .A2(n529), .ZN(n495) );
  XNOR2_X1 U566 ( .A(n495), .B(KEYINPUT46), .ZN(n496) );
  XNOR2_X1 U567 ( .A(n497), .B(KEYINPUT116), .ZN(n498) );
  NAND2_X1 U568 ( .A1(n498), .A2(n536), .ZN(n499) );
  XNOR2_X1 U569 ( .A(n499), .B(KEYINPUT47), .ZN(n506) );
  NAND2_X1 U570 ( .A1(n573), .A2(n576), .ZN(n501) );
  XNOR2_X1 U571 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n500) );
  XNOR2_X1 U572 ( .A(n501), .B(n500), .ZN(n503) );
  NAND2_X1 U573 ( .A1(n503), .A2(n502), .ZN(n504) );
  NOR2_X1 U574 ( .A1(n504), .A2(n569), .ZN(n505) );
  XNOR2_X1 U575 ( .A(n507), .B(KEYINPUT48), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n508), .B(KEYINPUT64), .ZN(n540) );
  NOR2_X1 U577 ( .A1(n540), .A2(n509), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n526), .A2(n510), .ZN(n511) );
  NOR2_X1 U579 ( .A1(n547), .A2(n511), .ZN(n520) );
  NAND2_X1 U580 ( .A1(n548), .A2(n520), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n512), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n514) );
  NAND2_X1 U583 ( .A1(n520), .A2(n554), .ZN(n513) );
  XNOR2_X1 U584 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U585 ( .A(G120GAT), .B(n515), .Z(G1341GAT) );
  XNOR2_X1 U586 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n519) );
  XOR2_X1 U587 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n517) );
  NAND2_X1 U588 ( .A1(n520), .A2(n573), .ZN(n516) );
  XNOR2_X1 U589 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U590 ( .A(n519), .B(n518), .ZN(G1342GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n522) );
  NAND2_X1 U592 ( .A1(n520), .A2(n558), .ZN(n521) );
  XNOR2_X1 U593 ( .A(n522), .B(n521), .ZN(n524) );
  XOR2_X1 U594 ( .A(G134GAT), .B(KEYINPUT120), .Z(n523) );
  XNOR2_X1 U595 ( .A(n524), .B(n523), .ZN(G1343GAT) );
  NAND2_X1 U596 ( .A1(n526), .A2(n525), .ZN(n535) );
  NOR2_X1 U597 ( .A1(n527), .A2(n535), .ZN(n528) );
  XOR2_X1 U598 ( .A(G141GAT), .B(n528), .Z(G1344GAT) );
  NOR2_X1 U599 ( .A1(n529), .A2(n535), .ZN(n531) );
  XNOR2_X1 U600 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n530) );
  XNOR2_X1 U601 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U602 ( .A(G148GAT), .B(n532), .ZN(G1345GAT) );
  INV_X1 U603 ( .A(n573), .ZN(n533) );
  NOR2_X1 U604 ( .A1(n533), .A2(n535), .ZN(n534) );
  XOR2_X1 U605 ( .A(G155GAT), .B(n534), .Z(G1346GAT) );
  NOR2_X1 U606 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U607 ( .A(KEYINPUT122), .B(n537), .Z(n538) );
  XNOR2_X1 U608 ( .A(G162GAT), .B(n538), .ZN(G1347GAT) );
  XOR2_X1 U609 ( .A(G169GAT), .B(KEYINPUT123), .Z(n550) );
  NOR2_X1 U610 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n541), .B(KEYINPUT54), .ZN(n543) );
  NAND2_X1 U612 ( .A1(n543), .A2(n542), .ZN(n563) );
  NOR2_X1 U613 ( .A1(n544), .A2(n563), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n545), .B(KEYINPUT55), .ZN(n546) );
  NAND2_X1 U615 ( .A1(n559), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n552) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(n553), .Z(n556) );
  NAND2_X1 U621 ( .A1(n559), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n573), .A2(n559), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(n562), .B(G190GAT), .Z(G1351GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n567) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n575), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n571) );
  NAND2_X1 U635 ( .A1(n575), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

