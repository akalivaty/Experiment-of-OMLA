

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  NOR2_X1 U322 ( .A1(n552), .A2(n551), .ZN(n563) );
  AND2_X1 U323 ( .A1(n546), .A2(n545), .ZN(n548) );
  AND2_X1 U324 ( .A1(n506), .A2(n579), .ZN(n290) );
  INV_X1 U325 ( .A(KEYINPUT64), .ZN(n547) );
  XNOR2_X1 U326 ( .A(n548), .B(n547), .ZN(n567) );
  XOR2_X1 U327 ( .A(n451), .B(n450), .Z(n569) );
  XOR2_X1 U328 ( .A(KEYINPUT102), .B(KEYINPUT34), .Z(n292) );
  XNOR2_X1 U329 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n291) );
  XNOR2_X1 U330 ( .A(n292), .B(n291), .ZN(n454) );
  XNOR2_X1 U331 ( .A(KEYINPUT91), .B(KEYINPUT2), .ZN(n293) );
  XNOR2_X1 U332 ( .A(n293), .B(G155GAT), .ZN(n294) );
  XOR2_X1 U333 ( .A(n294), .B(KEYINPUT92), .Z(n296) );
  XNOR2_X1 U334 ( .A(KEYINPUT3), .B(KEYINPUT93), .ZN(n295) );
  XNOR2_X1 U335 ( .A(n296), .B(n295), .ZN(n377) );
  XOR2_X1 U336 ( .A(G85GAT), .B(KEYINPUT1), .Z(n298) );
  XNOR2_X1 U337 ( .A(G162GAT), .B(KEYINPUT94), .ZN(n297) );
  XNOR2_X1 U338 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U339 ( .A(n377), .B(n299), .Z(n301) );
  NAND2_X1 U340 ( .A1(G225GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U341 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U342 ( .A(G148GAT), .B(G141GAT), .Z(n303) );
  XNOR2_X1 U343 ( .A(G29GAT), .B(G1GAT), .ZN(n302) );
  XNOR2_X1 U344 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U345 ( .A(n305), .B(n304), .Z(n314) );
  XNOR2_X1 U346 ( .A(G127GAT), .B(G134GAT), .ZN(n306) );
  XNOR2_X1 U347 ( .A(n306), .B(KEYINPUT83), .ZN(n307) );
  XOR2_X1 U348 ( .A(n307), .B(KEYINPUT0), .Z(n309) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(G120GAT), .ZN(n308) );
  XNOR2_X1 U350 ( .A(n309), .B(n308), .ZN(n368) );
  XOR2_X1 U351 ( .A(KEYINPUT6), .B(G57GAT), .Z(n311) );
  XNOR2_X1 U352 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n310) );
  XNOR2_X1 U353 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U354 ( .A(n368), .B(n312), .ZN(n313) );
  XNOR2_X1 U355 ( .A(n314), .B(n313), .ZN(n482) );
  XOR2_X1 U356 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n316) );
  XNOR2_X1 U357 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n315) );
  XNOR2_X1 U358 ( .A(n316), .B(n315), .ZN(n334) );
  XOR2_X1 U359 ( .A(G78GAT), .B(G211GAT), .Z(n318) );
  XNOR2_X1 U360 ( .A(G127GAT), .B(G183GAT), .ZN(n317) );
  XNOR2_X1 U361 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U362 ( .A(G64GAT), .B(G155GAT), .Z(n320) );
  XNOR2_X1 U363 ( .A(G22GAT), .B(G8GAT), .ZN(n319) );
  XNOR2_X1 U364 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U365 ( .A(n322), .B(n321), .Z(n332) );
  XOR2_X1 U366 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n324) );
  XNOR2_X1 U367 ( .A(G71GAT), .B(G57GAT), .ZN(n323) );
  XNOR2_X1 U368 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U369 ( .A(KEYINPUT72), .B(n325), .Z(n417) );
  XOR2_X1 U370 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n327) );
  XNOR2_X1 U371 ( .A(G15GAT), .B(G1GAT), .ZN(n326) );
  XNOR2_X1 U372 ( .A(n327), .B(n326), .ZN(n447) );
  XOR2_X1 U373 ( .A(n447), .B(KEYINPUT82), .Z(n329) );
  NAND2_X1 U374 ( .A1(G231GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U375 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U376 ( .A(n417), .B(n330), .ZN(n331) );
  XNOR2_X1 U377 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U378 ( .A(n334), .B(n333), .ZN(n560) );
  INV_X1 U379 ( .A(n560), .ZN(n579) );
  XOR2_X1 U380 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n336) );
  XNOR2_X1 U381 ( .A(KEYINPUT65), .B(KEYINPUT79), .ZN(n335) );
  XNOR2_X1 U382 ( .A(n336), .B(n335), .ZN(n353) );
  XOR2_X1 U383 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n338) );
  XNOR2_X1 U384 ( .A(G106GAT), .B(G92GAT), .ZN(n337) );
  XNOR2_X1 U385 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .Z(n394) );
  XOR2_X1 U387 ( .A(n339), .B(n394), .Z(n341) );
  XNOR2_X1 U388 ( .A(G134GAT), .B(G218GAT), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U390 ( .A(G99GAT), .B(G85GAT), .Z(n422) );
  XOR2_X1 U391 ( .A(n422), .B(KEYINPUT10), .Z(n343) );
  NAND2_X1 U392 ( .A1(G232GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U394 ( .A(n345), .B(n344), .Z(n351) );
  XOR2_X1 U395 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n347) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(G29GAT), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U398 ( .A(KEYINPUT7), .B(n348), .ZN(n450) );
  INV_X1 U399 ( .A(n450), .ZN(n349) );
  XOR2_X1 U400 ( .A(G50GAT), .B(G162GAT), .Z(n373) );
  XNOR2_X1 U401 ( .A(n349), .B(n373), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U403 ( .A(n353), .B(n352), .Z(n539) );
  INV_X1 U404 ( .A(n539), .ZN(n562) );
  NOR2_X1 U405 ( .A1(n579), .A2(n562), .ZN(n354) );
  XNOR2_X1 U406 ( .A(KEYINPUT16), .B(n354), .ZN(n415) );
  XOR2_X1 U407 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n356) );
  XNOR2_X1 U408 ( .A(KEYINPUT85), .B(KEYINPUT88), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n372) );
  XOR2_X1 U410 ( .A(G71GAT), .B(G190GAT), .Z(n358) );
  XNOR2_X1 U411 ( .A(G43GAT), .B(G99GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U413 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n360) );
  XNOR2_X1 U414 ( .A(G15GAT), .B(G176GAT), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U416 ( .A(n362), .B(n361), .Z(n370) );
  XOR2_X1 U417 ( .A(G183GAT), .B(KEYINPUT18), .Z(n364) );
  XNOR2_X1 U418 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n391) );
  XOR2_X1 U420 ( .A(G169GAT), .B(n391), .Z(n366) );
  NAND2_X1 U421 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n552) );
  XOR2_X1 U426 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n375) );
  XOR2_X1 U427 ( .A(G141GAT), .B(G22GAT), .Z(n434) );
  XNOR2_X1 U428 ( .A(n434), .B(n373), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U430 ( .A(n377), .B(n376), .Z(n379) );
  NAND2_X1 U431 ( .A1(G228GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U433 ( .A(G204GAT), .B(KEYINPUT24), .Z(n381) );
  XNOR2_X1 U434 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U436 ( .A(n383), .B(n382), .Z(n389) );
  XOR2_X1 U437 ( .A(G211GAT), .B(KEYINPUT21), .Z(n385) );
  XNOR2_X1 U438 ( .A(G197GAT), .B(G218GAT), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n396) );
  XOR2_X1 U440 ( .A(G78GAT), .B(G148GAT), .Z(n387) );
  XNOR2_X1 U441 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n426) );
  XNOR2_X1 U443 ( .A(n396), .B(n426), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n549) );
  XNOR2_X1 U445 ( .A(n549), .B(KEYINPUT66), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n390), .B(KEYINPUT28), .ZN(n489) );
  INV_X1 U447 ( .A(n482), .ZN(n545) );
  XOR2_X1 U448 ( .A(KEYINPUT95), .B(n391), .Z(n393) );
  NAND2_X1 U449 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U451 ( .A(n395), .B(n394), .Z(n398) );
  XOR2_X1 U452 ( .A(G169GAT), .B(G8GAT), .Z(n435) );
  XNOR2_X1 U453 ( .A(n435), .B(n396), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U455 ( .A(G92GAT), .B(G64GAT), .Z(n400) );
  XNOR2_X1 U456 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U458 ( .A(G204GAT), .B(n401), .Z(n418) );
  XNOR2_X1 U459 ( .A(n402), .B(n418), .ZN(n485) );
  INV_X1 U460 ( .A(n485), .ZN(n543) );
  XNOR2_X1 U461 ( .A(n543), .B(KEYINPUT27), .ZN(n407) );
  OR2_X1 U462 ( .A1(n545), .A2(n407), .ZN(n528) );
  NOR2_X1 U463 ( .A1(n489), .A2(n528), .ZN(n514) );
  NAND2_X1 U464 ( .A1(n552), .A2(n514), .ZN(n413) );
  NOR2_X1 U465 ( .A1(n543), .A2(n552), .ZN(n403) );
  NOR2_X1 U466 ( .A1(n549), .A2(n403), .ZN(n404) );
  XOR2_X1 U467 ( .A(n404), .B(KEYINPUT96), .Z(n405) );
  XNOR2_X1 U468 ( .A(KEYINPUT25), .B(n405), .ZN(n409) );
  NAND2_X1 U469 ( .A1(n552), .A2(n549), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n406), .B(KEYINPUT26), .ZN(n566) );
  NOR2_X1 U471 ( .A1(n566), .A2(n407), .ZN(n408) );
  NOR2_X1 U472 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n410), .B(KEYINPUT97), .ZN(n411) );
  NAND2_X1 U474 ( .A1(n411), .A2(n545), .ZN(n412) );
  NAND2_X1 U475 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n414), .B(KEYINPUT98), .ZN(n465) );
  NAND2_X1 U477 ( .A1(n415), .A2(n465), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n416), .B(KEYINPUT99), .ZN(n480) );
  XOR2_X1 U479 ( .A(n418), .B(n417), .Z(n430) );
  XOR2_X1 U480 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n420) );
  XNOR2_X1 U481 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U483 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U484 ( .A1(G230GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U486 ( .A(n425), .B(KEYINPUT33), .Z(n428) );
  XNOR2_X1 U487 ( .A(n426), .B(KEYINPUT76), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n574) );
  XOR2_X1 U490 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n432) );
  XNOR2_X1 U491 ( .A(G113GAT), .B(G197GAT), .ZN(n431) );
  XOR2_X1 U492 ( .A(n432), .B(n431), .Z(n438) );
  XOR2_X1 U493 ( .A(G36GAT), .B(G50GAT), .Z(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n442) );
  INV_X1 U497 ( .A(n442), .ZN(n440) );
  NAND2_X1 U498 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  INV_X1 U499 ( .A(n441), .ZN(n439) );
  NAND2_X1 U500 ( .A1(n440), .A2(n439), .ZN(n444) );
  NAND2_X1 U501 ( .A1(n442), .A2(n441), .ZN(n443) );
  NAND2_X1 U502 ( .A1(n444), .A2(n443), .ZN(n446) );
  INV_X1 U503 ( .A(KEYINPUT30), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n447), .B(KEYINPUT67), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n451) );
  INV_X1 U507 ( .A(n569), .ZN(n553) );
  AND2_X1 U508 ( .A1(n574), .A2(n553), .ZN(n467) );
  NAND2_X1 U509 ( .A1(n480), .A2(n467), .ZN(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT100), .B(n452), .Z(n462) );
  NAND2_X1 U511 ( .A1(n482), .A2(n462), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(G1324GAT) );
  XOR2_X1 U513 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n456) );
  NAND2_X1 U514 ( .A1(n462), .A2(n485), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U516 ( .A(G8GAT), .B(n457), .ZN(G1325GAT) );
  XOR2_X1 U517 ( .A(G15GAT), .B(KEYINPUT106), .Z(n459) );
  INV_X1 U518 ( .A(n552), .ZN(n515) );
  NAND2_X1 U519 ( .A1(n515), .A2(n462), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n460) );
  XNOR2_X1 U522 ( .A(n461), .B(n460), .ZN(G1326GAT) );
  NAND2_X1 U523 ( .A1(n462), .A2(n489), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U525 ( .A(KEYINPUT107), .B(KEYINPUT38), .Z(n469) );
  XNOR2_X1 U526 ( .A(n539), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U527 ( .A1(n583), .A2(n560), .ZN(n464) );
  NAND2_X1 U528 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U529 ( .A(KEYINPUT37), .B(n466), .ZN(n494) );
  NAND2_X1 U530 ( .A1(n494), .A2(n467), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n469), .B(n468), .ZN(n477) );
  NOR2_X1 U532 ( .A1(n477), .A2(n545), .ZN(n471) );
  XNOR2_X1 U533 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n471), .B(n470), .ZN(G1328GAT) );
  NOR2_X1 U535 ( .A1(n543), .A2(n477), .ZN(n472) );
  XOR2_X1 U536 ( .A(G36GAT), .B(n472), .Z(G1329GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n474) );
  XNOR2_X1 U538 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n473) );
  XNOR2_X1 U539 ( .A(n474), .B(n473), .ZN(n476) );
  NOR2_X1 U540 ( .A1(n477), .A2(n552), .ZN(n475) );
  XOR2_X1 U541 ( .A(n476), .B(n475), .Z(G1330GAT) );
  INV_X1 U542 ( .A(n489), .ZN(n501) );
  NOR2_X1 U543 ( .A1(n477), .A2(n501), .ZN(n478) );
  XOR2_X1 U544 ( .A(G50GAT), .B(n478), .Z(G1331GAT) );
  INV_X1 U545 ( .A(KEYINPUT41), .ZN(n479) );
  XNOR2_X1 U546 ( .A(n574), .B(n479), .ZN(n532) );
  XOR2_X1 U547 ( .A(KEYINPUT110), .B(n532), .Z(n555) );
  AND2_X1 U548 ( .A1(n569), .A2(n555), .ZN(n493) );
  NAND2_X1 U549 ( .A1(n493), .A2(n480), .ZN(n481) );
  XNOR2_X1 U550 ( .A(n481), .B(KEYINPUT111), .ZN(n490) );
  NAND2_X1 U551 ( .A1(n490), .A2(n482), .ZN(n483) );
  XNOR2_X1 U552 ( .A(n483), .B(KEYINPUT42), .ZN(n484) );
  XNOR2_X1 U553 ( .A(G57GAT), .B(n484), .ZN(G1332GAT) );
  NAND2_X1 U554 ( .A1(n485), .A2(n490), .ZN(n486) );
  XNOR2_X1 U555 ( .A(n486), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U556 ( .A1(n490), .A2(n515), .ZN(n487) );
  XNOR2_X1 U557 ( .A(n487), .B(KEYINPUT112), .ZN(n488) );
  XNOR2_X1 U558 ( .A(G71GAT), .B(n488), .ZN(G1334GAT) );
  XOR2_X1 U559 ( .A(G78GAT), .B(KEYINPUT43), .Z(n492) );
  NAND2_X1 U560 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U561 ( .A(n492), .B(n491), .ZN(G1335GAT) );
  NAND2_X1 U562 ( .A1(n494), .A2(n493), .ZN(n500) );
  NOR2_X1 U563 ( .A1(n545), .A2(n500), .ZN(n496) );
  XNOR2_X1 U564 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n495) );
  XNOR2_X1 U565 ( .A(n496), .B(n495), .ZN(G1336GAT) );
  NOR2_X1 U566 ( .A1(n543), .A2(n500), .ZN(n497) );
  XOR2_X1 U567 ( .A(G92GAT), .B(n497), .Z(G1337GAT) );
  NOR2_X1 U568 ( .A1(n552), .A2(n500), .ZN(n498) );
  XOR2_X1 U569 ( .A(KEYINPUT114), .B(n498), .Z(n499) );
  XNOR2_X1 U570 ( .A(G99GAT), .B(n499), .ZN(G1338GAT) );
  NOR2_X1 U571 ( .A1(n501), .A2(n500), .ZN(n502) );
  XOR2_X1 U572 ( .A(KEYINPUT44), .B(n502), .Z(n503) );
  XNOR2_X1 U573 ( .A(G106GAT), .B(n503), .ZN(G1339GAT) );
  NOR2_X1 U574 ( .A1(n569), .A2(n532), .ZN(n505) );
  XNOR2_X1 U575 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n504) );
  XNOR2_X1 U576 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U577 ( .A1(n539), .A2(n290), .ZN(n507) );
  XNOR2_X1 U578 ( .A(n507), .B(KEYINPUT47), .ZN(n512) );
  NOR2_X1 U579 ( .A1(n579), .A2(n583), .ZN(n508) );
  XNOR2_X1 U580 ( .A(n508), .B(KEYINPUT45), .ZN(n509) );
  NAND2_X1 U581 ( .A1(n509), .A2(n574), .ZN(n510) );
  NOR2_X1 U582 ( .A1(n510), .A2(n553), .ZN(n511) );
  NOR2_X1 U583 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U584 ( .A(n513), .B(KEYINPUT48), .ZN(n542) );
  NAND2_X1 U585 ( .A1(n515), .A2(n514), .ZN(n516) );
  NOR2_X1 U586 ( .A1(n542), .A2(n516), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n524), .A2(n553), .ZN(n517) );
  XNOR2_X1 U588 ( .A(n517), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n519) );
  NAND2_X1 U590 ( .A1(n524), .A2(n555), .ZN(n518) );
  XNOR2_X1 U591 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U592 ( .A(G120GAT), .B(n520), .ZN(G1341GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n522) );
  NAND2_X1 U594 ( .A1(n524), .A2(n560), .ZN(n521) );
  XNOR2_X1 U595 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n523), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n526) );
  NAND2_X1 U598 ( .A1(n524), .A2(n562), .ZN(n525) );
  XNOR2_X1 U599 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U600 ( .A(G134GAT), .B(n527), .ZN(G1343GAT) );
  INV_X1 U601 ( .A(n542), .ZN(n530) );
  NOR2_X1 U602 ( .A1(n566), .A2(n528), .ZN(n529) );
  NAND2_X1 U603 ( .A1(n530), .A2(n529), .ZN(n538) );
  NOR2_X1 U604 ( .A1(n569), .A2(n538), .ZN(n531) );
  XOR2_X1 U605 ( .A(G141GAT), .B(n531), .Z(G1344GAT) );
  NOR2_X1 U606 ( .A1(n538), .A2(n532), .ZN(n536) );
  XOR2_X1 U607 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n534) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n533) );
  XNOR2_X1 U609 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U610 ( .A(n536), .B(n535), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n579), .A2(n538), .ZN(n537) );
  XOR2_X1 U612 ( .A(G155GAT), .B(n537), .Z(G1346GAT) );
  NOR2_X1 U613 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U614 ( .A(KEYINPUT120), .B(n540), .Z(n541) );
  XNOR2_X1 U615 ( .A(G162GAT), .B(n541), .ZN(G1347GAT) );
  NOR2_X1 U616 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U617 ( .A(KEYINPUT54), .B(n544), .ZN(n546) );
  NOR2_X1 U618 ( .A1(n549), .A2(n567), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n550), .B(KEYINPUT55), .ZN(n551) );
  NAND2_X1 U620 ( .A1(n563), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT57), .Z(n557) );
  NAND2_X1 U623 ( .A1(n563), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n563), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT122), .B(n568), .Z(n584) );
  NOR2_X1 U634 ( .A1(n569), .A2(n584), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n584), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n584), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n582) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n586), .B(n585), .Z(G1355GAT) );
endmodule

