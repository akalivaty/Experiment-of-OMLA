//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n203), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n202), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  INV_X1    g0027(.A(new_n206), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n219), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(G20), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n212), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n227), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n216), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n219), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n202), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n215), .ZN(new_n251));
  INV_X1    g0051(.A(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  OAI21_X1  g0054(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G150), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OR3_X1    g0060(.A1(new_n259), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n255), .A2(new_n257), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n230), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n209), .B2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n219), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n268), .A2(KEYINPUT9), .A3(new_n270), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT72), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n265), .A2(new_n267), .B1(new_n219), .B2(new_n272), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT72), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT9), .A4(new_n270), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n262), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G223), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT67), .B(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G222), .ZN(new_n287));
  OAI221_X1 g0087(.A(new_n283), .B1(new_n284), .B2(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n289), .C1(G77), .C2(new_n283), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n289), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n295), .A2(new_n291), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G226), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n290), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G190), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n276), .A2(new_n270), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n301), .A2(new_n302), .B1(G200), .B2(new_n298), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n279), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT73), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n309), .A2(new_n279), .A3(new_n300), .A4(new_n303), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n299), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n298), .A2(new_n314), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n313), .A2(new_n315), .A3(new_n301), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n258), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n320));
  INV_X1    g0120(.A(new_n263), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n323), .A2(new_n267), .B1(new_n221), .B2(new_n272), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n269), .A2(G77), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(KEYINPUT69), .A2(G107), .ZN(new_n327));
  NOR2_X1   g0127(.A1(KEYINPUT69), .A2(G107), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n283), .B1(new_n214), .B2(new_n285), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n286), .A2(new_n224), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n289), .B1(new_n283), .B2(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n296), .A2(G244), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n294), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n314), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n326), .B(new_n335), .C1(G179), .C2(new_n334), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(G200), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT70), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n337), .B1(new_n338), .B2(new_n334), .C1(new_n326), .C2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT70), .B1(new_n324), .B2(new_n325), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT71), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G97), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT67), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT3), .A2(G33), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n344), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n293), .B1(new_n353), .B2(new_n289), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n296), .A2(G238), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n355), .B1(new_n354), .B2(new_n356), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT14), .B1(new_n360), .B2(new_n314), .ZN(new_n361));
  INV_X1    g0161(.A(new_n359), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n357), .A3(G179), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(G169), .C1(new_n358), .C2(new_n359), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n256), .A2(G50), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT74), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n321), .A2(new_n221), .B1(new_n210), .B2(G68), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n267), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XOR2_X1   g0170(.A(new_n370), .B(KEYINPUT11), .Z(new_n371));
  NAND4_X1  g0171(.A1(new_n209), .A2(new_n203), .A3(G13), .A4(G20), .ZN(new_n372));
  XOR2_X1   g0172(.A(new_n372), .B(KEYINPUT12), .Z(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(G68), .B2(new_n269), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n366), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n362), .A2(new_n357), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G200), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n376), .C1(new_n338), .C2(new_n379), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n260), .A2(new_n261), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n269), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n383), .B2(new_n271), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT76), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n352), .B2(new_n210), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n282), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n204), .A2(new_n205), .A3(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(G20), .B1(G159), .B2(new_n256), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n386), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI211_X1 g0196(.A(KEYINPUT76), .B(KEYINPUT16), .C1(new_n390), .C2(new_n393), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n281), .A2(new_n210), .A3(new_n282), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(KEYINPUT75), .A3(new_n388), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n388), .A2(KEYINPUT75), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(G68), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n393), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n405), .A2(new_n267), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n385), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n296), .A2(G232), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n286), .A2(new_n284), .B1(new_n220), .B2(new_n285), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(new_n283), .B1(G33), .B2(G87), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n294), .C1(new_n410), .C2(new_n295), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G200), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n411), .A2(new_n338), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n203), .B1(new_n401), .B2(new_n388), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n392), .A2(G20), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n256), .A2(G159), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n395), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT76), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n386), .B(new_n395), .C1(new_n415), .C2(new_n418), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n420), .A2(new_n267), .A3(new_n405), .A4(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n385), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n422), .A2(new_n413), .A3(new_n412), .A4(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n411), .A2(G169), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n348), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n429));
  INV_X1    g0229(.A(G87), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n429), .A2(new_n352), .B1(new_n262), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n289), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n432), .A2(G179), .A3(new_n408), .A4(new_n294), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT18), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  AOI221_X4 g0236(.A(new_n436), .B1(new_n428), .B2(new_n433), .C1(new_n422), .C2(new_n423), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n414), .B(new_n426), .C1(new_n435), .C2(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n318), .A2(new_n343), .A3(new_n382), .A4(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(G116), .B2(new_n263), .ZN(new_n441));
  OAI21_X1  g0241(.A(G20), .B1(new_n327), .B2(new_n328), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT81), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT23), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n442), .B2(KEYINPUT23), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n210), .B(G87), .C1(new_n350), .C2(new_n351), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT22), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n447), .B(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT24), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n442), .A2(KEYINPUT23), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT23), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n447), .B(KEYINPUT22), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT24), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .A4(new_n441), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n450), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n267), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n209), .A2(G33), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n271), .A2(new_n460), .A3(new_n230), .A4(new_n266), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n215), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n272), .A2(new_n215), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n464), .B(KEYINPUT25), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(G274), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n289), .B1(new_n470), .B2(new_n468), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G264), .ZN(new_n473));
  INV_X1    g0273(.A(G250), .ZN(new_n474));
  INV_X1    g0274(.A(G257), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n286), .A2(new_n474), .B1(new_n475), .B2(new_n285), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(new_n283), .B1(G33), .B2(G294), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n471), .B(new_n473), .C1(new_n477), .C2(new_n295), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n314), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(G179), .B2(new_n478), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n467), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n210), .C1(G33), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n252), .A2(G20), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n267), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT80), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(KEYINPUT80), .A2(KEYINPUT20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n489), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n485), .A2(new_n267), .A3(new_n492), .A4(new_n486), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n271), .A2(new_n252), .ZN(new_n495));
  INV_X1    g0295(.A(new_n461), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n252), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n314), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI221_X1 g0298(.A(new_n283), .B1(new_n216), .B2(new_n285), .C1(new_n286), .C2(new_n475), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n499), .B(new_n289), .C1(G303), .C2(new_n283), .ZN(new_n500));
  INV_X1    g0300(.A(new_n471), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(G270), .B2(new_n472), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(KEYINPUT21), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT21), .B1(new_n498), .B2(new_n503), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n494), .A2(new_n497), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(new_n502), .A3(G179), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n505), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n503), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n507), .B1(new_n512), .B2(G190), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n306), .B2(new_n512), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n482), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT19), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n210), .B1(new_n344), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT77), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n430), .B(new_n484), .C1(new_n327), .C2(new_n328), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT77), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n210), .C1(new_n344), .C2(new_n516), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT78), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT19), .B1(new_n263), .B2(G97), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n352), .A2(G20), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G68), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT78), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n518), .A2(new_n519), .A3(new_n527), .A4(new_n521), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n523), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n523), .A2(new_n526), .A3(KEYINPUT79), .A4(new_n528), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n267), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n322), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n496), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n322), .A2(new_n272), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n289), .B1(new_n292), .B2(new_n470), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(G250), .B2(new_n470), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n286), .A2(new_n214), .B1(new_n222), .B2(new_n285), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n283), .B1(G33), .B2(G116), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(new_n295), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(G179), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n314), .B2(new_n542), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n306), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G190), .B2(new_n542), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n496), .A2(G87), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n547), .A2(new_n533), .A3(new_n536), .A4(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n283), .A2(new_n348), .A3(G244), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT4), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n283), .A2(new_n348), .A3(KEYINPUT4), .A4(G244), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n285), .B1(new_n281), .B2(new_n282), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n289), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n475), .B(new_n289), .C1(new_n470), .C2(new_n468), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n557), .A2(new_n312), .A3(new_n471), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n256), .A2(G77), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT6), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n562), .A2(new_n484), .A3(G107), .ZN(new_n563));
  XNOR2_X1  g0363(.A(G97), .B(G107), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n561), .B1(new_n565), .B2(new_n210), .ZN(new_n566));
  INV_X1    g0366(.A(new_n329), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n401), .B2(new_n388), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n267), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n496), .A2(G97), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n272), .A2(new_n484), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n501), .B(new_n558), .C1(new_n556), .C2(new_n289), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n560), .B(new_n572), .C1(new_n573), .C2(G169), .ZN(new_n574));
  INV_X1    g0374(.A(new_n572), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n557), .A2(G190), .A3(new_n471), .A4(new_n559), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n306), .C2(new_n573), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n545), .A2(new_n549), .A3(new_n574), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n462), .B1(new_n458), .B2(new_n267), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n478), .A2(G200), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n478), .A2(new_n338), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n580), .A2(new_n466), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  AND4_X1   g0383(.A1(new_n439), .A2(new_n515), .A3(new_n579), .A4(new_n583), .ZN(G372));
  NAND2_X1  g0384(.A1(new_n378), .A2(new_n336), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n585), .A2(new_n426), .A3(new_n414), .A4(new_n381), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n435), .B2(new_n437), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n316), .B1(new_n587), .B2(new_n311), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n533), .A2(new_n536), .A3(new_n548), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(new_n547), .B1(new_n537), .B2(new_n544), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n574), .A2(KEYINPUT82), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n557), .A2(new_n471), .A3(new_n559), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n314), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(new_n572), .A4(new_n560), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT26), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n590), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n574), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n545), .A2(new_n599), .A3(new_n549), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT26), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n480), .B1(new_n580), .B2(new_n466), .ZN(new_n603));
  INV_X1    g0403(.A(new_n510), .ZN(new_n604));
  INV_X1    g0404(.A(new_n506), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n504), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n583), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n545), .B1(new_n607), .B2(new_n578), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n439), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n588), .A2(new_n610), .ZN(G369));
  NAND3_X1  g0411(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(G213), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G343), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n603), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n467), .A2(new_n617), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n603), .B1(new_n620), .B2(new_n583), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n606), .A2(new_n618), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT83), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(KEYINPUT83), .B(new_n619), .C1(new_n621), .C2(new_n622), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n606), .B1(new_n508), .B2(new_n618), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n511), .A2(new_n507), .A3(new_n617), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n514), .ZN(new_n630));
  INV_X1    g0430(.A(G330), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n619), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n621), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n622), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n627), .A2(new_n636), .ZN(G399));
  INV_X1    g0437(.A(new_n233), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(G41), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n229), .ZN(new_n640));
  INV_X1    g0440(.A(new_n639), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G1), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n519), .A2(G116), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT28), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n473), .B1(new_n477), .B2(new_n295), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n542), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(G179), .A3(new_n512), .A4(new_n573), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT30), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n573), .A2(new_n512), .A3(G179), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n478), .A3(new_n542), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n617), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT31), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n515), .A2(new_n579), .A3(new_n583), .A4(new_n618), .ZN(new_n658));
  XNOR2_X1  g0458(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n657), .B(new_n658), .C1(new_n655), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT29), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n609), .A2(new_n663), .A3(new_n618), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n590), .A2(new_n596), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n666));
  AOI211_X1 g0466(.A(new_n462), .B(new_n465), .C1(new_n458), .C2(new_n267), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n511), .B1(new_n667), .B2(new_n480), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n577), .A2(new_n574), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n590), .A3(new_n669), .A4(new_n583), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n590), .A2(new_n597), .A3(new_n599), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n666), .A2(new_n670), .A3(new_n545), .A4(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n672), .A2(new_n618), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n662), .B(new_n664), .C1(new_n663), .C2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n645), .B1(new_n675), .B2(G1), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT85), .ZN(G364));
  INV_X1    g0477(.A(G13), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G20), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n642), .B1(G45), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n632), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n630), .A2(new_n631), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n230), .B1(G20), .B2(new_n314), .ZN(new_n684));
  NOR3_X1   g0484(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n249), .A2(G45), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n638), .A2(new_n283), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n229), .B2(new_n469), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n686), .A2(new_n689), .B1(new_n252), .B2(new_n638), .ZN(new_n690));
  XOR2_X1   g0490(.A(G355), .B(KEYINPUT86), .Z(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n233), .A3(new_n283), .ZN(new_n692));
  AOI211_X1 g0492(.A(new_n684), .B(new_n685), .C1(new_n690), .C2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n680), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n685), .B(KEYINPUT89), .Z(new_n695));
  AOI211_X1 g0495(.A(new_n693), .B(new_n694), .C1(new_n630), .C2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n210), .A2(new_n312), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(G190), .A3(G200), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR4_X1   g0499(.A1(new_n210), .A2(new_n312), .A3(new_n338), .A4(G200), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n699), .A2(G50), .B1(new_n700), .B2(G58), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n338), .A2(G20), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT87), .ZN(new_n703));
  NOR2_X1   g0503(.A1(G179), .A2(G200), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G159), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n283), .B(new_n701), .C1(new_n707), .C2(KEYINPUT32), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n704), .A2(G190), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G20), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n707), .A2(KEYINPUT32), .B1(G97), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n306), .A2(G179), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT88), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(G20), .A3(G190), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G87), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n713), .A2(new_n703), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G107), .ZN(new_n718));
  NOR4_X1   g0518(.A1(new_n210), .A2(new_n312), .A3(new_n306), .A4(G190), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G68), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n711), .A2(new_n716), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n697), .A2(new_n338), .A3(new_n306), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI211_X1 g0523(.A(new_n708), .B(new_n721), .C1(G77), .C2(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n706), .A2(G329), .B1(G294), .B2(new_n710), .ZN(new_n725));
  INV_X1    g0525(.A(G311), .ZN(new_n726));
  INV_X1    g0526(.A(G322), .ZN(new_n727));
  INV_X1    g0527(.A(new_n700), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n725), .B1(new_n726), .B2(new_n722), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n719), .ZN(new_n730));
  INV_X1    g0530(.A(G317), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n730), .B1(KEYINPUT33), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(KEYINPUT33), .B2(new_n731), .ZN(new_n733));
  INV_X1    g0533(.A(G283), .ZN(new_n734));
  INV_X1    g0534(.A(new_n717), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n733), .B(new_n352), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G326), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n698), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G303), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n714), .A2(new_n739), .ZN(new_n740));
  NOR4_X1   g0540(.A1(new_n729), .A2(new_n736), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n684), .B1(new_n724), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n696), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n683), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(G396));
  NAND2_X1  g0545(.A1(new_n609), .A2(new_n618), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n336), .A2(new_n617), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n326), .A2(new_n617), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n340), .B2(new_n341), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(new_n749), .B2(new_n336), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n618), .B(new_n750), .C1(new_n602), .C2(new_n608), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n662), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n694), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G143), .A2(new_n700), .B1(new_n719), .B2(G150), .ZN(new_n758));
  INV_X1    g0558(.A(G137), .ZN(new_n759));
  INV_X1    g0559(.A(G159), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n758), .B1(new_n759), .B2(new_n698), .C1(new_n760), .C2(new_n722), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT90), .Z(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT34), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n735), .A2(new_n203), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n714), .A2(new_n219), .ZN(new_n765));
  INV_X1    g0565(.A(new_n710), .ZN(new_n766));
  INV_X1    g0566(.A(G132), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n283), .B1(new_n766), .B2(new_n202), .C1(new_n705), .C2(new_n767), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n763), .A2(new_n764), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n715), .A2(G107), .B1(G283), .B2(new_n719), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n430), .B2(new_n735), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n699), .A2(G303), .B1(G97), .B2(new_n710), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n772), .B(new_n352), .C1(new_n252), .C2(new_n722), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n705), .A2(new_n726), .ZN(new_n774));
  INV_X1    g0574(.A(G294), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n728), .A2(new_n775), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n771), .A2(new_n773), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n684), .B1(new_n769), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n684), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n221), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n751), .A2(new_n779), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n778), .A2(new_n680), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n757), .A2(new_n783), .ZN(G384));
  INV_X1    g0584(.A(new_n615), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n438), .A2(new_n427), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT95), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n428), .A2(new_n433), .A3(new_n615), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n424), .B1(new_n407), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT37), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT37), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n424), .B(new_n792), .C1(new_n407), .C2(new_n789), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT95), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n438), .A2(new_n795), .A3(new_n427), .A4(new_n785), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n787), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT38), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n405), .A2(new_n267), .ZN(new_n800));
  AOI21_X1  g0600(.A(KEYINPUT16), .B1(new_n404), .B2(new_n393), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n423), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n438), .A2(new_n785), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n788), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n424), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(KEYINPUT37), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT93), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n806), .A2(KEYINPUT93), .A3(new_n793), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n803), .A2(new_n807), .A3(KEYINPUT38), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n799), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT39), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n366), .A2(new_n377), .A3(new_n618), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT94), .Z(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n803), .A2(new_n807), .A3(new_n808), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n798), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(KEYINPUT39), .A3(new_n809), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n812), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT91), .ZN(new_n820));
  INV_X1    g0620(.A(new_n747), .ZN(new_n821));
  AND3_X1   g0621(.A1(new_n753), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n820), .B1(new_n753), .B2(new_n821), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n365), .A2(new_n363), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n364), .B1(new_n379), .B2(G169), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n377), .B(new_n617), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT92), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n366), .A2(KEYINPUT92), .A3(new_n377), .A4(new_n617), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n381), .B(new_n378), .C1(new_n376), .C2(new_n618), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n817), .A2(new_n809), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n824), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n437), .A2(new_n435), .A3(new_n785), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n819), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n664), .B1(new_n673), .B2(new_n663), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n439), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(new_n588), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n837), .B(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n809), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n798), .B2(new_n797), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n751), .B1(new_n831), .B2(new_n832), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n654), .A2(new_n656), .A3(new_n617), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n658), .A2(new_n655), .A3(new_n659), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT40), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n833), .A2(new_n750), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n845), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(new_n834), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n631), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n439), .A2(G330), .A3(new_n845), .A4(new_n846), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n848), .A2(new_n853), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n439), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n857), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n841), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n209), .B2(new_n679), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT35), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n210), .B(new_n230), .C1(new_n565), .C2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n864), .B(G116), .C1(new_n863), .C2(new_n565), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT36), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n229), .A2(G77), .A3(new_n391), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(G50), .B2(new_n203), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(G1), .A3(new_n678), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n862), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT96), .Z(G367));
  NOR2_X1   g0671(.A1(new_n684), .A2(new_n685), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n872), .B1(new_n233), .B2(new_n322), .C1(new_n245), .C2(new_n688), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n680), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT101), .Z(new_n875));
  INV_X1    g0675(.A(new_n695), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n533), .A2(new_n536), .A3(new_n548), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n617), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n537), .B2(new_n544), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT97), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n545), .A2(new_n549), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n878), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n881), .B1(new_n880), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n766), .A2(new_n203), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(G50), .B2(new_n723), .ZN(new_n888));
  INV_X1    g0688(.A(G150), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n728), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n735), .A2(new_n221), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n759), .B2(new_n705), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n352), .B(new_n893), .C1(G143), .C2(new_n699), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n894), .B1(new_n202), .B2(new_n714), .C1(new_n760), .C2(new_n730), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n715), .A2(G116), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT46), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n766), .A2(new_n567), .B1(new_n722), .B2(new_n734), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT102), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(G97), .B2(new_n717), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n283), .B1(new_n706), .B2(G317), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n719), .A2(G294), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n897), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n728), .A2(new_n739), .B1(new_n698), .B2(new_n726), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT103), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n895), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT47), .Z(new_n907));
  INV_X1    g0707(.A(new_n684), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n875), .B1(new_n876), .B2(new_n886), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n620), .A2(new_n583), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(new_n606), .A3(new_n482), .A4(new_n618), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n572), .A2(new_n617), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n669), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT42), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT42), .ZN(new_n915));
  INV_X1    g0715(.A(new_n913), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n634), .A2(new_n915), .A3(new_n635), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n633), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n599), .A2(new_n618), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n914), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT98), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT43), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n884), .B2(new_n885), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT98), .B1(new_n920), .B2(new_n924), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT99), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n920), .A2(new_n930), .A3(new_n924), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n929), .B1(new_n928), .B2(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n599), .A2(new_n617), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n913), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n933), .A2(new_n934), .B1(new_n636), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n927), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n920), .A2(KEYINPUT98), .A3(new_n924), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n931), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT99), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n636), .A2(new_n937), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n943), .A3(new_n932), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n209), .B1(new_n679), .B2(G45), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n937), .B1(new_n625), .B2(new_n626), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT45), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n625), .A2(new_n626), .A3(new_n937), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT44), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n636), .A3(new_n952), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n622), .B1(new_n621), .B2(new_n633), .C1(new_n630), .C2(new_n631), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n636), .A2(new_n954), .A3(new_n911), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n674), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n956), .A3(KEYINPUT100), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n675), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n639), .B(KEYINPUT41), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n947), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n909), .B1(new_n945), .B2(new_n960), .ZN(G387));
  OR2_X1    g0761(.A1(new_n673), .A2(new_n663), .ZN(new_n962));
  INV_X1    g0762(.A(new_n955), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n962), .A2(new_n664), .A3(new_n662), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n674), .A2(new_n955), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n965), .A3(new_n639), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G311), .A2(new_n719), .B1(new_n700), .B2(G317), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n739), .B2(new_n722), .C1(new_n727), .C2(new_n698), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT48), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n734), .B2(new_n766), .C1(new_n775), .C2(new_n714), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT49), .Z(new_n971));
  OAI221_X1 g0771(.A(new_n352), .B1(new_n737), .B2(new_n705), .C1(new_n735), .C2(new_n252), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n383), .A2(new_n730), .B1(new_n203), .B2(new_n722), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT105), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n715), .A2(G77), .B1(new_n706), .B2(G150), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(new_n484), .C2(new_n735), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n283), .B1(new_n766), .B2(new_n322), .C1(new_n728), .C2(new_n219), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n698), .A2(new_n760), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT104), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n684), .B1(new_n973), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n695), .B1(new_n621), .B2(new_n633), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n982), .A2(new_n680), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n319), .A2(new_n219), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT50), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n203), .A2(new_n221), .ZN(new_n987));
  NOR4_X1   g0787(.A1(new_n986), .A2(new_n643), .A3(G45), .A4(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n687), .B1(new_n242), .B2(new_n469), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n643), .A2(new_n233), .A3(new_n283), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n233), .A2(G107), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n872), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n984), .A2(new_n993), .B1(new_n947), .B2(new_n963), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n966), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT106), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT106), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n966), .A2(new_n997), .A3(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(G393));
  OR2_X1    g0799(.A1(new_n950), .A2(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n950), .A2(KEYINPUT44), .ZN(new_n1001));
  AND3_X1   g0801(.A1(new_n627), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT45), .B1(new_n627), .B2(new_n936), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1000), .B(new_n1001), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n636), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(new_n947), .A3(new_n953), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n937), .A2(new_n685), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n710), .A2(G77), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n728), .A2(new_n760), .B1(new_n698), .B2(new_n889), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT51), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1009), .B1(new_n714), .B2(new_n203), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n352), .B(new_n1012), .C1(new_n319), .C2(new_n723), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n706), .A2(G143), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n719), .A2(G50), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G87), .A2(new_n717), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n283), .B1(new_n715), .B2(G283), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n775), .B2(new_n722), .C1(new_n739), .C2(new_n730), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G322), .B2(new_n706), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n718), .C1(new_n252), .C2(new_n766), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n699), .A2(G317), .B1(new_n700), .B2(G311), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT52), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1017), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n684), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n253), .A2(new_n687), .B1(G97), .B2(new_n638), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n872), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n680), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT107), .Z(new_n1029));
  NAND3_X1  g0829(.A1(new_n1008), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n636), .B1(new_n949), .B2(new_n952), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n964), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n639), .A3(new_n957), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(KEYINPUT108), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT108), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1006), .A2(new_n953), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n641), .B1(new_n1037), .B2(new_n964), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1036), .B1(new_n1038), .B2(new_n957), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1007), .B(new_n1030), .C1(new_n1035), .C2(new_n1039), .ZN(G390));
  OAI21_X1  g0840(.A(new_n833), .B1(new_n822), .B2(new_n823), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n814), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n818), .B1(new_n843), .B2(KEYINPUT39), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n749), .A2(new_n336), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n672), .A2(new_n618), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n821), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n799), .A2(new_n809), .B1(new_n1046), .B2(new_n833), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1042), .A2(new_n1043), .B1(new_n814), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n846), .A2(G330), .A3(new_n845), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n849), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT109), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n755), .A2(new_n844), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT109), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n812), .A2(new_n818), .B1(new_n1041), .B2(new_n814), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1047), .A2(new_n814), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1055), .B(new_n1050), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1052), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT111), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1052), .A2(new_n1058), .A3(KEYINPUT111), .A4(new_n1054), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n839), .A2(new_n588), .A3(new_n856), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n833), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1049), .A2(KEYINPUT110), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n750), .B1(new_n1049), .B2(KEYINPUT110), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1046), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n1053), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n833), .B1(new_n755), .B2(new_n750), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n824), .B1(new_n1070), .B2(new_n1050), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1063), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1061), .A2(new_n1062), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT112), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1061), .A2(KEYINPUT112), .A3(new_n1062), .A4(new_n1073), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1052), .A2(new_n1058), .A3(new_n1072), .A4(new_n1054), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1076), .A2(new_n639), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1043), .A2(new_n779), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n383), .A2(new_n780), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT54), .B(G143), .Z(new_n1082));
  AOI22_X1  g0882(.A1(new_n723), .A2(new_n1082), .B1(new_n719), .B2(G137), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT113), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n714), .A2(new_n889), .ZN(new_n1085));
  XOR2_X1   g0885(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1086));
  OAI21_X1  g0886(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n706), .A2(G125), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n352), .B1(new_n700), .B2(G132), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n699), .A2(G128), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n735), .A2(new_n219), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n766), .A2(new_n760), .ZN(new_n1094));
  NOR4_X1   g0894(.A1(new_n1087), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n706), .A2(G294), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n283), .B1(new_n700), .B2(G116), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n716), .A2(new_n1096), .A3(new_n1009), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n730), .A2(new_n567), .B1(new_n484), .B2(new_n722), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT115), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n698), .A2(new_n734), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1098), .A2(new_n1100), .A3(new_n764), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n684), .B1(new_n1095), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1080), .A2(new_n680), .A3(new_n1081), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1059), .B2(new_n946), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT116), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1079), .A2(new_n1106), .ZN(G378));
  INV_X1    g0907(.A(new_n1063), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1078), .A2(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n819), .A2(new_n835), .A3(new_n836), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n318), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n301), .A2(new_n785), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1111), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n311), .A2(new_n317), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(new_n311), .B2(new_n317), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n316), .B(new_n1111), .C1(new_n308), .C2(new_n310), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1113), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1117), .A2(new_n1120), .A3(KEYINPUT120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT120), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n631), .B(new_n1123), .C1(new_n848), .C2(new_n853), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n858), .B2(G330), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1110), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1123), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n854), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1129), .B(new_n837), .C1(new_n854), .C2(new_n1125), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1109), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT57), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1109), .A2(new_n1131), .A3(KEYINPUT57), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n639), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1127), .A2(new_n1130), .A3(new_n947), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n717), .A2(G58), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT117), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n283), .B1(new_n706), .B2(G283), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n215), .C2(new_n728), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G77), .B2(new_n715), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n766), .A2(new_n203), .B1(new_n322), .B2(new_n722), .ZN(new_n1143));
  AOI211_X1 g0943(.A(G41), .B(new_n1143), .C1(G97), .C2(new_n719), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(new_n252), .C2(new_n698), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT58), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n219), .B1(new_n350), .B2(G41), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n766), .A2(new_n889), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n730), .A2(new_n767), .B1(new_n759), .B2(new_n722), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n715), .A2(new_n1082), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(KEYINPUT118), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n700), .A2(G128), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(KEYINPUT118), .C2(new_n1150), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1148), .B(new_n1153), .C1(G125), .C2(new_n699), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT59), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G33), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1157));
  AOI21_X1  g0957(.A(G41), .B1(new_n706), .B2(G124), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n760), .C2(new_n735), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1146), .B(new_n1147), .C1(new_n1156), .C2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT119), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n684), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n780), .A2(new_n219), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1123), .A2(new_n779), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1162), .A2(new_n680), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1137), .A2(KEYINPUT121), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT121), .B1(new_n1137), .B2(new_n1165), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1136), .A2(new_n1168), .ZN(G375));
  NAND3_X1  g0969(.A1(new_n1069), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n959), .B(KEYINPUT122), .Z(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1073), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n891), .B1(new_n329), .B2(new_n723), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n484), .B2(new_n714), .C1(new_n739), .C2(new_n705), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n730), .A2(new_n252), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n698), .A2(new_n775), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n352), .B1(new_n766), .B2(new_n322), .C1(new_n728), .C2(new_n734), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n715), .A2(G159), .B1(new_n706), .B2(G128), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1139), .B(new_n1180), .C1(new_n767), .C2(new_n698), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n722), .A2(new_n889), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n766), .A2(new_n219), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n352), .B1(new_n719), .B2(new_n1082), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n759), .B2(new_n728), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n684), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n779), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n680), .B(new_n1187), .C1(new_n833), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n203), .B2(new_n780), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n947), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1173), .A2(new_n1192), .ZN(G381));
  NOR2_X1   g0993(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1109), .A2(new_n1131), .A3(KEYINPUT57), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1109), .B2(new_n1131), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1194), .B1(new_n1197), .B2(new_n639), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1077), .A2(new_n639), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1078), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1105), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n909), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n942), .A2(new_n943), .A3(new_n932), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n943), .B1(new_n942), .B2(new_n932), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n958), .A2(new_n959), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n946), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1204), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(G381), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n996), .A2(new_n744), .A3(new_n998), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G390), .A2(G384), .A3(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1203), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(G407));
  INV_X1    g1014(.A(G213), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1203), .B2(new_n616), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(G407), .ZN(G409));
  NOR2_X1   g1017(.A1(new_n1215), .A2(G343), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1198), .A2(G378), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1105), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1137), .B(new_n1165), .C1(new_n1132), .C2(new_n1171), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1079), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1218), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n641), .B1(new_n1170), .B2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n1073), .C1(new_n1224), .C2(new_n1170), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1226), .A2(G384), .A3(new_n1192), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G384), .B1(new_n1226), .B2(new_n1192), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT63), .B1(new_n1223), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT116), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1105), .B(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1222), .B1(new_n1233), .B2(G375), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1218), .ZN(new_n1235));
  AND4_X1   g1035(.A1(KEYINPUT63), .A2(new_n1234), .A3(new_n1235), .A4(new_n1229), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1230), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1229), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(G2897), .A3(new_n1218), .ZN(new_n1239));
  INV_X1    g1039(.A(G2897), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1229), .B1(new_n1240), .B2(new_n1235), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(KEYINPUT123), .B1(new_n1223), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT123), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1198), .A2(G378), .B1(new_n1202), .B2(new_n1221), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1244), .B(new_n1245), .C1(new_n1246), .C2(new_n1218), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n998), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n997), .B1(new_n966), .B2(new_n994), .ZN(new_n1250));
  OAI21_X1  g1050(.A(G396), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n1212), .A3(KEYINPUT124), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(G390), .B2(new_n1210), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1251), .A2(new_n1212), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1030), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1034), .A2(KEYINPUT108), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1038), .A2(new_n1036), .A3(new_n957), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(G387), .A3(new_n1258), .A4(new_n1007), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1253), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G390), .A2(new_n1210), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1252), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT61), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT125), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1237), .A2(new_n1248), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1234), .A2(new_n1235), .A3(new_n1229), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1244), .B1(new_n1246), .B2(new_n1218), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1234), .A2(new_n1272), .A3(new_n1235), .A4(new_n1229), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1262), .A2(KEYINPUT126), .A3(new_n1264), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G387), .B1(new_n1258), .B2(new_n1007), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1278), .B2(new_n1263), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1274), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1267), .A2(new_n1281), .ZN(G405));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1275), .A2(new_n1283), .A3(new_n1279), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1229), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G375), .A2(new_n1202), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1219), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT126), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1278), .A2(new_n1276), .A3(new_n1263), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT127), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1275), .A2(new_n1279), .A3(new_n1283), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1238), .A3(new_n1292), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1286), .A2(new_n1288), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1288), .B1(new_n1286), .B2(new_n1293), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G402));
endmodule


