//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT67), .B(G244), .Z(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n203), .A2(G50), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n218), .A2(KEYINPUT1), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OR3_X1    g0024(.A1(new_n209), .A2(KEYINPUT65), .A3(G13), .ZN(new_n225));
  OAI21_X1  g0025(.A(KEYINPUT65), .B1(new_n209), .B2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT66), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n224), .B(new_n230), .C1(KEYINPUT1), .C2(new_n218), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n219), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n249), .B1(new_n250), .B2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G13), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n253), .A2(new_n220), .A3(G1), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n252), .B1(G50), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n220), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT72), .A2(G58), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n262), .B(new_n263), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n257), .B1(new_n258), .B2(new_n260), .C1(new_n261), .C2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n256), .B1(new_n265), .B2(new_n249), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT69), .ZN(new_n267));
  AND2_X1   g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n219), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G41), .A2(G45), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n272), .A2(KEYINPUT69), .A3(G1), .A4(G13), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n269), .A2(G274), .A3(new_n271), .A4(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT71), .B1(new_n270), .B2(G1), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT71), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n276), .B(new_n250), .C1(G41), .C2(G45), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n269), .A2(new_n275), .A3(new_n273), .A4(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(KEYINPUT70), .B(G226), .Z(new_n279));
  OAI21_X1  g0079(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1698), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G222), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n284), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n283), .B2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G223), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n286), .B1(new_n211), .B2(new_n287), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n280), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n298), .B1(KEYINPUT73), .B2(new_n301), .ZN(new_n302));
  AOI211_X1 g0102(.A(new_n266), .B(new_n302), .C1(KEYINPUT73), .C2(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n266), .A2(KEYINPUT9), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n304), .B(KEYINPUT75), .Z(new_n305));
  NAND2_X1  g0105(.A1(new_n295), .A2(G190), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT74), .B(G200), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n306), .B1(new_n307), .B2(new_n295), .C1(KEYINPUT9), .C2(new_n266), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n305), .A2(KEYINPUT10), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n305), .B2(new_n308), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT16), .ZN(new_n312));
  INV_X1    g0112(.A(G58), .ZN(new_n313));
  INV_X1    g0113(.A(G68), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(G20), .B1(new_n315), .B2(new_n202), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n259), .A2(G159), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n287), .B2(G20), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n314), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT79), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n319), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g0128(.A(KEYINPUT79), .B(new_n314), .C1(new_n321), .C2(new_n325), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n312), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n249), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n326), .A2(new_n318), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n264), .A2(new_n255), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n251), .B2(new_n264), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT80), .ZN(new_n337));
  INV_X1    g0137(.A(G232), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n274), .B1(new_n278), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT81), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G87), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n291), .A2(new_n288), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G226), .B2(new_n288), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n341), .B1(new_n343), .B2(new_n324), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n339), .A2(new_n340), .B1(new_n294), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(KEYINPUT81), .B(new_n274), .C1(new_n278), .C2(new_n338), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G190), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n339), .A2(new_n340), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n294), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G200), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n334), .A2(new_n337), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT17), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND4_X1   g0154(.A1(G179), .A2(new_n348), .A3(new_n346), .A4(new_n349), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n300), .B1(new_n345), .B2(new_n346), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT80), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n336), .B(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n330), .B2(new_n333), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT18), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n350), .A2(G169), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n296), .B2(new_n350), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n287), .A2(new_n320), .A3(G20), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT7), .B1(new_n324), .B2(new_n220), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n318), .B1(new_n366), .B2(KEYINPUT79), .ZN(new_n367));
  INV_X1    g0167(.A(new_n329), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT16), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(KEYINPUT16), .A3(new_n319), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n249), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n337), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n363), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n360), .A2(KEYINPUT17), .A3(new_n347), .A4(new_n351), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n354), .A2(new_n361), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n254), .A2(new_n314), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT12), .B1(new_n378), .B2(KEYINPUT76), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(KEYINPUT76), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(KEYINPUT76), .A3(KEYINPUT12), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n314), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n211), .B2(new_n261), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n249), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n386), .A2(new_n387), .B1(G68), .B2(new_n251), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n383), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G97), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G226), .A2(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n338), .B2(G1698), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n395), .B2(new_n287), .ZN(new_n396));
  INV_X1    g0196(.A(G238), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n293), .A2(new_n396), .B1(new_n278), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n274), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT13), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n278), .A2(new_n397), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n338), .A2(G1698), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G226), .B2(G1698), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n392), .B1(new_n404), .B2(new_n324), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n294), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n401), .A2(new_n402), .A3(new_n274), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT14), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n408), .B2(new_n296), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n409), .B1(new_n408), .B2(G169), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n391), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n274), .B1(new_n278), .B2(new_n210), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n285), .A2(G232), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n415), .B1(new_n206), .B2(new_n287), .C1(new_n290), .C2(new_n397), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(new_n294), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n417), .A2(G169), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT8), .B(G58), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n419), .A2(new_n260), .B1(new_n220), .B2(new_n211), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT15), .B(G87), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n261), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n249), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n251), .A2(G77), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n424), .C1(G77), .C2(new_n255), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n296), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n425), .B1(new_n417), .B2(G190), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n307), .B2(new_n417), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n311), .A2(new_n377), .A3(new_n413), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n400), .A2(new_n407), .A3(G190), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n390), .ZN(new_n435));
  INV_X1    g0235(.A(G200), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n400), .B2(new_n407), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n433), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n408), .A2(G200), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(KEYINPUT77), .A3(new_n434), .A4(new_n390), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT78), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n438), .B2(new_n440), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n432), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n269), .A2(new_n273), .ZN(new_n447));
  INV_X1    g0247(.A(G41), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n250), .B(G45), .C1(new_n448), .C2(KEYINPUT5), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(G264), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT83), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n450), .B1(new_n449), .B2(new_n453), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n447), .A2(G274), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(G250), .B(new_n288), .C1(new_n322), .C2(new_n323), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G294), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(G257), .B(G1698), .C1(new_n322), .C2(new_n323), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT88), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT88), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n287), .A2(new_n462), .A3(G257), .A4(G1698), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT89), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n294), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g0266(.A(KEYINPUT89), .B(new_n459), .C1(new_n461), .C2(new_n463), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n452), .B(new_n456), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n436), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n457), .A2(new_n458), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n462), .B1(new_n289), .B2(G257), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n460), .A2(KEYINPUT88), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n464), .A2(new_n465), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(new_n294), .ZN(new_n476));
  INV_X1    g0276(.A(G190), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n456), .A4(new_n452), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n469), .A2(KEYINPUT90), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n452), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n293), .B1(new_n473), .B2(KEYINPUT89), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n475), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT90), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n477), .A4(new_n456), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT23), .B1(new_n206), .B2(G20), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n485), .A2(new_n486), .B1(G20), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n220), .B(G87), .C1(new_n322), .C2(new_n323), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT22), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT22), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n287), .A2(new_n491), .A3(new_n220), .A4(G87), .ZN(new_n492));
  AOI211_X1 g0292(.A(KEYINPUT24), .B(new_n488), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n490), .A2(new_n492), .ZN(new_n495));
  INV_X1    g0295(.A(new_n488), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n249), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT87), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT87), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(new_n249), .C1(new_n493), .C2(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n250), .A2(G33), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n255), .A2(new_n331), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT25), .B1(new_n254), .B2(new_n206), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n505), .A2(G107), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n479), .A2(new_n484), .A3(new_n502), .A4(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n255), .A2(G97), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n504), .B2(new_n205), .ZN(new_n513));
  XNOR2_X1  g0313(.A(G97), .B(G107), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n515), .A2(new_n205), .A3(G107), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n520));
  OAI21_X1  g0320(.A(G107), .B1(new_n364), .B2(new_n365), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n513), .B1(new_n522), .B2(new_n249), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(G1698), .C1(new_n322), .C2(new_n323), .ZN(new_n525));
  OAI211_X1 g0325(.A(G244), .B(new_n288), .C1(new_n322), .C2(new_n323), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT4), .B1(new_n285), .B2(G244), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n294), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n447), .A2(G257), .A3(new_n451), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(G190), .A3(new_n456), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n456), .A2(new_n531), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT82), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n526), .A2(new_n527), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n537), .A3(new_n524), .A4(new_n525), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(KEYINPUT82), .A3(new_n294), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n533), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n523), .B(new_n532), .C1(new_n540), .C2(new_n436), .ZN(new_n541));
  INV_X1    g0341(.A(new_n533), .ZN(new_n542));
  INV_X1    g0342(.A(new_n539), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT82), .B1(new_n538), .B2(new_n294), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(new_n296), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n530), .A2(new_n456), .A3(new_n531), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n517), .B1(new_n515), .B2(new_n514), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n547), .A2(new_n220), .B1(new_n211), .B2(new_n260), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n206), .B1(new_n321), .B2(new_n325), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n249), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n511), .B1(new_n505), .B2(G97), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n546), .A2(new_n300), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n541), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n287), .A2(new_n220), .A3(G68), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n220), .B1(new_n392), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G87), .B2(new_n207), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n261), .B2(new_n205), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n249), .B1(new_n254), .B2(new_n421), .ZN(new_n561));
  INV_X1    g0361(.A(new_n421), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n505), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT85), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  INV_X1    g0367(.A(G45), .ZN(new_n568));
  OR3_X1    g0368(.A1(new_n568), .A2(G1), .A3(G274), .ZN(new_n569));
  INV_X1    g0369(.A(G250), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n568), .B2(G1), .ZN(new_n571));
  AND4_X1   g0371(.A1(new_n269), .A2(new_n569), .A3(new_n273), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n397), .A2(new_n288), .ZN(new_n573));
  INV_X1    g0373(.A(G244), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G1698), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n575), .C1(new_n322), .C2(new_n323), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n293), .B1(new_n576), .B2(new_n487), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n567), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n269), .A2(new_n569), .A3(new_n273), .A4(new_n571), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G238), .A2(G1698), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n574), .B2(G1698), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(new_n287), .B1(G33), .B2(G116), .ZN(new_n582));
  OAI211_X1 g0382(.A(KEYINPUT84), .B(new_n579), .C1(new_n582), .C2(new_n293), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n578), .A2(new_n296), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(G169), .B1(new_n578), .B2(new_n583), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n566), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(new_n583), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n300), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n578), .A2(new_n583), .A3(new_n296), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(KEYINPUT85), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n565), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n587), .A2(new_n477), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n505), .A2(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n561), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n307), .B1(new_n578), .B2(new_n583), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n554), .A2(new_n591), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n502), .A2(new_n509), .ZN(new_n598));
  INV_X1    g0398(.A(new_n468), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n296), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n468), .A2(new_n300), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n285), .A2(G257), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n289), .A2(G264), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n324), .A2(G303), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n294), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n447), .A2(G270), .A3(new_n451), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n456), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G169), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n255), .A2(G116), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n504), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n248), .A2(new_n219), .B1(G20), .B2(new_n614), .ZN(new_n616));
  AOI21_X1  g0416(.A(G20), .B1(G33), .B2(G283), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n282), .A2(G97), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT86), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT86), .B1(new_n617), .B2(new_n618), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(KEYINPUT20), .B(new_n616), .C1(new_n619), .C2(new_n620), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n615), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n603), .B1(new_n611), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n610), .A2(new_n296), .ZN(new_n627));
  INV_X1    g0427(.A(new_n615), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n624), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n630), .A2(KEYINPUT21), .A3(new_n610), .A4(G169), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n626), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n610), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G190), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n630), .B1(G200), .B2(new_n610), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n510), .A2(new_n597), .A3(new_n602), .A4(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n446), .A2(new_n638), .ZN(G372));
  NAND2_X1  g0439(.A1(new_n309), .A2(new_n310), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n354), .A2(new_n375), .ZN(new_n641));
  INV_X1    g0441(.A(new_n428), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n438), .A2(new_n440), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n644), .B2(new_n413), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n361), .A2(new_n374), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n303), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n446), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n586), .A2(new_n590), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n564), .ZN(new_n653));
  INV_X1    g0453(.A(new_n553), .ZN(new_n654));
  INV_X1    g0454(.A(new_n596), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT26), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n579), .B1(new_n582), .B2(new_n293), .ZN(new_n658));
  INV_X1    g0458(.A(new_n307), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n561), .A3(new_n593), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT91), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n578), .A2(new_n583), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G190), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n660), .A2(new_n561), .A3(new_n665), .A4(new_n593), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n561), .A2(new_n563), .B1(new_n300), .B2(new_n658), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n589), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n553), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n657), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n669), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n553), .A2(new_n541), .A3(new_n667), .A4(new_n669), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n484), .A2(new_n502), .A3(new_n509), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n679), .B2(new_n479), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n631), .A2(new_n632), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n602), .A2(new_n626), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n676), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n650), .B1(new_n651), .B2(new_n685), .ZN(G369));
  NAND3_X1  g0486(.A1(new_n250), .A2(new_n220), .A3(G13), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n598), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n510), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n602), .ZN(new_n695));
  INV_X1    g0495(.A(new_n602), .ZN(new_n696));
  INV_X1    g0496(.A(new_n692), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n637), .B1(new_n625), .B2(new_n697), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n633), .A2(new_n630), .A3(new_n692), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n696), .B1(new_n510), .B2(new_n693), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n633), .A2(new_n697), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n698), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0511(.A(new_n227), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n713), .A2(new_n250), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n223), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n713), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT28), .Z(new_n719));
  INV_X1    g0519(.A(KEYINPUT99), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n591), .A2(new_n553), .A3(new_n596), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT98), .B1(new_n721), .B2(KEYINPUT26), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT98), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n656), .A2(new_n723), .A3(new_n672), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n670), .A2(new_n672), .A3(new_n553), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n683), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n720), .B1(new_n728), .B2(new_n697), .ZN(new_n729));
  AOI211_X1 g0529(.A(KEYINPUT99), .B(new_n692), .C1(new_n727), .C2(new_n683), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT29), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n692), .B1(new_n675), .B2(new_n683), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n476), .A2(KEYINPUT94), .A3(new_n663), .A4(new_n452), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(new_n627), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT95), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT94), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n452), .B1(new_n466), .B2(new_n467), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n587), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n546), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n737), .A2(new_n738), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n741), .A2(new_n627), .A3(new_n736), .A4(new_n743), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n546), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n741), .A2(new_n627), .A3(new_n748), .A4(new_n736), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n742), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT96), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n658), .A2(new_n296), .ZN(new_n753));
  NOR4_X1   g0553(.A1(new_n599), .A2(new_n634), .A3(new_n540), .A4(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n749), .A2(KEYINPUT96), .A3(new_n742), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n747), .A2(new_n752), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT31), .B1(new_n757), .B2(new_n692), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT97), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n749), .A2(KEYINPUT96), .A3(new_n742), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT96), .B1(new_n749), .B2(new_n742), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n754), .B1(new_n744), .B2(new_n746), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n697), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(KEYINPUT97), .B1(new_n765), .B2(KEYINPUT31), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n747), .A2(new_n755), .A3(new_n750), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n638), .A2(new_n697), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n760), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G330), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n735), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n719), .B1(new_n772), .B2(G1), .ZN(G364));
  NOR2_X1   g0573(.A1(new_n253), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n250), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n713), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n703), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n701), .A2(new_n700), .A3(new_n702), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n777), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n220), .A2(G190), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(new_n296), .A3(new_n436), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT101), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT101), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n659), .A2(G20), .A3(new_n296), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n477), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n787), .A2(G329), .B1(new_n789), .B2(G303), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n296), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n782), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n324), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(G20), .A3(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n794), .B1(G322), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n788), .A2(G190), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n790), .B(new_n797), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n220), .A2(new_n296), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G190), .ZN(new_n804));
  INV_X1    g0604(.A(G317), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(KEYINPUT33), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n805), .A2(KEYINPUT33), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n477), .A2(G179), .A3(G200), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n220), .ZN(new_n811));
  INV_X1    g0611(.A(G326), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n803), .A2(new_n477), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n808), .B1(new_n809), .B2(new_n811), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  OR3_X1    g0616(.A1(new_n786), .A2(KEYINPUT32), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT32), .B1(new_n786), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n804), .A2(G68), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n811), .A2(new_n205), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G50), .B2(new_n813), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n789), .A2(G87), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n799), .A2(G107), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n796), .A2(G58), .ZN(new_n825));
  INV_X1    g0625(.A(new_n792), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n324), .B1(new_n826), .B2(G77), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n801), .A2(new_n815), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n219), .B1(G20), .B2(new_n300), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(G13), .A2(G33), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(G20), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n830), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n712), .A2(new_n287), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(G45), .B2(new_n223), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n243), .B2(G45), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT100), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n227), .A2(new_n287), .ZN(new_n840));
  INV_X1    g0640(.A(G355), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n840), .A2(new_n841), .B1(G116), .B2(new_n227), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n838), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n839), .B2(new_n842), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n781), .B(new_n831), .C1(new_n835), .C2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n701), .A2(new_n702), .A3(new_n834), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n780), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  NOR2_X1   g0649(.A1(new_n830), .A2(new_n832), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT102), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n799), .A2(G87), .ZN(new_n852));
  INV_X1    g0652(.A(new_n789), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n206), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n324), .B1(new_n792), .B2(new_n614), .C1(new_n809), .C2(new_n795), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n820), .B(new_n855), .C1(G303), .C2(new_n813), .ZN(new_n856));
  INV_X1    g0656(.A(new_n804), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n856), .B1(new_n861), .B2(new_n798), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n854), .B(new_n862), .C1(G311), .C2(new_n787), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n796), .A2(G143), .B1(new_n826), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n864), .B1(new_n857), .B2(new_n258), .C1(new_n865), .C2(new_n814), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT104), .Z(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n868));
  INV_X1    g0668(.A(G132), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n287), .B1(new_n786), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT105), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n789), .A2(G50), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n872), .B1(new_n313), .B2(new_n811), .C1(new_n800), .C2(new_n314), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n868), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n863), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n830), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n777), .B1(G77), .B2(new_n851), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n642), .A2(new_n697), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n425), .A2(new_n692), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n430), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n428), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n878), .B1(new_n832), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n883), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n732), .B(new_n885), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n771), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n777), .B1(new_n771), .B2(new_n886), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(G384));
  NOR2_X1   g0690(.A1(new_n774), .A2(new_n250), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n757), .A2(new_n768), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n597), .A2(new_n637), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(new_n510), .A3(new_n602), .A4(new_n697), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n892), .B(new_n894), .C1(new_n765), .C2(KEYINPUT31), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n390), .A2(new_n697), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n413), .A2(new_n643), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n411), .A2(new_n412), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n443), .B2(new_n444), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n902), .B2(new_n896), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n883), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n312), .B1(new_n326), .B2(new_n318), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n370), .A3(new_n249), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n336), .ZN(new_n908));
  INV_X1    g0708(.A(new_n690), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n376), .A2(new_n905), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n905), .B1(new_n376), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n908), .B1(new_n356), .B2(new_n355), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n352), .A2(new_n915), .A3(new_n910), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT37), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT107), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(KEYINPUT107), .A3(KEYINPUT37), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n363), .A2(new_n372), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n372), .A2(new_n909), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT37), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n352), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n914), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n376), .A2(new_n911), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT106), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n376), .A2(new_n905), .A3(new_n911), .ZN(new_n929));
  AND4_X1   g0729(.A1(KEYINPUT38), .A2(new_n925), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n895), .B(new_n904), .C1(new_n926), .C2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT110), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT110), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n925), .A2(new_n928), .A3(KEYINPUT38), .A4(new_n929), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT38), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n360), .A2(new_n690), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT37), .B1(new_n940), .B2(KEYINPUT108), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n921), .A2(new_n922), .A3(new_n352), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n376), .A2(new_n940), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n932), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n643), .A2(KEYINPUT78), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n900), .B1(new_n949), .B2(new_n442), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n898), .B1(new_n950), .B2(new_n897), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n885), .ZN(new_n952));
  INV_X1    g0752(.A(new_n758), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n638), .A2(new_n697), .B1(new_n757), .B2(new_n768), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n948), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n937), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n892), .A2(new_n894), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n758), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n651), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n700), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT111), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n963), .A2(new_n964), .B1(new_n957), .B2(new_n961), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n963), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n731), .A2(new_n446), .A3(new_n734), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT109), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n731), .A2(KEYINPUT109), .A3(new_n446), .A4(new_n734), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n649), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n925), .A2(new_n928), .A3(new_n929), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n939), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(KEYINPUT39), .A3(new_n938), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT39), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n946), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n900), .A2(new_n391), .A3(new_n697), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n974), .A2(new_n938), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(G200), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n523), .A2(new_n532), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n983), .A2(new_n984), .B1(new_n545), .B2(new_n552), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n667), .A2(new_n669), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n469), .A2(KEYINPUT90), .A3(new_n478), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n985), .B(new_n986), .C1(new_n987), .C2(new_n678), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n502), .A2(new_n509), .B1(new_n300), .B2(new_n468), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n633), .B1(new_n989), .B2(new_n600), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n669), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n885), .B(new_n697), .C1(new_n991), .C2(new_n674), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n903), .B1(new_n992), .B2(new_n879), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n981), .A2(new_n993), .B1(new_n646), .B2(new_n690), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n980), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n972), .B(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n891), .B1(new_n967), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n997), .B2(new_n967), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n614), .B(new_n222), .C1(new_n519), .C2(KEYINPUT35), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT35), .B2(new_n519), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT36), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n223), .A2(new_n211), .A3(new_n315), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n201), .A2(new_n314), .ZN(new_n1004));
  OAI211_X1 g0804(.A(G1), .B(new_n253), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n999), .A2(new_n1002), .A3(new_n1005), .ZN(G367));
  NOR3_X1   g0806(.A1(new_n238), .A2(new_n712), .A3(new_n287), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n835), .B1(new_n227), .B2(new_n421), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n777), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT46), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n789), .A2(G116), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n860), .A2(G294), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1013));
  INV_X1    g0813(.A(G303), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n324), .B1(new_n795), .B2(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n814), .A2(new_n793), .B1(new_n206), .B2(new_n811), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G283), .C2(new_n826), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n799), .A2(G97), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n805), .C2(new_n786), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n799), .A2(G77), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n786), .B2(new_n865), .C1(new_n853), .C2(new_n313), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n811), .A2(new_n314), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n201), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n287), .B1(new_n258), .B2(new_n795), .C1(new_n1023), .C2(new_n792), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(G143), .C2(new_n813), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n861), .B2(new_n816), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1013), .A2(new_n1019), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1009), .B1(new_n1028), .B2(new_n830), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n834), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n594), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(new_n697), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n670), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n676), .A2(new_n1032), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1029), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT112), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n985), .B1(new_n523), .B2(new_n697), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n654), .A2(new_n692), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n709), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT44), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n709), .A2(KEYINPUT44), .A3(new_n1041), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT45), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n709), .B2(new_n1041), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT92), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n707), .B(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(new_n695), .A3(new_n698), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1051), .A2(KEYINPUT45), .A3(new_n698), .A4(new_n1040), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1037), .B(new_n705), .C1(new_n1046), .C2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1044), .A2(new_n1045), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n704), .B1(new_n1055), .B2(KEYINPUT112), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n699), .B(new_n1050), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(new_n703), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1059), .A2(new_n771), .A3(new_n735), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n772), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n713), .B(KEYINPUT41), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n776), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1035), .A2(KEYINPUT43), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n699), .A2(new_n1050), .A3(new_n1040), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT42), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n696), .A2(new_n541), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n692), .B1(new_n1067), .B2(new_n553), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1065), .B2(KEYINPUT42), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1064), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1035), .A2(KEYINPUT43), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n704), .B2(new_n1041), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1073), .A2(new_n705), .A3(new_n1040), .A4(new_n1074), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1036), .B1(new_n1063), .B2(new_n1078), .ZN(G387));
  NAND2_X1  g0879(.A1(new_n1059), .A2(new_n776), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n324), .B1(new_n786), .B2(new_n812), .C1(new_n800), .C2(new_n614), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n811), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n789), .A2(G294), .B1(G283), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n796), .A2(G317), .B1(new_n826), .B2(G303), .ZN(new_n1084));
  INV_X1    g0884(.A(G322), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n814), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n860), .B2(G311), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT48), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT114), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(KEYINPUT48), .B2(new_n1087), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1092), .A2(KEYINPUT49), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(KEYINPUT49), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1081), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n324), .B1(new_n796), .B2(G50), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1018), .B(new_n1096), .C1(new_n314), .C2(new_n792), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n789), .A2(G77), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n258), .B2(new_n786), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n264), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1100), .A2(new_n804), .B1(new_n813), .B2(G159), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n421), .B2(new_n811), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1097), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n830), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(G45), .B(new_n715), .C1(G68), .C2(G77), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT113), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n419), .A2(G50), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT50), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1105), .A2(KEYINPUT113), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n836), .B1(new_n568), .B2(new_n235), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(G107), .B2(new_n227), .C1(new_n714), .C2(new_n840), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n781), .B1(new_n1112), .B2(new_n835), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1104), .B(new_n1113), .C1(new_n699), .C2(new_n1030), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1060), .A2(new_n713), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n772), .A2(new_n1059), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1080), .B(new_n1114), .C1(new_n1115), .C2(new_n1116), .ZN(G393));
  XNOR2_X1  g0917(.A(new_n1055), .B(new_n704), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1118), .A2(new_n775), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n836), .A2(new_n246), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n835), .C1(new_n205), .C2(new_n227), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT115), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n781), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n853), .A2(new_n798), .B1(new_n1085), .B2(new_n786), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n287), .B1(new_n826), .B2(G294), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n824), .B(new_n1127), .C1(new_n614), .C2(new_n811), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(G303), .C2(new_n860), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n813), .A2(G317), .B1(new_n796), .B2(G311), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT52), .Z(new_n1131));
  OAI22_X1  g0931(.A1(new_n814), .A2(new_n258), .B1(new_n816), .B2(new_n795), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n201), .C2(new_n860), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n787), .A2(G143), .B1(new_n789), .B2(G68), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n811), .A2(new_n211), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n419), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n324), .B1(new_n826), .B2(new_n1140), .ZN(new_n1141));
  AND4_X1   g0941(.A1(new_n852), .A2(new_n1137), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1129), .A2(new_n1131), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1125), .B1(new_n877), .B2(new_n1143), .C1(new_n1040), .C2(new_n1030), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n713), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1118), .A2(new_n1060), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1119), .B(new_n1144), .C1(new_n1145), .C2(new_n1146), .ZN(G390));
  AOI21_X1  g0947(.A(new_n596), .B1(new_n652), .B2(new_n564), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT26), .B1(new_n1148), .B2(new_n654), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n725), .B1(new_n1149), .B2(new_n723), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n991), .B1(new_n722), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT99), .B1(new_n1151), .B2(new_n692), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n728), .A2(new_n720), .A3(new_n697), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n879), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n951), .B(KEYINPUT117), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n882), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n947), .A2(new_n979), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n975), .A2(new_n977), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n993), .A2(new_n979), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1156), .A2(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n770), .A2(G330), .A3(new_n885), .A4(new_n951), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n959), .A2(new_n700), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n904), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1154), .A2(new_n882), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n895), .A2(G330), .A3(new_n885), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n903), .B(KEYINPUT117), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1166), .A2(new_n1161), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n769), .B1(new_n758), .B2(new_n759), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n765), .A2(KEYINPUT97), .A3(KEYINPUT31), .ZN(new_n1172));
  OAI211_X1 g0972(.A(G330), .B(new_n885), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1173), .A2(new_n903), .B1(new_n1163), .B2(new_n904), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n992), .A2(new_n879), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1170), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n651), .A2(new_n700), .A3(new_n959), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n972), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1165), .A2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n649), .B(new_n1178), .C1(new_n970), .C2(new_n971), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1159), .A2(new_n1158), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n904), .A3(new_n1163), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1182), .A2(new_n1186), .A3(new_n1162), .A4(new_n1177), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1181), .A2(new_n1187), .A3(new_n713), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1183), .A2(new_n1184), .A3(new_n1161), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1158), .A2(new_n832), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n777), .B1(new_n851), .B2(new_n1100), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n860), .A2(G107), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n787), .A2(G294), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G68), .A2(new_n799), .B1(new_n789), .B2(G87), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n324), .B1(new_n792), .B2(new_n205), .C1(new_n614), .C2(new_n795), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1138), .B(new_n1197), .C1(G283), .C2(new_n813), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n811), .A2(new_n816), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT54), .B(G143), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n287), .B1(new_n792), .B2(new_n1201), .C1(new_n869), .C2(new_n795), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G128), .C2(new_n813), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n787), .A2(G125), .B1(new_n799), .B2(new_n201), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n865), .C2(new_n861), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n789), .A2(G150), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT53), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1199), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1193), .B1(new_n1208), .B2(new_n830), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1191), .A2(new_n776), .B1(new_n1192), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1188), .A2(new_n1210), .ZN(G378));
  NOR2_X1   g1011(.A1(new_n266), .A2(new_n690), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT121), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n311), .B(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1215));
  XOR2_X1   g1015(.A(new_n1214), .B(new_n1215), .Z(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n700), .B1(new_n948), .B2(new_n955), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n995), .B1(new_n937), .B2(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(KEYINPUT110), .B(KEYINPUT40), .C1(new_n955), .C2(new_n981), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n935), .B1(new_n931), .B2(new_n932), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n995), .B(new_n1218), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1217), .B1(new_n1219), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n996), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1222), .A3(new_n1216), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n776), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n796), .A2(G107), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT118), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n814), .A2(new_n614), .B1(new_n205), .B2(new_n857), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n324), .A2(new_n448), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1233), .B(new_n1022), .C1(new_n562), .C2(new_n826), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n787), .A2(G283), .B1(new_n799), .B2(G58), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1098), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT58), .ZN(new_n1237));
  AOI21_X1  g1037(.A(G50), .B1(new_n282), .B2(new_n448), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1236), .A2(new_n1237), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT119), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1201), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n789), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n804), .A2(G132), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G150), .A2(new_n1082), .B1(new_n813), .B2(G125), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n796), .A2(G128), .B1(new_n826), .B2(G137), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT59), .Z(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(KEYINPUT120), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(KEYINPUT120), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n799), .A2(G159), .ZN(new_n1250));
  AOI211_X1 g1050(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1240), .B1(new_n1237), .B2(new_n1236), .C1(new_n1248), .C2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n830), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n851), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n781), .B1(new_n1255), .B2(new_n1023), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(new_n1216), .C2(new_n833), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1228), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1227), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1216), .B1(new_n1226), .B2(new_n1222), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1187), .A2(new_n1182), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT57), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1224), .A2(KEYINPUT57), .A3(new_n1227), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n733), .B1(new_n1265), .B2(KEYINPUT29), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT109), .B1(new_n1266), .B2(new_n446), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n971), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n650), .B(new_n1179), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1191), .B2(new_n1177), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n713), .B1(new_n1264), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1258), .B1(new_n1263), .B2(new_n1271), .ZN(G375));
  AOI21_X1  g1072(.A(new_n781), .B1(new_n1255), .B2(new_n314), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n861), .A2(new_n614), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n1020), .B1(new_n786), .B2(new_n1014), .C1(new_n853), .C2(new_n205), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n324), .B1(new_n792), .B2(new_n206), .C1(new_n798), .C2(new_n795), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n814), .A2(new_n809), .B1(new_n421), .B2(new_n811), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1279), .A2(KEYINPUT122), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n814), .A2(new_n869), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n853), .A2(new_n816), .B1(new_n1281), .B2(KEYINPUT123), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(KEYINPUT123), .B2(new_n1281), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n860), .A2(new_n1241), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n287), .B1(new_n792), .B2(new_n258), .C1(new_n865), .C2(new_n795), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(G50), .B2(new_n1082), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n787), .A2(G128), .B1(new_n799), .B2(G58), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1283), .A2(new_n1284), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1279), .A2(KEYINPUT122), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1280), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n1273), .B1(new_n877), .B2(new_n1290), .C1(new_n1155), .C2(new_n833), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1173), .A2(new_n903), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1164), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1154), .A2(new_n882), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1293), .A2(new_n1175), .B1(new_n1161), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1291), .B1(new_n1295), .B2(new_n775), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1180), .A2(new_n1062), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1182), .A2(new_n1177), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(G381));
  INV_X1    g1100(.A(G390), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n889), .ZN(new_n1302));
  OR2_X1    g1102(.A1(G393), .A2(G396), .ZN(new_n1303));
  NOR4_X1   g1103(.A1(new_n1302), .A2(G387), .A3(G381), .A4(new_n1303), .ZN(new_n1304));
  XOR2_X1   g1104(.A(new_n1304), .B(KEYINPUT124), .Z(new_n1305));
  OR2_X1    g1105(.A1(G375), .A2(G378), .ZN(new_n1306));
  OR2_X1    g1106(.A1(new_n1305), .A2(new_n1306), .ZN(G407));
  OAI211_X1 g1107(.A(G407), .B(G213), .C1(G343), .C2(new_n1306), .ZN(G409));
  AND2_X1   g1108(.A1(new_n691), .A2(G213), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(G2897), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1182), .B2(new_n1177), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n713), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1182), .B2(new_n1177), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1269), .A2(KEYINPUT60), .A3(new_n1295), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT125), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT125), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1313), .A2(new_n1315), .A3(new_n1319), .A4(new_n1316), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(G384), .B1(new_n1321), .B2(new_n1297), .ZN(new_n1322));
  AOI211_X1 g1122(.A(new_n889), .B(new_n1296), .C1(new_n1318), .C2(new_n1320), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1311), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1180), .A2(new_n713), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT60), .B1(new_n1269), .B2(new_n1295), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1319), .B1(new_n1327), .B2(new_n1316), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1320), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1297), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n889), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1321), .A2(G384), .A3(new_n1297), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1331), .A2(new_n1332), .A3(new_n1310), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(G375), .A2(G378), .ZN(new_n1334));
  AND4_X1   g1134(.A1(new_n1188), .A2(new_n1210), .A3(new_n1228), .A4(new_n1257), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1261), .A2(new_n1062), .A3(new_n1262), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1309), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1334), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1324), .A2(new_n1333), .A3(new_n1338), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1334), .A2(new_n1331), .A3(new_n1332), .A4(new_n1337), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(KEYINPUT62), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1343), .A2(new_n1344), .A3(new_n1334), .A4(new_n1337), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1339), .A2(new_n1341), .A3(new_n1342), .A4(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(G387), .A2(new_n1301), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(G393), .B(new_n848), .ZN(new_n1348));
  OAI211_X1 g1148(.A(G390), .B(new_n1036), .C1(new_n1063), .C2(new_n1078), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1347), .A2(new_n1348), .A3(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1348), .B1(new_n1347), .B2(new_n1349), .ZN(new_n1351));
  OR2_X1    g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1346), .A2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT126), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1339), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT63), .ZN(new_n1356));
  OR2_X1    g1156(.A1(new_n1340), .A2(new_n1356), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1342), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1359), .B1(new_n1340), .B2(new_n1356), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1324), .A2(new_n1333), .A3(new_n1338), .A4(KEYINPUT126), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1355), .A2(new_n1357), .A3(new_n1360), .A4(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1353), .A2(new_n1362), .ZN(G405));
  XOR2_X1   g1163(.A(G375), .B(G378), .Z(new_n1364));
  OAI21_X1  g1164(.A(KEYINPUT127), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT127), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1352), .B1(new_n1343), .B2(new_n1367), .ZN(new_n1368));
  NOR4_X1   g1168(.A1(new_n1358), .A2(KEYINPUT127), .A3(new_n1322), .A4(new_n1323), .ZN(new_n1369));
  NOR3_X1   g1169(.A1(new_n1366), .A2(new_n1368), .A3(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1343), .A2(new_n1367), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(new_n1358), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1352), .A2(new_n1343), .A3(new_n1367), .ZN(new_n1373));
  AOI22_X1  g1173(.A1(new_n1372), .A2(new_n1373), .B1(new_n1365), .B2(new_n1364), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1370), .A2(new_n1374), .ZN(G402));
endmodule


