//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G101), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n475), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n474), .A2(G136), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n469), .A2(G2105), .A3(new_n472), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  MUX2_X1   g064(.A(G100), .B(G112), .S(G2105), .Z(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2104), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT70), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n470), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n470), .A2(G102), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n469), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n500), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT71), .B1(new_n500), .B2(new_n501), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(new_n470), .A3(G138), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n478), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n469), .A2(G138), .A3(new_n470), .A4(new_n472), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT4), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n502), .A2(new_n503), .A3(new_n508), .ZN(G164));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT72), .B(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT73), .B(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n516), .A2(new_n517), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT75), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n523), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n512), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n515), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n523), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n516), .A2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n515), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(new_n511), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n538), .A2(new_n539), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(G43), .A2(new_n523), .B1(new_n516), .B2(G81), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT76), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n515), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(new_n511), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND3_X1  g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  OR2_X1    g135(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(G91), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT78), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n531), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n523), .A2(new_n567), .A3(G53), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n515), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n566), .A2(new_n568), .B1(G651), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n561), .A2(new_n573), .A3(G91), .A4(new_n562), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n564), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(G299));
  OR2_X1    g152(.A1(new_n533), .A2(new_n536), .ZN(G286));
  NAND3_X1  g153(.A1(new_n561), .A2(G87), .A3(new_n562), .ZN(new_n579));
  INV_X1    g154(.A(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n515), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n523), .A2(G49), .B1(G651), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT80), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n579), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  NAND3_X1  g163(.A1(new_n561), .A2(G86), .A3(new_n562), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n515), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n523), .A2(G48), .B1(new_n511), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n523), .A2(G47), .ZN(new_n595));
  INV_X1    g170(.A(new_n516), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT81), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n515), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n511), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G290));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G301), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n561), .A2(new_n562), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n523), .B(KEYINPUT82), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n515), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n613), .A2(G54), .B1(G651), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n606), .B1(new_n619), .B2(new_n605), .ZN(G284));
  XNOR2_X1  g195(.A(G284), .B(KEYINPUT83), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n605), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(new_n605), .B2(G168), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n552), .A2(new_n605), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n625), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT84), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n629), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g206(.A1(new_n482), .A2(new_n472), .A3(new_n477), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  MUX2_X1   g210(.A(G99), .B(G111), .S(G2105), .Z(new_n636));
  AOI22_X1  g211(.A1(new_n488), .A2(G123), .B1(G2104), .B2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n473), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2427), .ZN(new_n646));
  INV_X1    g221(.A(G2430), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(KEYINPUT17), .ZN(new_n666));
  INV_X1    g241(.A(new_n660), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n667), .A2(new_n663), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n660), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n671));
  INV_X1    g246(.A(new_n662), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n663), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n671), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n640), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n683), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  AOI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n680), .C2(new_n684), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT88), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT89), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n692), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G16), .A2(G19), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n553), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1341), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(G171), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G5), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1961), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G32), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT26), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  AOI22_X1  g286(.A1(G105), .A2(new_n482), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G141), .ZN(new_n713));
  INV_X1    g288(.A(G129), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n712), .B1(new_n473), .B2(new_n713), .C1(new_n714), .C2(new_n487), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n707), .B1(new_n715), .B2(G29), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT27), .B(G1996), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n703), .A2(new_n704), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(new_n717), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n705), .A2(new_n718), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT99), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n639), .A2(new_n706), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT30), .B(G28), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n723), .B(new_n724), .C1(new_n706), .C2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NOR2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n706), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n484), .B2(new_n706), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n726), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n701), .A2(G21), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G168), .B2(new_n701), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1966), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n721), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2078), .ZN(new_n739));
  NAND2_X1  g314(.A1(G164), .A2(G29), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G27), .B2(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n706), .A2(G26), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT28), .Z(new_n743));
  MUX2_X1   g318(.A(G104), .B(G116), .S(G2105), .Z(new_n744));
  AOI22_X1  g319(.A1(new_n488), .A2(G128), .B1(G2104), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n474), .A2(G140), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n745), .A2(KEYINPUT95), .A3(new_n746), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n743), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT96), .B(G2067), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n738), .B1(new_n739), .B2(new_n741), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n619), .B2(G16), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n700), .B(new_n754), .C1(G1348), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G35), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G162), .B2(G29), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT29), .Z(new_n760));
  INV_X1    g335(.A(G2090), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT100), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  INV_X1    g339(.A(new_n756), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(G299), .A2(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n701), .A2(G20), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT23), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G1956), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  INV_X1    g349(.A(G139), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n473), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT97), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n472), .A2(new_n477), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n778), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n777), .B1(new_n470), .B2(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G2072), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT98), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n760), .A2(new_n761), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n752), .A2(new_n753), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n741), .A2(new_n739), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n781), .A2(G2072), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n757), .A2(new_n766), .A3(new_n772), .A4(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G6), .B(G305), .S(G16), .Z(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  XOR2_X1   g367(.A(new_n791), .B(new_n792), .Z(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(new_n583), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT33), .B(G1976), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT92), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n796), .B(new_n798), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n701), .A2(G22), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT93), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G303), .B2(G16), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1971), .Z(new_n803));
  NOR3_X1   g378(.A1(new_n793), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n701), .A2(G24), .ZN(new_n808));
  XNOR2_X1  g383(.A(G290), .B(KEYINPUT91), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n701), .ZN(new_n810));
  INV_X1    g385(.A(G1986), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G25), .A2(G29), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n474), .A2(G131), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT90), .ZN(new_n815));
  MUX2_X1   g390(.A(G95), .B(G107), .S(G2105), .Z(new_n816));
  AOI22_X1  g391(.A1(new_n488), .A2(G119), .B1(G2104), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n813), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n806), .A2(new_n807), .A3(new_n812), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n790), .B1(new_n824), .B2(new_n825), .ZN(G311));
  INV_X1    g401(.A(new_n790), .ZN(new_n827));
  INV_X1    g402(.A(new_n825), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n823), .ZN(G150));
  NAND2_X1  g404(.A1(new_n523), .A2(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n596), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n515), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n511), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  INV_X1    g417(.A(new_n839), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n552), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n839), .B1(new_n547), .B2(new_n551), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n619), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n840), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n842), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT102), .ZN(G145));
  MUX2_X1   g428(.A(G106), .B(G118), .S(G2105), .Z(new_n854));
  AOI22_X1  g429(.A1(new_n488), .A2(G130), .B1(G2104), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n474), .A2(G142), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n633), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n818), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n751), .B(new_n715), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n500), .A2(new_n501), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n508), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n780), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n861), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n639), .B(KEYINPUT103), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n492), .B(new_n484), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n868), .B2(new_n865), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n870), .B(KEYINPUT104), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(G395));
  NOR2_X1   g453(.A1(new_n843), .A2(G868), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n629), .B(new_n846), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g456(.A1(G299), .A2(new_n618), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(G299), .A2(new_n618), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(G299), .A2(new_n618), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(KEYINPUT106), .A3(new_n882), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n883), .B2(new_n884), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n880), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G290), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n583), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n583), .B(KEYINPUT107), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(G290), .ZN(new_n900));
  XNOR2_X1  g475(.A(G305), .B(G166), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n898), .B2(new_n900), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT108), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n898), .A2(new_n900), .ZN(new_n906));
  INV_X1    g481(.A(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n909), .A3(new_n902), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n902), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(KEYINPUT42), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n894), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n879), .B1(new_n915), .B2(G868), .ZN(G295));
  AOI21_X1  g491(.A(new_n879), .B1(new_n915), .B2(G868), .ZN(G331));
  XNOR2_X1  g492(.A(G168), .B(G171), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n844), .B2(new_n845), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT109), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n844), .A2(new_n918), .A3(new_n845), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n923), .B(new_n918), .C1(new_n844), .C2(new_n845), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n891), .A2(new_n892), .A3(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n886), .A2(new_n882), .A3(new_n922), .A4(new_n919), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n911), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n927), .ZN(new_n932));
  INV_X1    g507(.A(new_n911), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(KEYINPUT43), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n921), .B1(KEYINPUT109), .B2(new_n919), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n885), .A2(new_n887), .A3(new_n937), .A4(new_n924), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n922), .A2(new_n919), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n891), .A2(new_n892), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n911), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n936), .B1(new_n930), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT44), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n931), .A2(new_n936), .A3(new_n934), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT110), .B1(new_n930), .B2(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n933), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n929), .A4(new_n928), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n944), .B1(new_n950), .B2(new_n936), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n943), .B1(new_n951), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g527(.A(KEYINPUT111), .B(G1384), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT45), .B1(new_n863), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G40), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n484), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n895), .A2(new_n811), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT112), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n811), .B2(new_n895), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n751), .A2(G2067), .ZN(new_n962));
  INV_X1    g537(.A(G2067), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n749), .A2(new_n963), .A3(new_n750), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n818), .A2(new_n820), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n818), .A2(new_n820), .ZN(new_n967));
  INV_X1    g542(.A(G1996), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n715), .B(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n957), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n972), .B(new_n973), .C1(new_n508), .C2(new_n862), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT113), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n503), .A2(new_n508), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n500), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n975), .B1(new_n978), .B2(new_n972), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT113), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n956), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT114), .B1(new_n981), .B2(G2090), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n978), .A2(KEYINPUT45), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n863), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n956), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(G1971), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n980), .A2(new_n956), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n988), .A2(new_n989), .A3(new_n761), .A4(new_n979), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n982), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(G303), .A2(G8), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT115), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n992), .B2(new_n993), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(G8), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n508), .A2(new_n862), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(G1384), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n956), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n584), .A4(new_n586), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT116), .B1(new_n795), .B2(G1976), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1006), .A2(new_n1007), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n584), .A2(new_n1005), .A3(new_n586), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(new_n1008), .A3(new_n1007), .A4(new_n1004), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n589), .A2(new_n1012), .A3(new_n593), .ZN(new_n1013));
  INV_X1    g588(.A(new_n593), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n516), .A2(G86), .ZN(new_n1015));
  OAI21_X1  g590(.A(G1981), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1013), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1004), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1011), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1009), .A2(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n999), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1001), .A2(KEYINPUT50), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(KEYINPUT50), .B2(new_n978), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n956), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n987), .B1(G2090), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n998), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n983), .A2(new_n985), .A3(G2078), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(KEYINPUT53), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n739), .A2(KEYINPUT53), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT71), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n862), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n1039));
  INV_X1    g614(.A(new_n506), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n977), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1036), .B1(new_n1042), .B2(new_n973), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1036), .B(new_n973), .C1(new_n508), .C2(new_n862), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n956), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1034), .B1(new_n1035), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1961), .B1(new_n988), .B2(new_n979), .ZN(new_n1048));
  OAI21_X1  g623(.A(G171), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G286), .A2(G8), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT121), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n1055));
  INV_X1    g630(.A(G1966), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1046), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n979), .A2(new_n731), .A3(new_n956), .A4(new_n980), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1059), .B2(G8), .ZN(new_n1060));
  AOI211_X1 g635(.A(KEYINPUT122), .B(new_n1003), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1054), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1052), .A2(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(G8), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1052), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1003), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT123), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT51), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT124), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1069), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1052), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1068), .B2(KEYINPUT123), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1053), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n1063), .A4(new_n1062), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1071), .A2(KEYINPUT62), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT62), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1050), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1048), .A2(KEYINPUT125), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1033), .A2(KEYINPUT53), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n985), .A2(new_n954), .A3(new_n1035), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1048), .A2(KEYINPUT125), .ZN(new_n1085));
  AOI21_X1  g660(.A(G301), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1047), .A2(G171), .A3(new_n1048), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT54), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(G301), .A3(new_n1085), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1049), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n983), .A2(new_n985), .A3(G1996), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT58), .B(G1341), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1002), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n553), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1095), .A2(KEYINPUT59), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(KEYINPUT59), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n981), .A2(new_n764), .B1(new_n963), .B2(new_n1002), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n618), .A2(KEYINPUT60), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1096), .A2(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1027), .A2(new_n771), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT120), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n986), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n575), .A2(KEYINPUT119), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n575), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1105), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1101), .A2(new_n1108), .A3(new_n1104), .A4(new_n1109), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1098), .A2(new_n618), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1098), .A2(new_n618), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT60), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(KEYINPUT61), .A3(new_n1112), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1100), .A2(new_n1115), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1112), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1121), .A2(new_n1111), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1088), .A2(new_n1091), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1071), .A2(new_n1077), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1032), .B1(new_n1080), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1023), .A2(G8), .A3(new_n998), .A4(new_n991), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1021), .A2(new_n1005), .A3(new_n587), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1013), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1004), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1127), .A2(KEYINPUT117), .A3(new_n1130), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1065), .A2(G286), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1031), .A2(new_n999), .A3(new_n1023), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n991), .A2(G8), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1030), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1024), .A2(KEYINPUT63), .A3(new_n1136), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1135), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT118), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1135), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n971), .B1(new_n1126), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n959), .A2(new_n957), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1150), .A2(KEYINPUT48), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(KEYINPUT48), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n970), .A2(new_n957), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n965), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n957), .B1(new_n1155), .B2(new_n715), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n957), .A2(new_n1157), .A3(KEYINPUT46), .A4(new_n968), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n957), .B(new_n968), .C1(new_n1157), .C2(KEYINPUT46), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT46), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1159), .B1(KEYINPUT126), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1156), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n965), .A2(new_n969), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n964), .B1(new_n1164), .B2(new_n967), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n957), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1154), .A2(new_n1163), .A3(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT127), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1149), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g744(.A1(new_n935), .A2(new_n942), .ZN(new_n1171));
  NOR3_X1   g745(.A1(G227), .A2(new_n463), .A3(G401), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n696), .A2(new_n1172), .ZN(new_n1173));
  NOR3_X1   g747(.A1(new_n872), .A2(new_n1171), .A3(new_n1173), .ZN(G308));
  INV_X1    g748(.A(G308), .ZN(G225));
endmodule


