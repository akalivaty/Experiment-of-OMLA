//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT69), .A2(G237), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT69), .A2(G237), .ZN(new_n191));
  OAI211_X1 g005(.A(G210), .B(new_n188), .C1(new_n190), .C2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT27), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT69), .B(G237), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT27), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G210), .A4(new_n188), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G101), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n193), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n193), .B2(new_n196), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n203), .A2(new_n204), .B1(KEYINPUT2), .B2(G113), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G116), .ZN(new_n207));
  INV_X1    g021(.A(G116), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n210), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT2), .A2(G113), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT2), .A2(G113), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n216), .B2(new_n202), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT30), .ZN(new_n220));
  XNOR2_X1  g034(.A(G134), .B(G137), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  INV_X1    g038(.A(G134), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT11), .A3(G134), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(G137), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n226), .A2(new_n228), .A3(new_n222), .A4(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n225), .A2(G137), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n227), .A2(G134), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n231), .B(G131), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n223), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G143), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n241), .B(KEYINPUT1), .C1(new_n238), .C2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G128), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n241), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n240), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  AND4_X1   g060(.A1(new_n246), .A2(new_n237), .A3(new_n239), .A4(G128), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G131), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n230), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n237), .A2(new_n239), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT0), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT65), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(KEYINPUT0), .B2(G128), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n257), .A2(new_n259), .B1(KEYINPUT0), .B2(G128), .ZN(new_n260));
  INV_X1    g074(.A(new_n240), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n254), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n235), .A2(new_n249), .B1(new_n252), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n220), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n252), .A2(new_n262), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT1), .B1(new_n238), .B2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT67), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(G128), .A3(new_n242), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n247), .B1(new_n269), .B2(new_n240), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n223), .A2(new_n230), .A3(new_n234), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n266), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n219), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n266), .B(new_n219), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n201), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n235), .A2(new_n249), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n219), .B1(new_n279), .B2(new_n266), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n278), .B(KEYINPUT28), .C1(new_n276), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n211), .A2(new_n218), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n270), .A2(new_n271), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n257), .A2(new_n259), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n253), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n240), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n287), .A2(new_n254), .B1(new_n230), .B2(new_n251), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n283), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n282), .B1(new_n289), .B2(new_n275), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n275), .A2(new_n282), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n281), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n187), .B(new_n277), .C1(new_n294), .C2(new_n201), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n289), .A2(new_n296), .A3(new_n275), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n280), .A2(KEYINPUT73), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(KEYINPUT28), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n297), .A2(KEYINPUT74), .A3(KEYINPUT28), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n291), .A2(KEYINPUT29), .A3(new_n200), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n295), .B1(new_n305), .B2(KEYINPUT75), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n307));
  AOI211_X1 g121(.A(new_n307), .B(G902), .C1(new_n303), .C2(new_n304), .ZN(new_n308));
  OAI21_X1  g122(.A(G472), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT31), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n275), .A2(KEYINPUT70), .A3(new_n200), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT70), .B1(new_n275), .B2(new_n200), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n311), .B1(new_n314), .B2(new_n274), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n275), .A2(new_n200), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n275), .A2(KEYINPUT70), .A3(new_n200), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n263), .A2(new_n264), .A3(new_n220), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT30), .B1(new_n272), .B2(KEYINPUT64), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n283), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n323), .A3(KEYINPUT31), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n201), .A2(new_n294), .B1(new_n315), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(G472), .A2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n310), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT32), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n315), .A2(new_n324), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n281), .B(new_n201), .C1(new_n290), .C2(new_n292), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT72), .A3(new_n326), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n325), .A2(new_n329), .A3(new_n327), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n309), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n256), .A2(G119), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n206), .A2(G128), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n256), .A2(KEYINPUT23), .A3(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n338), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT24), .B(G110), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n343), .A2(G110), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G125), .ZN(new_n350));
  INV_X1    g164(.A(G125), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G140), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT16), .ZN(new_n353));
  OR3_X1    g167(.A1(new_n351), .A2(KEYINPUT16), .A3(G140), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(G146), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(G146), .B1(new_n353), .B2(new_n354), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n348), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n344), .A2(new_n346), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT76), .ZN(new_n360));
  INV_X1    g174(.A(G110), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n340), .A2(new_n342), .A3(new_n361), .A4(new_n341), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n344), .A2(new_n346), .A3(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n360), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n350), .A2(new_n352), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G125), .B(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT77), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n370), .A3(new_n236), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n355), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n365), .A2(KEYINPUT78), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n371), .A2(new_n355), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n360), .A2(new_n362), .A3(new_n364), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n358), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G137), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n358), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT78), .B1(new_n365), .B2(new_n372), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n375), .A2(new_n374), .A3(new_n376), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n381), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n382), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT25), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n382), .A2(new_n389), .A3(KEYINPUT25), .A4(new_n383), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G217), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(G234), .B2(new_n383), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n387), .A2(new_n388), .ZN(new_n399));
  AOI211_X1 g213(.A(new_n381), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n396), .A2(G902), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n397), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n396), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n392), .B2(new_n393), .ZN(new_n406));
  INV_X1    g220(.A(new_n403), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT79), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G104), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT3), .B1(new_n411), .B2(G107), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n413));
  INV_X1    g227(.A(G107), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(G104), .ZN(new_n415));
  INV_X1    g229(.A(G101), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(G107), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n412), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n411), .A2(G107), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n414), .A2(G104), .ZN(new_n420));
  OAI21_X1  g234(.A(G101), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT83), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n249), .A2(new_n423), .A3(KEYINPUT10), .A4(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT10), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n267), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n237), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(G128), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n247), .B1(new_n431), .B2(new_n240), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n427), .B1(new_n432), .B2(new_n422), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n251), .A2(new_n230), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n412), .A2(new_n415), .A3(new_n417), .ZN(new_n435));
  AND2_X1   g249(.A1(KEYINPUT81), .A2(G101), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT4), .A3(new_n418), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n435), .A2(KEYINPUT81), .A3(new_n439), .A4(G101), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n262), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n426), .A2(new_n433), .A3(new_n434), .A4(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n245), .A2(new_n422), .A3(new_n248), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n432), .B2(new_n422), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT12), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(new_n434), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n444), .A2(new_n447), .A3(new_n252), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n252), .B2(new_n444), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n442), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G140), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n188), .A2(G227), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n451), .B(new_n452), .Z(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n442), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n426), .A2(new_n433), .A3(new_n441), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n252), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n450), .A2(new_n453), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G469), .B1(new_n458), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(G469), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n448), .A2(new_n449), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n442), .A2(new_n454), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n454), .B1(new_n457), .B2(new_n442), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n460), .B(new_n383), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT9), .B(G234), .ZN(new_n467));
  OAI21_X1  g281(.A(G221), .B1(new_n467), .B2(G902), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n468), .B(KEYINPUT80), .Z(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G210), .B1(G237), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n283), .A2(new_n438), .A3(new_n440), .ZN(new_n473));
  INV_X1    g287(.A(G113), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n208), .A2(G119), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT5), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT5), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n217), .A2(new_n212), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n423), .A2(new_n479), .A3(new_n425), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G122), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n473), .A2(new_n480), .A3(new_n482), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n245), .A2(new_n248), .A3(new_n351), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n351), .B2(new_n262), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n188), .A2(G224), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT85), .Z(new_n490));
  XNOR2_X1  g304(.A(new_n488), .B(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n481), .A2(new_n492), .A3(new_n483), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n486), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n487), .B(KEYINPUT87), .C1(new_n351), .C2(new_n262), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(KEYINPUT7), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n495), .B(new_n496), .C1(KEYINPUT87), .C2(new_n487), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n489), .A2(KEYINPUT88), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n489), .A2(KEYINPUT88), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(KEYINPUT7), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n488), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n418), .A2(new_n421), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n479), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n482), .B(KEYINPUT8), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n479), .B2(new_n503), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n497), .A2(new_n501), .A3(new_n485), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n383), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n472), .B1(new_n494), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n485), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n488), .A2(new_n500), .B1(new_n504), .B2(new_n506), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n513), .B2(new_n497), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n486), .A2(new_n491), .A3(new_n493), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n471), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G952), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(G953), .ZN(new_n519));
  NAND2_X1  g333(.A1(G234), .A2(G237), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(G902), .A3(G953), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT21), .B(G898), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(G214), .B1(G237), .B2(G902), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n466), .A2(new_n470), .A3(new_n517), .A4(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(G214), .B(new_n188), .C1(new_n190), .C2(new_n191), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n238), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n194), .A2(G143), .A3(G214), .A4(new_n188), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G131), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT89), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT89), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n538), .A3(G131), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n532), .A2(new_n533), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n222), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n356), .A2(new_n357), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n538), .B1(new_n534), .B2(G131), .ZN(new_n544));
  AOI211_X1 g358(.A(KEYINPUT89), .B(new_n222), .C1(new_n532), .C2(new_n533), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT17), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G113), .B(G122), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n411), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT18), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n540), .B1(new_n550), .B2(new_n222), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n534), .A2(KEYINPUT18), .A3(G131), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n371), .B1(new_n236), .B2(new_n369), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n547), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n549), .B1(new_n547), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n383), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  XNOR2_X1  g372(.A(G116), .B(G122), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(new_n414), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n238), .A2(G128), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT13), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n256), .A2(G143), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  OAI21_X1  g380(.A(G134), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(new_n564), .A3(new_n225), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n560), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n188), .A2(G217), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n467), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n561), .A2(new_n564), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G134), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n575), .A2(new_n568), .B1(new_n414), .B2(new_n559), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n208), .A2(KEYINPUT14), .A3(G122), .ZN(new_n577));
  XOR2_X1   g391(.A(G116), .B(G122), .Z(new_n578));
  OAI211_X1 g392(.A(G107), .B(new_n577), .C1(new_n578), .C2(KEYINPUT14), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n569), .A2(new_n573), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n573), .B1(new_n569), .B2(new_n580), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n383), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G478), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n585), .A2(KEYINPUT15), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n584), .B(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT20), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n547), .A2(new_n549), .A3(new_n554), .ZN(new_n589));
  INV_X1    g403(.A(new_n549), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT90), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n368), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n367), .B1(new_n593), .B2(KEYINPUT90), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n592), .A2(new_n593), .B1(new_n369), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n355), .B1(new_n595), .B2(G146), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n544), .A2(new_n545), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n597), .B2(new_n541), .ZN(new_n598));
  INV_X1    g412(.A(new_n554), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n590), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n589), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(G475), .A2(G902), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n588), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n602), .ZN(new_n604));
  AOI211_X1 g418(.A(KEYINPUT20), .B(new_n604), .C1(new_n589), .C2(new_n600), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n558), .B(new_n587), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n530), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n337), .A2(new_n410), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  OAI21_X1  g423(.A(G472), .B1(new_n325), .B2(G902), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n328), .A2(new_n610), .A3(new_n333), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n409), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n469), .B1(new_n459), .B2(new_n465), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT92), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n471), .B1(new_n514), .B2(new_n515), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n528), .B1(new_n616), .B2(KEYINPUT93), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n510), .A2(new_n618), .A3(new_n516), .ZN(new_n619));
  INV_X1    g433(.A(new_n526), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n601), .A2(new_n602), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT20), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n601), .A2(new_n588), .A3(new_n602), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n623), .A2(new_n624), .B1(G475), .B2(new_n557), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n569), .A2(new_n580), .ZN(new_n627));
  INV_X1    g441(.A(new_n573), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n581), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n569), .A2(new_n573), .A3(new_n580), .A4(KEYINPUT94), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT95), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n626), .B1(new_n582), .B2(new_n583), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT95), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n629), .A2(new_n631), .A3(new_n636), .A4(new_n632), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n585), .A2(G902), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n634), .A2(new_n635), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n637), .A2(new_n635), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n642), .A2(KEYINPUT96), .A3(new_n634), .A4(new_n638), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT97), .B(G478), .Z(new_n644));
  AOI22_X1  g458(.A1(new_n641), .A2(new_n643), .B1(new_n584), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT98), .B1(new_n625), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n558), .B1(new_n603), .B2(new_n605), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n641), .A2(new_n643), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n584), .A2(new_n644), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n621), .B1(new_n646), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n615), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  INV_X1    g470(.A(new_n587), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n625), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n621), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n615), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  OAI21_X1  g476(.A(new_n378), .B1(KEYINPUT36), .B2(new_n381), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n381), .A2(KEYINPUT36), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n387), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n394), .A2(new_n396), .B1(new_n402), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n530), .A2(new_n606), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n611), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n402), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n397), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(new_n613), .A3(new_n619), .A4(new_n617), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n521), .B1(G900), .B2(new_n523), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n625), .A2(new_n657), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n337), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT99), .B(G128), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G30));
  NOR2_X1   g495(.A1(new_n314), .A2(new_n274), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n297), .A2(new_n201), .A3(new_n298), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n383), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G472), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n334), .A2(new_n336), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n647), .A2(new_n657), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n517), .B(KEYINPUT38), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n527), .A3(new_n667), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n613), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n676), .B(KEYINPUT39), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT100), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n613), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n690), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n238), .ZN(G45));
  NAND3_X1  g519(.A1(new_n647), .A2(new_n650), .A3(new_n676), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n675), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n337), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NOR2_X1   g523(.A1(new_n463), .A2(new_n464), .ZN(new_n710));
  OAI21_X1  g524(.A(G469), .B1(new_n710), .B2(G902), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n470), .A3(new_n465), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n409), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n653), .A2(new_n337), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND3_X1  g530(.A1(new_n337), .A2(new_n659), .A3(new_n713), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT102), .B(G116), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G18));
  NAND2_X1  g533(.A1(new_n617), .A2(new_n619), .ZN(new_n720));
  NOR4_X1   g534(.A1(new_n720), .A2(new_n712), .A3(new_n667), .A4(new_n526), .ZN(new_n721));
  INV_X1    g535(.A(new_n606), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n337), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  AOI21_X1  g538(.A(new_n200), .B1(new_n303), .B2(new_n291), .ZN(new_n725));
  INV_X1    g539(.A(new_n330), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n326), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n406), .A2(new_n407), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n610), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT103), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n610), .A2(new_n727), .A3(new_n731), .A4(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n687), .A2(KEYINPUT104), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n647), .A2(new_n735), .A3(new_n657), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n720), .A2(new_n712), .A3(new_n526), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n733), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n733), .A2(new_n737), .A3(KEYINPUT105), .A4(new_n738), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND3_X1  g558(.A1(new_n610), .A2(new_n674), .A3(new_n727), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n706), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n720), .A2(new_n712), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NAND3_X1  g563(.A1(new_n510), .A2(new_n516), .A3(new_n527), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n510), .A2(new_n516), .A3(KEYINPUT106), .A4(new_n527), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n613), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n754), .A2(new_n706), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT32), .B1(new_n332), .B2(new_n326), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n335), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n309), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT108), .B1(new_n759), .B2(new_n728), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  INV_X1    g575(.A(new_n728), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n761), .B(new_n762), .C1(new_n309), .C2(new_n758), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n756), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n754), .A2(new_n706), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n337), .A2(new_n410), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(KEYINPUT107), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n337), .A2(new_n765), .A3(new_n768), .A4(new_n410), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n755), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n764), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NOR2_X1   g586(.A1(new_n677), .A2(new_n754), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n337), .A2(new_n410), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  NAND2_X1  g589(.A1(new_n752), .A2(new_n753), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n458), .A2(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n458), .A2(KEYINPUT45), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(G469), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(G469), .A2(G902), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT46), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n465), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n780), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n470), .B(new_n692), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n558), .B(KEYINPUT109), .C1(new_n603), .C2(new_n605), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n786), .B(new_n787), .C1(new_n647), .C2(new_n645), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n625), .B(new_n650), .C1(KEYINPUT109), .C2(KEYINPUT43), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n669), .B(new_n667), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n776), .B(new_n785), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n337), .A2(new_n410), .A3(new_n706), .A4(new_n776), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n784), .A2(new_n781), .A3(new_n782), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n469), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT47), .B(new_n470), .C1(new_n783), .C2(new_n784), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n799), .A2(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n800), .A2(new_n799), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n521), .B1(new_n788), .B2(new_n789), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n688), .A2(new_n527), .A3(new_n712), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n733), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n733), .A2(new_n810), .A3(KEYINPUT50), .A4(new_n811), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n711), .A2(new_n465), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(new_n752), .A3(new_n470), .A4(new_n753), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n521), .B(new_n819), .C1(new_n789), .C2(new_n788), .ZN(new_n820));
  INV_X1    g634(.A(new_n745), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n334), .A2(new_n336), .A3(new_n685), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n404), .A2(new_n408), .A3(new_n522), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n647), .A2(new_n650), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT114), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n819), .A2(new_n824), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n686), .A2(new_n828), .A3(new_n826), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n822), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n809), .B1(new_n817), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n825), .A2(KEYINPUT114), .A3(new_n826), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n830), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n834), .A2(new_n835), .B1(new_n821), .B2(new_n820), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(KEYINPUT115), .A3(new_n816), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n818), .A2(new_n469), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n803), .A2(new_n804), .A3(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n733), .A2(new_n810), .A3(new_n752), .A4(new_n753), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n833), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n836), .A2(new_n841), .A3(new_n816), .A4(KEYINPUT51), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n733), .A2(new_n810), .A3(new_n747), .ZN(new_n846));
  INV_X1    g660(.A(new_n825), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n646), .A2(new_n652), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n846), .B(new_n519), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n762), .B1(new_n309), .B2(new_n758), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT108), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT48), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n820), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n820), .B1(new_n763), .B2(new_n760), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT48), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n849), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n845), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT116), .B1(new_n844), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n860), .B(new_n857), .C1(new_n842), .C2(new_n843), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n714), .A2(new_n723), .A3(new_n717), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n741), .B2(new_n742), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n647), .A2(new_n650), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n530), .B1(new_n658), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n612), .A2(new_n867), .B1(new_n668), .B2(new_n669), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n674), .A2(new_n676), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n754), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n337), .A2(new_n722), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n868), .A2(new_n608), .A3(new_n774), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n873));
  INV_X1    g687(.A(new_n754), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n746), .B2(new_n874), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n745), .A2(new_n754), .A3(new_n706), .A4(KEYINPUT112), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n865), .A2(new_n878), .A3(new_n771), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n679), .A2(new_n708), .A3(new_n748), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n667), .A2(new_n613), .A3(new_n676), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n823), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n720), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n734), .A2(new_n883), .A3(new_n736), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT52), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n678), .A2(new_n337), .B1(new_n746), .B2(new_n747), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n737), .A2(new_n883), .A3(new_n823), .A4(new_n881), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(new_n887), .A3(new_n888), .A4(new_n708), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n863), .B1(new_n879), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT113), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n886), .A2(new_n892), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n879), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n894), .A2(new_n895), .B1(new_n897), .B2(KEYINPUT53), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n879), .A2(new_n896), .A3(KEYINPUT113), .A4(new_n863), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT54), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n893), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n865), .A2(new_n878), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT53), .A4(new_n771), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n863), .B1(new_n879), .B2(new_n896), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n862), .A2(KEYINPUT117), .A3(new_n900), .A4(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n894), .A2(new_n895), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n897), .A2(KEYINPUT53), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n899), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n906), .B1(new_n911), .B2(new_n904), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n836), .A2(new_n816), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n913), .A2(new_n809), .B1(new_n839), .B2(new_n840), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT51), .B1(new_n914), .B2(new_n837), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n860), .B1(new_n915), .B2(new_n857), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n844), .A2(KEYINPUT116), .A3(new_n858), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n908), .B1(new_n912), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n518), .A2(new_n188), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n907), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n818), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(KEYINPUT49), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(KEYINPUT49), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n762), .A2(new_n469), .A3(new_n528), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n647), .A2(new_n645), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OR4_X1    g742(.A1(new_n823), .A2(new_n926), .A3(new_n688), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n921), .A2(new_n929), .ZN(G75));
  NOR2_X1   g744(.A1(new_n188), .A2(G952), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT120), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n903), .A2(new_n905), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n934), .A2(G210), .A3(G902), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n486), .A2(new_n493), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n491), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n494), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(KEYINPUT118), .ZN(new_n942));
  OR3_X1    g756(.A1(new_n935), .A2(KEYINPUT56), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT119), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n939), .B1(new_n935), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n933), .B1(new_n943), .B2(new_n946), .ZN(G51));
  NAND2_X1  g761(.A1(new_n934), .A2(KEYINPUT54), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n906), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n780), .B(KEYINPUT57), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n710), .B(KEYINPUT121), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n934), .ZN(new_n954));
  OR3_X1    g768(.A1(new_n954), .A2(new_n383), .A3(new_n779), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n931), .B1(new_n953), .B2(new_n955), .ZN(G54));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n383), .ZN(new_n957));
  AND2_X1   g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n601), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n959), .A2(KEYINPUT122), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT122), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n957), .A2(new_n601), .A3(new_n958), .ZN(new_n963));
  INV_X1    g777(.A(new_n931), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n961), .A2(new_n962), .A3(new_n965), .ZN(G60));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n642), .A2(new_n634), .ZN(new_n968));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT59), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n912), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n968), .A2(new_n971), .ZN(new_n973));
  INV_X1    g787(.A(new_n906), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n904), .B1(new_n903), .B2(new_n905), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n932), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n967), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n933), .B1(new_n949), .B2(new_n973), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n970), .B1(new_n900), .B2(new_n906), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n979), .B(KEYINPUT123), .C1(new_n980), .C2(new_n968), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(G63));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT60), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n903), .B2(new_n905), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n932), .B1(new_n986), .B2(new_n401), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  INV_X1    g804(.A(new_n985), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n934), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n401), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n933), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n666), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n995), .B(new_n985), .C1(new_n903), .C2(new_n905), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n987), .A2(KEYINPUT125), .A3(new_n996), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n989), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT61), .B1(new_n994), .B2(KEYINPUT124), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT125), .B1(new_n987), .B2(new_n996), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n994), .A2(new_n990), .A3(new_n997), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1000), .A2(new_n1004), .ZN(G66));
  INV_X1    g819(.A(new_n525), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n188), .B1(new_n1006), .B2(G224), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n865), .A2(new_n608), .A3(new_n868), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n188), .ZN(new_n1009));
  INV_X1    g823(.A(G898), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n936), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1009), .B(new_n1011), .ZN(G69));
  AOI22_X1  g826(.A1(new_n795), .A2(new_n796), .B1(new_n805), .B2(new_n806), .ZN(new_n1013));
  INV_X1    g827(.A(new_n880), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n702), .A2(new_n703), .A3(new_n1014), .ZN(new_n1015));
  OR2_X1    g829(.A1(new_n1015), .A2(KEYINPUT62), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(KEYINPUT62), .ZN(new_n1017));
  INV_X1    g831(.A(new_n697), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n776), .B1(new_n658), .B2(new_n866), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1018), .A2(new_n337), .A3(new_n410), .A4(new_n1019), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n188), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n265), .A2(new_n273), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(new_n595), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n785), .A2(new_n884), .ZN(new_n1025));
  AOI21_X1  g839(.A(KEYINPUT127), .B1(new_n1025), .B2(new_n851), .ZN(new_n1026));
  INV_X1    g840(.A(new_n774), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n1026), .A2(new_n1027), .A3(new_n880), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1025), .A2(new_n851), .A3(KEYINPUT127), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1013), .A2(new_n188), .A3(new_n771), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1024), .B1(G900), .B2(G953), .ZN(new_n1032));
  AOI22_X1  g846(.A1(new_n1022), .A2(new_n1024), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT126), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1033), .B(new_n1036), .ZN(G72));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT63), .Z(new_n1039));
  NAND3_X1  g853(.A1(new_n1013), .A2(new_n771), .A3(new_n1030), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1039), .B1(new_n1040), .B2(new_n1008), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n274), .A2(new_n276), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1041), .A2(new_n201), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1039), .B1(new_n1021), .B2(new_n1008), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1042), .A2(new_n201), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1043), .A2(new_n1046), .A3(new_n964), .ZN(new_n1047));
  INV_X1    g861(.A(new_n277), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1039), .B1(new_n1048), .B2(new_n682), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n911), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1047), .A2(new_n1050), .ZN(G57));
endmodule


