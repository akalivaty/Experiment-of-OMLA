

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U556 ( .A1(n809), .A2(n686), .ZN(n732) );
  INV_X1 U557 ( .A(n732), .ZN(n704) );
  NAND2_X1 U558 ( .A1(n748), .A2(n747), .ZN(n767) );
  NOR2_X2 U559 ( .A1(n542), .A2(n541), .ZN(G160) );
  OR2_X1 U560 ( .A1(n815), .A2(n814), .ZN(n522) );
  XNOR2_X1 U561 ( .A(n690), .B(KEYINPUT93), .ZN(n691) );
  XNOR2_X1 U562 ( .A(n692), .B(n691), .ZN(n694) );
  AND2_X1 U563 ( .A1(n744), .A2(n722), .ZN(n723) );
  XNOR2_X1 U564 ( .A(n741), .B(KEYINPUT32), .ZN(n748) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n809) );
  NOR2_X2 U566 ( .A1(n526), .A2(n527), .ZN(n883) );
  NAND2_X1 U567 ( .A1(n816), .A2(n522), .ZN(n817) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XOR2_X1 U569 ( .A(KEYINPUT68), .B(n523), .Z(n524) );
  XNOR2_X2 U570 ( .A(KEYINPUT17), .B(n524), .ZN(n880) );
  NAND2_X1 U571 ( .A1(n880), .A2(G138), .ZN(n525) );
  XNOR2_X1 U572 ( .A(n525), .B(KEYINPUT84), .ZN(n533) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  AND2_X1 U574 ( .A1(n885), .A2(G114), .ZN(n531) );
  XOR2_X1 U575 ( .A(G2104), .B(KEYINPUT65), .Z(n526) );
  INV_X1 U576 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U577 ( .A1(G126), .A2(n883), .ZN(n529) );
  AND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n613) );
  NAND2_X1 U579 ( .A1(G102), .A2(n613), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  AND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(G164) );
  AND2_X1 U583 ( .A1(G125), .A2(n883), .ZN(n534) );
  XNOR2_X1 U584 ( .A(KEYINPUT66), .B(n534), .ZN(n537) );
  NAND2_X1 U585 ( .A1(G101), .A2(n613), .ZN(n535) );
  XNOR2_X1 U586 ( .A(KEYINPUT23), .B(n535), .ZN(n536) );
  NOR2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n539) );
  NAND2_X1 U588 ( .A1(G137), .A2(n880), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U590 ( .A1(G113), .A2(n885), .ZN(n540) );
  XNOR2_X1 U591 ( .A(KEYINPUT67), .B(n540), .ZN(n541) );
  INV_X1 U592 ( .A(G651), .ZN(n547) );
  NOR2_X1 U593 ( .A1(G543), .A2(n547), .ZN(n543) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n543), .Z(n653) );
  NAND2_X1 U595 ( .A1(G64), .A2(n653), .ZN(n546) );
  XOR2_X1 U596 ( .A(KEYINPUT0), .B(G543), .Z(n654) );
  NOR2_X1 U597 ( .A1(G651), .A2(n654), .ZN(n544) );
  XNOR2_X1 U598 ( .A(KEYINPUT64), .B(n544), .ZN(n649) );
  NAND2_X1 U599 ( .A1(G52), .A2(n649), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n553) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n640) );
  NAND2_X1 U602 ( .A1(G90), .A2(n640), .ZN(n549) );
  NOR2_X1 U603 ( .A1(n654), .A2(n547), .ZN(n643) );
  NAND2_X1 U604 ( .A1(G77), .A2(n643), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U606 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  XNOR2_X1 U607 ( .A(KEYINPUT69), .B(n551), .ZN(n552) );
  NOR2_X1 U608 ( .A1(n553), .A2(n552), .ZN(G171) );
  INV_X1 U609 ( .A(G108), .ZN(G238) );
  INV_X1 U610 ( .A(G120), .ZN(G236) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  NAND2_X1 U612 ( .A1(G62), .A2(n653), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G50), .A2(n649), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT80), .B(n556), .Z(n560) );
  NAND2_X1 U616 ( .A1(G88), .A2(n640), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G75), .A2(n643), .ZN(n557) );
  AND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(G303) );
  NAND2_X1 U620 ( .A1(G89), .A2(n640), .ZN(n561) );
  XOR2_X1 U621 ( .A(KEYINPUT75), .B(n561), .Z(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G76), .A2(n643), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U625 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U626 ( .A1(G63), .A2(n653), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G51), .A2(n649), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U631 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(n572) );
  XNOR2_X1 U633 ( .A(KEYINPUT76), .B(n572), .ZN(G286) );
  NAND2_X1 U634 ( .A1(G94), .A2(G452), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT70), .B(n573), .Z(G173) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n574), .B(KEYINPUT10), .ZN(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT72), .B(n575), .ZN(G223) );
  INV_X1 U639 ( .A(G567), .ZN(n680) );
  NOR2_X1 U640 ( .A1(G223), .A2(n680), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U642 ( .A(G860), .ZN(n606) );
  NAND2_X1 U643 ( .A1(G56), .A2(n653), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(n577), .Z(n583) );
  NAND2_X1 U645 ( .A1(n640), .A2(G81), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G68), .A2(n643), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U649 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G43), .A2(n649), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n1010) );
  NOR2_X1 U653 ( .A1(n606), .A2(n1010), .ZN(n586) );
  XNOR2_X1 U654 ( .A(n586), .B(KEYINPUT73), .ZN(G153) );
  INV_X1 U655 ( .A(G171), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U657 ( .A1(G54), .A2(n649), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G66), .A2(n653), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G79), .A2(n643), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n640), .A2(G92), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT74), .B(n589), .Z(n590) );
  NOR2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U665 ( .A(KEYINPUT15), .B(n594), .Z(n1012) );
  INV_X1 U666 ( .A(G868), .ZN(n665) );
  NAND2_X1 U667 ( .A1(n1012), .A2(n665), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G91), .A2(n640), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G78), .A2(n643), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U672 ( .A(KEYINPUT71), .B(n599), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n649), .A2(G53), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G65), .A2(n653), .ZN(n600) );
  AND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(G299) );
  NAND2_X1 U677 ( .A1(G868), .A2(G286), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G299), .A2(n665), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n606), .A2(G559), .ZN(n607) );
  INV_X1 U681 ( .A(n1012), .ZN(n631) );
  NAND2_X1 U682 ( .A1(n607), .A2(n631), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n1010), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n631), .A2(G868), .ZN(n609) );
  NOR2_X1 U686 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G123), .A2(n883), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT18), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G111), .A2(n885), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G99), .A2(n613), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U693 ( .A1(G135), .A2(n880), .ZN(n616) );
  XNOR2_X1 U694 ( .A(KEYINPUT77), .B(n616), .ZN(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U697 ( .A(KEYINPUT78), .B(n621), .Z(n985) );
  XNOR2_X1 U698 ( .A(n985), .B(G2096), .ZN(n623) );
  INV_X1 U699 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G67), .A2(n653), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G93), .A2(n640), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G80), .A2(n643), .ZN(n626) );
  XNOR2_X1 U705 ( .A(KEYINPUT79), .B(n626), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G55), .A2(n649), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n666) );
  NAND2_X1 U709 ( .A1(G559), .A2(n631), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n632), .B(n1010), .ZN(n663) );
  NOR2_X1 U711 ( .A1(G860), .A2(n663), .ZN(n633) );
  XOR2_X1 U712 ( .A(n666), .B(n633), .Z(G145) );
  AND2_X1 U713 ( .A1(n653), .A2(G60), .ZN(n637) );
  NAND2_X1 U714 ( .A1(G85), .A2(n640), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G72), .A2(n643), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U718 ( .A1(G47), .A2(n649), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G61), .A2(n653), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G86), .A2(n640), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U726 ( .A1(G48), .A2(n649), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(G305) );
  NAND2_X1 U728 ( .A1(G651), .A2(G74), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G49), .A2(n649), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n654), .A2(G87), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(G288) );
  INV_X1 U734 ( .A(G299), .ZN(n1020) );
  XNOR2_X1 U735 ( .A(n1020), .B(G303), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n657), .B(n666), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n658), .B(G290), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n659), .B(G305), .ZN(n660) );
  XNOR2_X1 U739 ( .A(KEYINPUT19), .B(n660), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n661), .B(G288), .ZN(n906) );
  XOR2_X1 U741 ( .A(KEYINPUT81), .B(n906), .Z(n662) );
  XNOR2_X1 U742 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n664), .A2(G868), .ZN(n668) );
  NAND2_X1 U744 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U750 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U752 ( .A1(G132), .A2(G82), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n673), .B(KEYINPUT22), .ZN(n674) );
  XNOR2_X1 U754 ( .A(n674), .B(KEYINPUT82), .ZN(n675) );
  NOR2_X1 U755 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G96), .A2(n676), .ZN(n835) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n835), .ZN(n677) );
  XNOR2_X1 U758 ( .A(n677), .B(KEYINPUT83), .ZN(n682) );
  NOR2_X1 U759 ( .A1(G236), .A2(G238), .ZN(n678) );
  NAND2_X1 U760 ( .A1(G69), .A2(n678), .ZN(n679) );
  NOR2_X1 U761 ( .A1(G237), .A2(n679), .ZN(n834) );
  NOR2_X1 U762 ( .A1(n680), .A2(n834), .ZN(n681) );
  NOR2_X1 U763 ( .A1(n682), .A2(n681), .ZN(G319) );
  INV_X1 U764 ( .A(G319), .ZN(n684) );
  NAND2_X1 U765 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U766 ( .A1(n684), .A2(n683), .ZN(n833) );
  NAND2_X1 U767 ( .A1(n833), .A2(G36), .ZN(G176) );
  OR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n813) );
  NAND2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n685) );
  NAND2_X1 U770 ( .A1(n813), .A2(n685), .ZN(n1008) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n808) );
  INV_X1 U772 ( .A(n808), .ZN(n686) );
  INV_X1 U773 ( .A(G1961), .ZN(n950) );
  NAND2_X1 U774 ( .A1(n732), .A2(n950), .ZN(n689) );
  XNOR2_X1 U775 ( .A(G2078), .B(KEYINPUT25), .ZN(n687) );
  XNOR2_X1 U776 ( .A(n687), .B(KEYINPUT92), .ZN(n938) );
  NAND2_X1 U777 ( .A1(n704), .A2(n938), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n725) );
  NAND2_X1 U779 ( .A1(n725), .A2(G171), .ZN(n720) );
  NAND2_X1 U780 ( .A1(G2072), .A2(n704), .ZN(n692) );
  INV_X1 U781 ( .A(KEYINPUT27), .ZN(n690) );
  INV_X1 U782 ( .A(G1956), .ZN(n952) );
  NOR2_X1 U783 ( .A1(n704), .A2(n952), .ZN(n693) );
  NOR2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U785 ( .A1(n697), .A2(n1020), .ZN(n696) );
  XOR2_X1 U786 ( .A(KEYINPUT94), .B(KEYINPUT28), .Z(n695) );
  XNOR2_X1 U787 ( .A(n696), .B(n695), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n697), .A2(n1020), .ZN(n715) );
  XOR2_X1 U789 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n705) );
  NOR2_X1 U790 ( .A1(G1996), .A2(n705), .ZN(n698) );
  NOR2_X1 U791 ( .A1(n698), .A2(n1010), .ZN(n702) );
  NAND2_X1 U792 ( .A1(G1348), .A2(n732), .ZN(n700) );
  NAND2_X1 U793 ( .A1(G2067), .A2(n704), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n711) );
  NAND2_X1 U795 ( .A1(n1012), .A2(n711), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n710) );
  INV_X1 U797 ( .A(G1341), .ZN(n1011) );
  NAND2_X1 U798 ( .A1(n1011), .A2(n705), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n703), .A2(n732), .ZN(n708) );
  AND2_X1 U800 ( .A1(G1996), .A2(n704), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n713) );
  NOR2_X1 U804 ( .A1(n711), .A2(n1012), .ZN(n712) );
  NOR2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U808 ( .A(KEYINPUT29), .B(n718), .Z(n719) );
  NAND2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n730) );
  NAND2_X1 U810 ( .A1(G8), .A2(n732), .ZN(n815) );
  NOR2_X1 U811 ( .A1(n815), .A2(G1966), .ZN(n721) );
  XNOR2_X1 U812 ( .A(n721), .B(KEYINPUT91), .ZN(n744) );
  INV_X1 U813 ( .A(G8), .ZN(n738) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n732), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n738), .A2(n742), .ZN(n722) );
  XOR2_X1 U816 ( .A(KEYINPUT30), .B(n723), .Z(n724) );
  NOR2_X1 U817 ( .A1(G168), .A2(n724), .ZN(n727) );
  NOR2_X1 U818 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U820 ( .A(KEYINPUT31), .B(n728), .Z(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n743) );
  AND2_X1 U822 ( .A1(G286), .A2(G8), .ZN(n731) );
  NAND2_X1 U823 ( .A1(n743), .A2(n731), .ZN(n740) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n732), .ZN(n733) );
  XNOR2_X1 U825 ( .A(n733), .B(KEYINPUT96), .ZN(n735) );
  NOR2_X1 U826 ( .A1(n815), .A2(G1971), .ZN(n734) );
  NOR2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U828 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  AND2_X1 U830 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U831 ( .A1(G8), .A2(n742), .ZN(n746) );
  AND2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n1018) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n749) );
  XOR2_X1 U836 ( .A(n749), .B(KEYINPUT97), .Z(n750) );
  NOR2_X1 U837 ( .A1(n1018), .A2(n750), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n767), .A2(n751), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(KEYINPUT98), .ZN(n754) );
  INV_X1 U840 ( .A(n815), .ZN(n753) );
  AND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n758) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n1015) );
  INV_X1 U843 ( .A(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n753), .A2(n1018), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n760), .A2(n755), .ZN(n756) );
  XNOR2_X1 U846 ( .A(n756), .B(KEYINPUT99), .ZN(n759) );
  AND2_X1 U847 ( .A1(n1015), .A2(n759), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n763) );
  INV_X1 U849 ( .A(n759), .ZN(n761) );
  OR2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n1008), .A2(n764), .ZN(n818) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n765) );
  XNOR2_X1 U854 ( .A(KEYINPUT100), .B(n765), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n766), .A2(G8), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n769), .A2(n815), .ZN(n812) );
  XNOR2_X1 U858 ( .A(G2067), .B(KEYINPUT37), .ZN(n770) );
  XOR2_X1 U859 ( .A(n770), .B(KEYINPUT86), .Z(n805) );
  NAND2_X1 U860 ( .A1(G140), .A2(n880), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n613), .A2(G104), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U863 ( .A(KEYINPUT34), .B(n773), .ZN(n778) );
  NAND2_X1 U864 ( .A1(G128), .A2(n883), .ZN(n775) );
  NAND2_X1 U865 ( .A1(G116), .A2(n885), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U867 ( .A(KEYINPUT35), .B(n776), .Z(n777) );
  NOR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U869 ( .A(KEYINPUT36), .B(n779), .Z(n897) );
  NOR2_X1 U870 ( .A1(n805), .A2(n897), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n780), .B(KEYINPUT103), .ZN(n996) );
  NAND2_X1 U872 ( .A1(n613), .A2(G105), .ZN(n781) );
  XNOR2_X1 U873 ( .A(n781), .B(KEYINPUT38), .ZN(n783) );
  NAND2_X1 U874 ( .A1(G129), .A2(n883), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G117), .A2(n885), .ZN(n784) );
  XNOR2_X1 U877 ( .A(KEYINPUT89), .B(n784), .ZN(n785) );
  NOR2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U879 ( .A(n787), .B(KEYINPUT90), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G141), .A2(n880), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n898) );
  NOR2_X1 U882 ( .A1(G1996), .A2(n898), .ZN(n790) );
  XOR2_X1 U883 ( .A(KEYINPUT101), .B(n790), .Z(n992) );
  XNOR2_X1 U884 ( .A(KEYINPUT87), .B(G1991), .ZN(n929) );
  NAND2_X1 U885 ( .A1(G131), .A2(n880), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n613), .A2(G95), .ZN(n791) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G119), .A2(n883), .ZN(n794) );
  NAND2_X1 U889 ( .A1(G107), .A2(n885), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n878) );
  AND2_X1 U892 ( .A1(n929), .A2(n878), .ZN(n989) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n797) );
  XNOR2_X1 U894 ( .A(KEYINPUT102), .B(n797), .ZN(n798) );
  NOR2_X1 U895 ( .A1(n989), .A2(n798), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n878), .A2(n929), .ZN(n799) );
  XOR2_X1 U897 ( .A(KEYINPUT88), .B(n799), .Z(n801) );
  NAND2_X1 U898 ( .A1(G1996), .A2(n898), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n801), .A2(n800), .ZN(n821) );
  NOR2_X1 U900 ( .A1(n802), .A2(n821), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n992), .A2(n803), .ZN(n804) );
  XNOR2_X1 U902 ( .A(n804), .B(KEYINPUT39), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n805), .A2(n897), .ZN(n820) );
  NAND2_X1 U904 ( .A1(n806), .A2(n820), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n996), .A2(n807), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U907 ( .A(KEYINPUT85), .B(n810), .Z(n823) );
  NAND2_X1 U908 ( .A1(n811), .A2(n823), .ZN(n819) );
  AND2_X1 U909 ( .A1(n812), .A2(n819), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n813), .B(KEYINPUT24), .ZN(n814) );
  OR2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n828) );
  INV_X1 U912 ( .A(n819), .ZN(n826) );
  INV_X1 U913 ( .A(n820), .ZN(n822) );
  NOR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n987) );
  XOR2_X1 U915 ( .A(G1986), .B(G290), .Z(n1005) );
  NAND2_X1 U916 ( .A1(n987), .A2(n1005), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  OR2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n827) );
  AND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U920 ( .A(KEYINPUT40), .B(n829), .ZN(G329) );
  INV_X1 U921 ( .A(G223), .ZN(n830) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U924 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U927 ( .A(n834), .ZN(n836) );
  NOR2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G325) );
  XNOR2_X1 U929 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U931 ( .A(G132), .ZN(G219) );
  INV_X1 U932 ( .A(G82), .ZN(G220) );
  INV_X1 U933 ( .A(G303), .ZN(G166) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n838) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n840) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U940 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1961), .B(G1966), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n856) );
  XOR2_X1 U946 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1981), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1956), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U953 ( .A(KEYINPUT110), .B(G2474), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n883), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n857), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U958 ( .A1(G112), .A2(n885), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G100), .A2(n613), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G136), .A2(n880), .ZN(n860) );
  XNOR2_X1 U962 ( .A(KEYINPUT111), .B(n860), .ZN(n861) );
  NOR2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(KEYINPUT112), .B(n865), .Z(G162) );
  XOR2_X1 U966 ( .A(KEYINPUT117), .B(KEYINPUT113), .Z(n867) );
  XNOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G130), .A2(n883), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G118), .A2(n885), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G106), .A2(n613), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G142), .A2(n880), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(n872), .B(KEYINPUT45), .Z(n873) );
  NOR2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(n876), .B(n875), .Z(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n894) );
  XNOR2_X1 U979 ( .A(G160), .B(G164), .ZN(n892) );
  NAND2_X1 U980 ( .A1(n613), .A2(G103), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n879), .B(KEYINPUT114), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n891) );
  NAND2_X1 U984 ( .A1(n883), .A2(G127), .ZN(n884) );
  XOR2_X1 U985 ( .A(KEYINPUT115), .B(n884), .Z(n887) );
  NAND2_X1 U986 ( .A1(n885), .A2(G115), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT116), .B(n888), .Z(n889) );
  XNOR2_X1 U989 ( .A(KEYINPUT47), .B(n889), .ZN(n890) );
  NOR2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n979) );
  XNOR2_X1 U991 ( .A(n892), .B(n979), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n895), .B(G162), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n896), .B(n985), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U997 ( .A1(G37), .A2(n901), .ZN(G395) );
  XOR2_X1 U998 ( .A(n1012), .B(n1010), .Z(n902) );
  XNOR2_X1 U999 ( .A(G286), .B(n902), .ZN(n908) );
  XOR2_X1 U1000 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n904) );
  XNOR2_X1 U1001 ( .A(G171), .B(KEYINPUT118), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1003 ( .A(n906), .B(n905), .Z(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1006 ( .A(G2451), .B(KEYINPUT106), .Z(n911) );
  XNOR2_X1 U1007 ( .A(G2443), .B(G2446), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1009 ( .A(G2435), .B(KEYINPUT105), .Z(n913) );
  XNOR2_X1 U1010 ( .A(G2438), .B(G2454), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1012 ( .A(n915), .B(n914), .Z(n917) );
  XNOR2_X1 U1013 ( .A(G2427), .B(KEYINPUT104), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n917), .B(n916), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(G1348), .B(G2430), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n918), .B(n1011), .ZN(n919) );
  XOR2_X1 U1017 ( .A(n920), .B(n919), .Z(n921) );
  NAND2_X1 U1018 ( .A1(G14), .A2(n921), .ZN(n927) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G69), .ZN(G235) );
  INV_X1 U1027 ( .A(G96), .ZN(G221) );
  INV_X1 U1028 ( .A(n927), .ZN(G401) );
  XNOR2_X1 U1029 ( .A(G2090), .B(G35), .ZN(n943) );
  XNOR2_X1 U1030 ( .A(G32), .B(G1996), .ZN(n928) );
  XNOR2_X1 U1031 ( .A(n928), .B(KEYINPUT123), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(G2067), .B(G26), .ZN(n931) );
  XOR2_X1 U1033 ( .A(G25), .B(n929), .Z(n930) );
  NOR2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1035 ( .A1(G28), .A2(n932), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(KEYINPUT122), .B(G2072), .ZN(n933) );
  XNOR2_X1 U1037 ( .A(G33), .B(n933), .ZN(n934) );
  NOR2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n940) );
  XOR2_X1 U1040 ( .A(n938), .B(G27), .Z(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(KEYINPUT53), .B(n941), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1044 ( .A(G2084), .B(G34), .Z(n944) );
  XNOR2_X1 U1045 ( .A(KEYINPUT54), .B(n944), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(G29), .A2(KEYINPUT55), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n949), .A2(n947), .ZN(n948) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n948), .ZN(n978) );
  INV_X1 U1050 ( .A(KEYINPUT55), .ZN(n1000) );
  OR2_X1 U1051 ( .A1(n1000), .A2(n949), .ZN(n976) );
  XNOR2_X1 U1052 ( .A(G5), .B(n950), .ZN(n964) );
  XNOR2_X1 U1053 ( .A(KEYINPUT59), .B(G1348), .ZN(n951) );
  XNOR2_X1 U1054 ( .A(n951), .B(G4), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n1011), .B(G19), .ZN(n954) );
  XNOR2_X1 U1056 ( .A(n952), .B(G20), .ZN(n953) );
  NAND2_X1 U1057 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1058 ( .A(G6), .B(G1981), .ZN(n955) );
  NOR2_X1 U1059 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1060 ( .A1(n958), .A2(n957), .ZN(n960) );
  XOR2_X1 U1061 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n959) );
  XNOR2_X1 U1062 ( .A(n960), .B(n959), .ZN(n962) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G21), .ZN(n961) );
  NOR2_X1 U1064 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1065 ( .A1(n964), .A2(n963), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(G1971), .B(G22), .ZN(n966) );
  XNOR2_X1 U1067 ( .A(G23), .B(G1976), .ZN(n965) );
  NOR2_X1 U1068 ( .A1(n966), .A2(n965), .ZN(n968) );
  XOR2_X1 U1069 ( .A(G1986), .B(G24), .Z(n967) );
  NAND2_X1 U1070 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1071 ( .A(KEYINPUT58), .B(n969), .ZN(n970) );
  NOR2_X1 U1072 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1073 ( .A(KEYINPUT61), .B(n972), .ZN(n974) );
  INV_X1 U1074 ( .A(G16), .ZN(n973) );
  NAND2_X1 U1075 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1076 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n1004) );
  XOR2_X1 U1078 ( .A(G2072), .B(n979), .Z(n981) );
  XOR2_X1 U1079 ( .A(G164), .B(G2078), .Z(n980) );
  NOR2_X1 U1080 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1081 ( .A(KEYINPUT50), .B(n982), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(G2084), .B(G160), .ZN(n983) );
  XNOR2_X1 U1083 ( .A(KEYINPUT121), .B(n983), .ZN(n984) );
  NOR2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1085 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1086 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n998) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1089 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1090 ( .A(KEYINPUT51), .B(n994), .Z(n995) );
  NAND2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(KEYINPUT52), .B(n999), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(G29), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1034) );
  XOR2_X1 U1097 ( .A(G16), .B(KEYINPUT56), .Z(n1032) );
  XNOR2_X1 U1098 ( .A(G171), .B(G1961), .ZN(n1006) );
  NAND2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1029) );
  XOR2_X1 U1100 ( .A(G168), .B(G1966), .Z(n1007) );
  NOR2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1102 ( .A(KEYINPUT57), .B(n1009), .Z(n1027) );
  XNOR2_X1 U1103 ( .A(n1011), .B(n1010), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(G1348), .B(n1012), .Z(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1025) );
  XNOR2_X1 U1106 ( .A(G166), .B(G1971), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1109 ( .A(KEYINPUT124), .B(n1019), .Z(n1022) );
  XOR2_X1 U1110 ( .A(n1020), .B(G1956), .Z(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1112 ( .A(n1023), .B(KEYINPUT125), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(KEYINPUT126), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1119 ( .A(n1035), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

