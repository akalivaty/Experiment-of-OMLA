

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U557 ( .A1(n766), .A2(n765), .ZN(n767) );
  AND2_X1 U558 ( .A1(n757), .A2(n756), .ZN(n766) );
  INV_X2 U559 ( .A(n729), .ZN(n717) );
  NOR2_X1 U560 ( .A1(n947), .A2(n701), .ZN(n696) );
  AND2_X1 U561 ( .A1(n749), .A2(n740), .ZN(n739) );
  NOR2_X1 U562 ( .A1(G651), .A2(n642), .ZN(n647) );
  XOR2_X1 U563 ( .A(KEYINPUT30), .B(n733), .Z(n523) );
  INV_X1 U564 ( .A(KEYINPUT31), .ZN(n737) );
  XNOR2_X1 U565 ( .A(n738), .B(n737), .ZN(n748) );
  AND2_X1 U566 ( .A1(n749), .A2(n748), .ZN(n754) );
  INV_X1 U567 ( .A(G651), .ZN(n537) );
  NOR2_X2 U568 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  AND2_X1 U569 ( .A1(n531), .A2(G2104), .ZN(n891) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n639) );
  AND2_X1 U571 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U572 ( .A1(n530), .A2(n529), .ZN(n689) );
  INV_X1 U573 ( .A(G2105), .ZN(n531) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n531), .ZN(n895) );
  NAND2_X1 U575 ( .A1(G125), .A2(n895), .ZN(n530) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n524), .Z(n890) );
  NAND2_X1 U577 ( .A1(G137), .A2(n890), .ZN(n527) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n898) );
  NAND2_X1 U579 ( .A1(n898), .A2(G113), .ZN(n525) );
  XNOR2_X1 U580 ( .A(n525), .B(KEYINPUT64), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U582 ( .A(n528), .B(KEYINPUT65), .ZN(n529) );
  NAND2_X1 U583 ( .A1(G101), .A2(n891), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT23), .B(n532), .Z(n687) );
  AND2_X1 U585 ( .A1(n689), .A2(n687), .ZN(G160) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n642) );
  NAND2_X1 U587 ( .A1(G47), .A2(n647), .ZN(n536) );
  NOR2_X1 U588 ( .A1(G543), .A2(n537), .ZN(n533) );
  XOR2_X1 U589 ( .A(KEYINPUT66), .B(n533), .Z(n534) );
  XNOR2_X2 U590 ( .A(KEYINPUT1), .B(n534), .ZN(n646) );
  NAND2_X1 U591 ( .A1(G60), .A2(n646), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n541) );
  NAND2_X1 U593 ( .A1(G85), .A2(n639), .ZN(n539) );
  NOR2_X1 U594 ( .A1(n642), .A2(n537), .ZN(n635) );
  NAND2_X1 U595 ( .A1(G72), .A2(n635), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U597 ( .A1(n541), .A2(n540), .ZN(G290) );
  NAND2_X1 U598 ( .A1(G99), .A2(n891), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G111), .A2(n898), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G135), .A2(n890), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n895), .A2(G123), .ZN(n544) );
  XOR2_X1 U603 ( .A(KEYINPUT18), .B(n544), .Z(n545) );
  NOR2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U606 ( .A(n549), .B(KEYINPUT82), .ZN(n992) );
  XNOR2_X1 U607 ( .A(n992), .B(G2096), .ZN(n550) );
  OR2_X1 U608 ( .A1(G2100), .A2(n550), .ZN(G156) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  INV_X1 U610 ( .A(G69), .ZN(G235) );
  INV_X1 U611 ( .A(G108), .ZN(G238) );
  INV_X1 U612 ( .A(G120), .ZN(G236) );
  NAND2_X1 U613 ( .A1(G52), .A2(n647), .ZN(n551) );
  XNOR2_X1 U614 ( .A(n551), .B(KEYINPUT67), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G90), .A2(n639), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G77), .A2(n635), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(KEYINPUT9), .ZN(n556) );
  NAND2_X1 U619 ( .A1(G64), .A2(n646), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U621 ( .A1(n558), .A2(n557), .ZN(G171) );
  NAND2_X1 U622 ( .A1(n639), .A2(G89), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G76), .A2(n635), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT5), .ZN(n569) );
  XNOR2_X1 U627 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n567) );
  NAND2_X1 U628 ( .A1(G63), .A2(n646), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT76), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G51), .A2(n647), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT79), .B(KEYINPUT7), .Z(n570) );
  XNOR2_X1 U635 ( .A(KEYINPUT78), .B(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(G168) );
  XOR2_X1 U637 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U638 ( .A1(G94), .A2(G452), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT68), .B(n573), .Z(G173) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT10), .ZN(n575) );
  XNOR2_X1 U642 ( .A(KEYINPUT70), .B(n575), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n834) );
  NAND2_X1 U644 ( .A1(n834), .A2(G567), .ZN(n576) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  INV_X1 U646 ( .A(G860), .ZN(n617) );
  NAND2_X1 U647 ( .A1(n639), .A2(G81), .ZN(n577) );
  XNOR2_X1 U648 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G68), .A2(n635), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n581) );
  XOR2_X1 U651 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n580) );
  XNOR2_X1 U652 ( .A(n581), .B(n580), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n646), .A2(G56), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT14), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT71), .ZN(n584) );
  NOR2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n647), .A2(G43), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n927) );
  NOR2_X1 U659 ( .A1(n617), .A2(n927), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n588), .B(KEYINPUT73), .ZN(G153) );
  INV_X1 U661 ( .A(G171), .ZN(G301) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G92), .A2(n639), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G66), .A2(n646), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U666 ( .A(KEYINPUT74), .B(n591), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G79), .A2(n635), .ZN(n593) );
  NAND2_X1 U668 ( .A1(G54), .A2(n647), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U671 ( .A(KEYINPUT15), .B(n596), .Z(n597) );
  XNOR2_X1 U672 ( .A(KEYINPUT75), .B(n597), .ZN(n947) );
  INV_X1 U673 ( .A(G868), .ZN(n657) );
  NAND2_X1 U674 ( .A1(n947), .A2(n657), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U676 ( .A1(G53), .A2(n647), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G65), .A2(n646), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G91), .A2(n639), .ZN(n603) );
  NAND2_X1 U680 ( .A1(G78), .A2(n635), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n930) );
  XNOR2_X1 U683 ( .A(n930), .B(KEYINPUT69), .ZN(G299) );
  XOR2_X1 U684 ( .A(G868), .B(KEYINPUT80), .Z(n606) );
  NOR2_X1 U685 ( .A1(G286), .A2(n606), .ZN(n607) );
  XOR2_X1 U686 ( .A(KEYINPUT81), .B(n607), .Z(n609) );
  NOR2_X1 U687 ( .A1(G868), .A2(G299), .ZN(n608) );
  NOR2_X1 U688 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n617), .A2(G559), .ZN(n610) );
  INV_X1 U690 ( .A(n947), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n610), .A2(n615), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(G868), .A2(n927), .ZN(n614) );
  NAND2_X1 U694 ( .A1(G868), .A2(n615), .ZN(n612) );
  NOR2_X1 U695 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U696 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U697 ( .A1(G559), .A2(n615), .ZN(n616) );
  XOR2_X1 U698 ( .A(n927), .B(n616), .Z(n655) );
  NAND2_X1 U699 ( .A1(n617), .A2(n655), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G93), .A2(n639), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G55), .A2(n647), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G67), .A2(n646), .ZN(n620) );
  XNOR2_X1 U704 ( .A(KEYINPUT83), .B(n620), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n635), .A2(G80), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n658) );
  XNOR2_X1 U708 ( .A(n625), .B(n658), .ZN(G145) );
  NAND2_X1 U709 ( .A1(G50), .A2(n647), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G62), .A2(n646), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U712 ( .A(KEYINPUT84), .B(n628), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G88), .A2(n639), .ZN(n630) );
  NAND2_X1 U714 ( .A1(G75), .A2(n635), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U716 ( .A1(n632), .A2(n631), .ZN(G166) );
  NAND2_X1 U717 ( .A1(G48), .A2(n647), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G61), .A2(n646), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n639), .A2(G86), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U725 ( .A1(G87), .A2(n642), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n647), .A2(G49), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(G288) );
  XNOR2_X1 U731 ( .A(G166), .B(G299), .ZN(n654) );
  XNOR2_X1 U732 ( .A(G305), .B(G290), .ZN(n652) );
  XOR2_X1 U733 ( .A(KEYINPUT19), .B(G288), .Z(n650) );
  XNOR2_X1 U734 ( .A(n658), .B(n650), .ZN(n651) );
  XNOR2_X1 U735 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U736 ( .A(n654), .B(n653), .ZN(n861) );
  XNOR2_X1 U737 ( .A(n655), .B(n861), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(G295) );
  XOR2_X1 U741 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n664) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n661) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U744 ( .A1(n662), .A2(G2090), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G2072), .A2(n665), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U748 ( .A1(G132), .A2(G82), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n666), .B(KEYINPUT86), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n667), .B(KEYINPUT22), .ZN(n668) );
  NOR2_X1 U751 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U752 ( .A1(G96), .A2(n669), .ZN(n838) );
  NAND2_X1 U753 ( .A1(G2106), .A2(n838), .ZN(n670) );
  XNOR2_X1 U754 ( .A(KEYINPUT87), .B(n670), .ZN(n676) );
  NOR2_X1 U755 ( .A1(G236), .A2(G238), .ZN(n672) );
  NOR2_X1 U756 ( .A1(G235), .A2(G237), .ZN(n671) );
  NAND2_X1 U757 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U758 ( .A(KEYINPUT88), .B(n673), .ZN(n839) );
  NAND2_X1 U759 ( .A1(n839), .A2(G567), .ZN(n674) );
  XNOR2_X1 U760 ( .A(KEYINPUT89), .B(n674), .ZN(n675) );
  NOR2_X1 U761 ( .A1(n676), .A2(n675), .ZN(G319) );
  INV_X1 U762 ( .A(G319), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U764 ( .A1(n678), .A2(n677), .ZN(n837) );
  NAND2_X1 U765 ( .A1(n837), .A2(G36), .ZN(n679) );
  XNOR2_X1 U766 ( .A(KEYINPUT90), .B(n679), .ZN(G176) );
  NAND2_X1 U767 ( .A1(n890), .A2(G138), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G102), .A2(n891), .ZN(n680) );
  XOR2_X1 U769 ( .A(KEYINPUT91), .B(n680), .Z(n681) );
  NAND2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U771 ( .A1(G114), .A2(n898), .ZN(n684) );
  NAND2_X1 U772 ( .A1(G126), .A2(n895), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U774 ( .A1(n686), .A2(n685), .ZN(G164) );
  XOR2_X1 U775 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  XOR2_X1 U776 ( .A(G1981), .B(G305), .Z(n942) );
  AND2_X1 U777 ( .A1(G40), .A2(n687), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n818) );
  INV_X1 U779 ( .A(n818), .ZN(n690) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n819) );
  NAND2_X1 U781 ( .A1(n690), .A2(n819), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n717), .A2(G1996), .ZN(n691) );
  XNOR2_X1 U783 ( .A(KEYINPUT26), .B(n691), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n729), .A2(G1341), .ZN(n692) );
  XNOR2_X1 U785 ( .A(n692), .B(KEYINPUT101), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n927), .A2(n693), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n701) );
  XOR2_X1 U788 ( .A(n696), .B(KEYINPUT102), .Z(n700) );
  NOR2_X1 U789 ( .A1(G2067), .A2(n729), .ZN(n698) );
  NOR2_X1 U790 ( .A1(n717), .A2(G1348), .ZN(n697) );
  NOR2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n947), .A2(n701), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n708) );
  NAND2_X1 U795 ( .A1(n717), .A2(G2072), .ZN(n704) );
  XNOR2_X1 U796 ( .A(n704), .B(KEYINPUT27), .ZN(n706) );
  INV_X1 U797 ( .A(G1956), .ZN(n1015) );
  NOR2_X1 U798 ( .A1(n1015), .A2(n717), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n930), .A2(n710), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U802 ( .A(KEYINPUT103), .B(n709), .ZN(n714) );
  NOR2_X1 U803 ( .A1(n930), .A2(n710), .ZN(n711) );
  XNOR2_X1 U804 ( .A(KEYINPUT100), .B(n711), .ZN(n712) );
  XNOR2_X1 U805 ( .A(KEYINPUT28), .B(n712), .ZN(n713) );
  NOR2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U807 ( .A(n715), .B(KEYINPUT29), .ZN(n721) );
  XOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  NOR2_X1 U809 ( .A1(n961), .A2(n729), .ZN(n716) );
  XNOR2_X1 U810 ( .A(n716), .B(KEYINPUT99), .ZN(n719) );
  OR2_X1 U811 ( .A1(G1961), .A2(n717), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n734) );
  NAND2_X1 U813 ( .A1(G171), .A2(n734), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n749) );
  INV_X1 U815 ( .A(G8), .ZN(n728) );
  NAND2_X1 U816 ( .A1(n729), .A2(G8), .ZN(n722) );
  XOR2_X2 U817 ( .A(KEYINPUT97), .B(n722), .Z(n779) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n779), .ZN(n723) );
  XNOR2_X1 U819 ( .A(n723), .B(KEYINPUT106), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n729), .A2(G2090), .ZN(n724) );
  NOR2_X1 U821 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U822 ( .A1(n726), .A2(G303), .ZN(n727) );
  OR2_X1 U823 ( .A1(n728), .A2(n727), .ZN(n740) );
  NOR2_X1 U824 ( .A1(G1966), .A2(n779), .ZN(n751) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n729), .ZN(n750) );
  NOR2_X1 U826 ( .A1(n751), .A2(n750), .ZN(n730) );
  XNOR2_X1 U827 ( .A(n730), .B(KEYINPUT104), .ZN(n731) );
  NAND2_X1 U828 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U829 ( .A(n732), .B(KEYINPUT105), .ZN(n733) );
  NOR2_X1 U830 ( .A1(n523), .A2(G168), .ZN(n736) );
  NOR2_X1 U831 ( .A1(G171), .A2(n734), .ZN(n735) );
  NOR2_X1 U832 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U833 ( .A1(n739), .A2(n748), .ZN(n744) );
  INV_X1 U834 ( .A(n740), .ZN(n742) );
  AND2_X1 U835 ( .A1(G286), .A2(G8), .ZN(n741) );
  OR2_X1 U836 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U837 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U838 ( .A(n745), .B(KEYINPUT32), .ZN(n773) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n931) );
  INV_X1 U840 ( .A(n931), .ZN(n746) );
  OR2_X1 U841 ( .A1(n779), .A2(n746), .ZN(n760) );
  INV_X1 U842 ( .A(n760), .ZN(n747) );
  AND2_X1 U843 ( .A1(n773), .A2(n747), .ZN(n757) );
  AND2_X1 U844 ( .A1(G8), .A2(n750), .ZN(n752) );
  OR2_X1 U845 ( .A1(n752), .A2(n751), .ZN(n753) );
  OR2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n774) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n759), .A2(KEYINPUT33), .ZN(n755) );
  OR2_X1 U849 ( .A1(n779), .A2(n755), .ZN(n764) );
  AND2_X1 U850 ( .A1(n774), .A2(n764), .ZN(n756) );
  NOR2_X1 U851 ( .A1(G303), .A2(G1971), .ZN(n758) );
  NOR2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n936) );
  OR2_X1 U853 ( .A1(n760), .A2(n936), .ZN(n762) );
  INV_X1 U854 ( .A(KEYINPUT33), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n763) );
  AND2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n942), .A2(n767), .ZN(n769) );
  INV_X1 U858 ( .A(KEYINPUT107), .ZN(n768) );
  XNOR2_X1 U859 ( .A(n769), .B(n768), .ZN(n824) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n770) );
  XOR2_X1 U861 ( .A(n770), .B(KEYINPUT24), .Z(n771) );
  NOR2_X1 U862 ( .A1(n779), .A2(n771), .ZN(n772) );
  XNOR2_X1 U863 ( .A(n772), .B(KEYINPUT98), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n777) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n775) );
  NAND2_X1 U866 ( .A1(G8), .A2(n775), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n778) );
  AND2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n822) );
  NAND2_X1 U870 ( .A1(G117), .A2(n898), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G141), .A2(n890), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n891), .A2(G105), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n895), .A2(G129), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n885) );
  NOR2_X1 U878 ( .A1(n885), .A2(G1996), .ZN(n789) );
  XNOR2_X1 U879 ( .A(n789), .B(KEYINPUT108), .ZN(n984) );
  NAND2_X1 U880 ( .A1(G1996), .A2(n885), .ZN(n790) );
  XNOR2_X1 U881 ( .A(n790), .B(KEYINPUT96), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G131), .A2(n890), .ZN(n792) );
  NAND2_X1 U883 ( .A1(G95), .A2(n891), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G107), .A2(n898), .ZN(n794) );
  NAND2_X1 U886 ( .A1(G119), .A2(n895), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n873) );
  NAND2_X1 U889 ( .A1(G1991), .A2(n873), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n989) );
  NOR2_X1 U891 ( .A1(G1991), .A2(n873), .ZN(n990) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n990), .A2(n799), .ZN(n800) );
  NOR2_X1 U894 ( .A1(n989), .A2(n800), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n984), .A2(n801), .ZN(n802) );
  XNOR2_X1 U896 ( .A(n802), .B(KEYINPUT39), .ZN(n814) );
  XNOR2_X1 U897 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NAND2_X1 U898 ( .A1(n891), .A2(G104), .ZN(n803) );
  XNOR2_X1 U899 ( .A(n803), .B(KEYINPUT94), .ZN(n805) );
  NAND2_X1 U900 ( .A1(G140), .A2(n890), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n806), .ZN(n811) );
  NAND2_X1 U903 ( .A1(G116), .A2(n898), .ZN(n808) );
  NAND2_X1 U904 ( .A1(G128), .A2(n895), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U906 ( .A(KEYINPUT35), .B(n809), .Z(n810) );
  NOR2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U908 ( .A(n812), .B(KEYINPUT95), .ZN(n813) );
  XOR2_X1 U909 ( .A(n813), .B(KEYINPUT36), .Z(n904) );
  OR2_X1 U910 ( .A1(n815), .A2(n904), .ZN(n988) );
  NAND2_X1 U911 ( .A1(n814), .A2(n988), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n815), .A2(n904), .ZN(n987) );
  NAND2_X1 U913 ( .A1(n816), .A2(n987), .ZN(n817) );
  XOR2_X1 U914 ( .A(KEYINPUT109), .B(n817), .Z(n821) );
  NOR2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U916 ( .A(KEYINPUT93), .B(n820), .Z(n827) );
  NAND2_X1 U917 ( .A1(n821), .A2(n827), .ZN(n825) );
  AND2_X1 U918 ( .A1(n822), .A2(n825), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n832) );
  INV_X1 U920 ( .A(n825), .ZN(n830) );
  XNOR2_X1 U921 ( .A(G1986), .B(G290), .ZN(n938) );
  NOR2_X1 U922 ( .A1(n989), .A2(n938), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n826), .A2(n988), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n828), .A2(n827), .ZN(n829) );
  OR2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U933 ( .A(G132), .ZN(G219) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XOR2_X1 U937 ( .A(KEYINPUT114), .B(G1991), .Z(n841) );
  XNOR2_X1 U938 ( .A(G1956), .B(G1996), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U940 ( .A(n842), .B(KEYINPUT41), .Z(n844) );
  XNOR2_X1 U941 ( .A(G1971), .B(G1986), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(G1976), .B(G1981), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1961), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U947 ( .A(KEYINPUT115), .B(G2474), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(G229) );
  XOR2_X1 U949 ( .A(KEYINPUT113), .B(G2067), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2078), .B(G2072), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n853), .B(G2100), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2084), .B(G2090), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U955 ( .A(G2096), .B(G2678), .Z(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n859), .B(n858), .Z(G227) );
  XNOR2_X1 U959 ( .A(G171), .B(n927), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(G286), .ZN(n863) );
  XOR2_X1 U961 ( .A(n947), .B(n861), .Z(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  NOR2_X1 U963 ( .A1(G37), .A2(n864), .ZN(G397) );
  NAND2_X1 U964 ( .A1(n895), .A2(G124), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n890), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U968 ( .A(KEYINPUT116), .B(n868), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G112), .A2(n898), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G100), .A2(n891), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U972 ( .A1(n872), .A2(n871), .ZN(G162) );
  XNOR2_X1 U973 ( .A(KEYINPUT119), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n873), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n887) );
  NAND2_X1 U976 ( .A1(G139), .A2(n890), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G103), .A2(n891), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G115), .A2(n898), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G127), .A2(n895), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U982 ( .A(KEYINPUT118), .B(n880), .Z(n881) );
  XNOR2_X1 U983 ( .A(KEYINPUT47), .B(n881), .ZN(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n977) );
  XOR2_X1 U985 ( .A(n977), .B(n992), .Z(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U987 ( .A(n887), .B(n886), .Z(n889) );
  XNOR2_X1 U988 ( .A(G164), .B(G160), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n903) );
  NAND2_X1 U990 ( .A1(G142), .A2(n890), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G106), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n894), .B(KEYINPUT45), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n901) );
  NAND2_X1 U996 ( .A1(G118), .A2(n898), .ZN(n899) );
  XNOR2_X1 U997 ( .A(KEYINPUT117), .B(n899), .ZN(n900) );
  NOR2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U999 ( .A(n903), .B(n902), .Z(n906) );
  XOR2_X1 U1000 ( .A(n904), .B(G162), .Z(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1002 ( .A1(n907), .A2(G37), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n908), .B(KEYINPUT120), .ZN(G395) );
  XOR2_X1 U1004 ( .A(KEYINPUT112), .B(G2438), .Z(n910) );
  XNOR2_X1 U1005 ( .A(G2451), .B(KEYINPUT111), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1007 ( .A(G2443), .B(KEYINPUT110), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G2430), .B(G2454), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1011 ( .A(G2435), .B(G2427), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n919) );
  XOR2_X1 U1013 ( .A(G1348), .B(G1341), .Z(n917) );
  XNOR2_X1 U1014 ( .A(G2446), .B(n917), .ZN(n918) );
  XOR2_X1 U1015 ( .A(n919), .B(n918), .Z(n920) );
  NAND2_X1 U1016 ( .A1(G14), .A2(n920), .ZN(n926) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n926), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(G397), .A2(G395), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G96), .ZN(G221) );
  INV_X1 U1025 ( .A(n926), .ZN(G401) );
  XNOR2_X1 U1026 ( .A(KEYINPUT56), .B(G16), .ZN(n951) );
  XNOR2_X1 U1027 ( .A(G301), .B(G1961), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(n927), .B(G1341), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n941) );
  XNOR2_X1 U1030 ( .A(n930), .B(G1956), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n934) );
  AND2_X1 U1032 ( .A1(G303), .A2(G1971), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(n939), .B(KEYINPUT124), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G1966), .B(G168), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1040 ( .A(KEYINPUT57), .B(n944), .Z(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1042 ( .A(G1348), .B(n947), .Z(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(KEYINPUT125), .B(n952), .ZN(n976) );
  XNOR2_X1 U1046 ( .A(G2072), .B(G33), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1049 ( .A(G2067), .B(G26), .Z(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G25), .B(G1991), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G27), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT53), .B(n964), .Z(n967) );
  XOR2_X1 U1058 ( .A(KEYINPUT54), .B(G34), .Z(n965) );
  XNOR2_X1 U1059 ( .A(G2084), .B(n965), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G35), .B(G2090), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(n970), .B(KEYINPUT55), .ZN(n972) );
  INV_X1 U1064 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n973), .ZN(n974) );
  XOR2_X1 U1067 ( .A(KEYINPUT123), .B(n974), .Z(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n1004) );
  XOR2_X1 U1069 ( .A(G2072), .B(n977), .Z(n979) );
  XOR2_X1 U1070 ( .A(G164), .B(G2078), .Z(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(KEYINPUT50), .B(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G160), .B(G2084), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n998) );
  XOR2_X1 U1075 ( .A(G2090), .B(G162), .Z(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT121), .B(n985), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n986), .B(KEYINPUT51), .ZN(n996) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n994) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(KEYINPUT52), .B(n999), .ZN(n1001) );
  INV_X1 U1086 ( .A(KEYINPUT55), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(G29), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1030) );
  XOR2_X1 U1090 ( .A(G1986), .B(G24), .Z(n1008) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G22), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1010), .B(n1009), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G5), .B(G1961), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1025) );
  XNOR2_X1 U1101 ( .A(G20), .B(n1015), .ZN(n1019) );
  XNOR2_X1 U1102 ( .A(G1341), .B(G19), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G6), .B(G1981), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XOR2_X1 U1106 ( .A(KEYINPUT59), .B(G1348), .Z(n1020) );
  XNOR2_X1 U1107 ( .A(G4), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(KEYINPUT60), .B(n1023), .Z(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1026), .Z(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT126), .B(G16), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(n1031), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

