

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U548 ( .A(n737), .B(KEYINPUT32), .ZN(n755) );
  AND2_X2 U549 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X2 U550 ( .A(KEYINPUT1), .B(n536), .Z(n643) );
  NOR2_X2 U551 ( .A1(n684), .A2(n789), .ZN(n693) );
  INV_X1 U552 ( .A(KEYINPUT105), .ZN(n749) );
  NOR2_X1 U553 ( .A1(n748), .A2(n747), .ZN(n750) );
  AND2_X1 U554 ( .A1(n766), .A2(n512), .ZN(n767) );
  AND2_X1 U555 ( .A1(n765), .A2(n515), .ZN(n512) );
  AND2_X1 U556 ( .A1(n804), .A2(n818), .ZN(n513) );
  OR2_X1 U557 ( .A1(n805), .A2(n513), .ZN(n514) );
  OR2_X1 U558 ( .A1(n764), .A2(n763), .ZN(n515) );
  NOR2_X1 U559 ( .A1(n761), .A2(n764), .ZN(n516) );
  INV_X1 U560 ( .A(n693), .ZN(n728) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X1 U562 ( .A(KEYINPUT15), .B(n601), .Z(n964) );
  NOR2_X1 U563 ( .A1(G651), .A2(n628), .ZN(n646) );
  BUF_X1 U564 ( .A(n680), .Z(G160) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n517), .Z(n883) );
  NAND2_X1 U566 ( .A1(n883), .A2(G137), .ZN(n519) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U568 ( .A1(n879), .A2(G113), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n519), .A2(n518), .ZN(n526) );
  INV_X1 U570 ( .A(G2104), .ZN(n520) );
  NOR2_X1 U571 ( .A1(n520), .A2(G2105), .ZN(n547) );
  NAND2_X1 U572 ( .A1(n547), .A2(G101), .ZN(n521) );
  XOR2_X1 U573 ( .A(n521), .B(KEYINPUT23), .Z(n523) );
  AND2_X1 U574 ( .A1(n520), .A2(G2105), .ZN(n878) );
  NAND2_X1 U575 ( .A1(n878), .A2(G125), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(n524), .Z(n525) );
  NOR2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n680) );
  XOR2_X1 U579 ( .A(G2443), .B(G2446), .Z(n528) );
  XNOR2_X1 U580 ( .A(G2427), .B(G2451), .ZN(n527) );
  XNOR2_X1 U581 ( .A(n528), .B(n527), .ZN(n534) );
  XOR2_X1 U582 ( .A(G2430), .B(G2454), .Z(n530) );
  XNOR2_X1 U583 ( .A(G1348), .B(G1341), .ZN(n529) );
  XNOR2_X1 U584 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U585 ( .A(G2435), .B(G2438), .Z(n531) );
  XNOR2_X1 U586 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U587 ( .A(n534), .B(n533), .Z(n535) );
  AND2_X1 U588 ( .A1(G14), .A2(n535), .ZN(G401) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  NAND2_X1 U590 ( .A1(n646), .A2(G52), .ZN(n538) );
  XNOR2_X1 U591 ( .A(KEYINPUT67), .B(G651), .ZN(n539) );
  NOR2_X1 U592 ( .A1(G543), .A2(n539), .ZN(n536) );
  NAND2_X1 U593 ( .A1(G64), .A2(n643), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n545) );
  NOR2_X1 U595 ( .A1(n628), .A2(n539), .ZN(n647) );
  NAND2_X1 U596 ( .A1(G77), .A2(n647), .ZN(n540) );
  XNOR2_X1 U597 ( .A(n540), .B(KEYINPUT68), .ZN(n542) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U599 ( .A1(G90), .A2(n642), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n543), .Z(n544) );
  NOR2_X1 U602 ( .A1(n545), .A2(n544), .ZN(G171) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U604 ( .A1(n879), .A2(G111), .ZN(n546) );
  XOR2_X1 U605 ( .A(KEYINPUT77), .B(n546), .Z(n549) );
  BUF_X1 U606 ( .A(n547), .Z(n886) );
  NAND2_X1 U607 ( .A1(n886), .A2(G99), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U609 ( .A(KEYINPUT78), .B(n550), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n878), .A2(G123), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT18), .B(n551), .Z(n552) );
  NOR2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n883), .A2(G135), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n924) );
  XNOR2_X1 U615 ( .A(G2096), .B(n924), .ZN(n556) );
  OR2_X1 U616 ( .A1(G2100), .A2(n556), .ZN(G156) );
  NAND2_X1 U617 ( .A1(n646), .A2(G53), .ZN(n558) );
  NAND2_X1 U618 ( .A1(G65), .A2(n643), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G91), .A2(n642), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G78), .A2(n647), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n970) );
  INV_X1 U624 ( .A(n970), .ZN(G299) );
  INV_X1 U625 ( .A(G82), .ZN(G220) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G120), .ZN(G236) );
  NAND2_X1 U628 ( .A1(n886), .A2(G102), .ZN(n565) );
  NAND2_X1 U629 ( .A1(G114), .A2(n879), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT87), .B(n563), .Z(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G126), .A2(n878), .ZN(n567) );
  NAND2_X1 U633 ( .A1(G138), .A2(n883), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(G164) );
  NAND2_X1 U636 ( .A1(G89), .A2(n642), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT74), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT4), .B(n571), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G76), .A2(n647), .ZN(n572) );
  XOR2_X1 U640 ( .A(KEYINPUT75), .B(n572), .Z(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT5), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n646), .A2(G51), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G63), .A2(n643), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U646 ( .A(KEYINPUT6), .B(n578), .Z(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U649 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U650 ( .A1(G7), .A2(G661), .ZN(n582) );
  XOR2_X1 U651 ( .A(n582), .B(KEYINPUT10), .Z(n823) );
  NAND2_X1 U652 ( .A1(n823), .A2(G567), .ZN(n583) );
  XOR2_X1 U653 ( .A(KEYINPUT11), .B(n583), .Z(G234) );
  XOR2_X1 U654 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n585) );
  NAND2_X1 U655 ( .A1(G56), .A2(n643), .ZN(n584) );
  XNOR2_X1 U656 ( .A(n585), .B(n584), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n642), .A2(G81), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G68), .A2(n647), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U661 ( .A(KEYINPUT13), .B(n589), .Z(n590) );
  NOR2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n646), .A2(G43), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n960) );
  XNOR2_X1 U665 ( .A(G860), .B(KEYINPUT71), .ZN(n607) );
  OR2_X1 U666 ( .A1(n960), .A2(n607), .ZN(G153) );
  NAND2_X1 U667 ( .A1(G868), .A2(G171), .ZN(n603) );
  NAND2_X1 U668 ( .A1(G66), .A2(n643), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n642), .A2(G92), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n596), .B(KEYINPUT72), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n646), .A2(G54), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G79), .A2(n647), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  INV_X1 U676 ( .A(G868), .ZN(n662) );
  NAND2_X1 U677 ( .A1(n964), .A2(n662), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT73), .ZN(G284) );
  NOR2_X1 U680 ( .A1(G286), .A2(n662), .ZN(n606) );
  NOR2_X1 U681 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U682 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U683 ( .A1(G559), .A2(n607), .ZN(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT76), .B(n608), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n609), .A2(n964), .ZN(n610) );
  XNOR2_X1 U686 ( .A(KEYINPUT16), .B(n610), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n960), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G868), .A2(n964), .ZN(n611) );
  NOR2_X1 U689 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U690 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U691 ( .A1(n646), .A2(G50), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G62), .A2(n643), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U694 ( .A(KEYINPUT82), .B(n616), .ZN(n620) );
  NAND2_X1 U695 ( .A1(G88), .A2(n642), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G75), .A2(n647), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U698 ( .A1(n620), .A2(n619), .ZN(G166) );
  INV_X1 U699 ( .A(G166), .ZN(G303) );
  NAND2_X1 U700 ( .A1(G60), .A2(n643), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G72), .A2(n647), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n642), .A2(G85), .ZN(n623) );
  XOR2_X1 U704 ( .A(KEYINPUT66), .B(n623), .Z(n624) );
  NOR2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n646), .A2(G47), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(G290) );
  NAND2_X1 U708 ( .A1(G87), .A2(n628), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U711 ( .A1(n643), .A2(n631), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n646), .A2(G49), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U714 ( .A1(n647), .A2(G73), .ZN(n634) );
  XNOR2_X1 U715 ( .A(n634), .B(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(G86), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G61), .A2(n643), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G48), .A2(n646), .ZN(n637) );
  XNOR2_X1 U720 ( .A(KEYINPUT81), .B(n637), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U723 ( .A1(n642), .A2(G93), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G67), .A2(n643), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n646), .A2(G55), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G80), .A2(n647), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U730 ( .A(KEYINPUT80), .B(n652), .Z(n829) );
  XOR2_X1 U731 ( .A(G303), .B(n829), .Z(n658) );
  XNOR2_X1 U732 ( .A(KEYINPUT19), .B(G290), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n653), .B(G288), .ZN(n654) );
  XNOR2_X1 U734 ( .A(KEYINPUT83), .B(n654), .ZN(n656) );
  XOR2_X1 U735 ( .A(G305), .B(G299), .Z(n655) );
  XNOR2_X1 U736 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n658), .B(n657), .ZN(n897) );
  XNOR2_X1 U738 ( .A(n960), .B(KEYINPUT79), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n964), .A2(G559), .ZN(n659) );
  XOR2_X1 U740 ( .A(n660), .B(n659), .Z(n827) );
  XNOR2_X1 U741 ( .A(n897), .B(n827), .ZN(n661) );
  NOR2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n664) );
  NOR2_X1 U743 ( .A1(n829), .A2(G868), .ZN(n663) );
  NOR2_X1 U744 ( .A1(n664), .A2(n663), .ZN(G295) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n666) );
  NAND2_X1 U746 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U752 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U753 ( .A1(G236), .A2(G237), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G69), .A2(n670), .ZN(n671) );
  XNOR2_X1 U755 ( .A(KEYINPUT85), .B(n671), .ZN(n672) );
  NAND2_X1 U756 ( .A1(n672), .A2(G108), .ZN(n830) );
  NAND2_X1 U757 ( .A1(G567), .A2(n830), .ZN(n673) );
  XNOR2_X1 U758 ( .A(n673), .B(KEYINPUT86), .ZN(n678) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U761 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U762 ( .A1(G96), .A2(n676), .ZN(n831) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n831), .ZN(n677) );
  NAND2_X1 U764 ( .A1(n678), .A2(n677), .ZN(n832) );
  NAND2_X1 U765 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U766 ( .A1(n832), .A2(n679), .ZN(n826) );
  NAND2_X1 U767 ( .A1(n826), .A2(G36), .ZN(G176) );
  INV_X1 U768 ( .A(KEYINPUT98), .ZN(n682) );
  AND2_X1 U769 ( .A1(G40), .A2(n680), .ZN(n681) );
  XNOR2_X1 U770 ( .A(n681), .B(KEYINPUT88), .ZN(n790) );
  XNOR2_X1 U771 ( .A(n682), .B(n790), .ZN(n684) );
  NOR2_X1 U772 ( .A1(G1384), .A2(G164), .ZN(n683) );
  XOR2_X1 U773 ( .A(n683), .B(KEYINPUT64), .Z(n789) );
  NAND2_X1 U774 ( .A1(G8), .A2(n728), .ZN(n764) );
  NOR2_X1 U775 ( .A1(G1966), .A2(n764), .ZN(n740) );
  NOR2_X1 U776 ( .A1(G2084), .A2(n728), .ZN(n738) );
  NOR2_X1 U777 ( .A1(n740), .A2(n738), .ZN(n685) );
  NAND2_X1 U778 ( .A1(G8), .A2(n685), .ZN(n686) );
  XNOR2_X1 U779 ( .A(KEYINPUT30), .B(n686), .ZN(n687) );
  NOR2_X1 U780 ( .A1(G168), .A2(n687), .ZN(n691) );
  XNOR2_X1 U781 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NOR2_X1 U782 ( .A1(n728), .A2(n943), .ZN(n689) );
  INV_X1 U783 ( .A(G1961), .ZN(n845) );
  NOR2_X1 U784 ( .A1(n693), .A2(n845), .ZN(n688) );
  NOR2_X1 U785 ( .A1(n689), .A2(n688), .ZN(n720) );
  NOR2_X1 U786 ( .A1(G171), .A2(n720), .ZN(n690) );
  NOR2_X1 U787 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U788 ( .A(KEYINPUT31), .B(n692), .ZN(n724) );
  AND2_X1 U789 ( .A1(n693), .A2(G1996), .ZN(n694) );
  XNOR2_X1 U790 ( .A(n694), .B(KEYINPUT26), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n728), .A2(G1341), .ZN(n696) );
  INV_X1 U792 ( .A(n960), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n700) );
  NOR2_X1 U795 ( .A1(n700), .A2(n964), .ZN(n699) );
  XNOR2_X1 U796 ( .A(n699), .B(KEYINPUT101), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n700), .A2(n964), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n693), .A2(G1348), .ZN(n702) );
  NOR2_X1 U799 ( .A1(G2067), .A2(n728), .ZN(n701) );
  NOR2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n712) );
  NAND2_X1 U803 ( .A1(G1956), .A2(n728), .ZN(n707) );
  XNOR2_X1 U804 ( .A(KEYINPUT99), .B(n707), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n693), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U806 ( .A(KEYINPUT27), .B(n708), .ZN(n709) );
  NOR2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U808 ( .A1(n713), .A2(n970), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U810 ( .A1(n713), .A2(n970), .ZN(n715) );
  XOR2_X1 U811 ( .A(KEYINPUT100), .B(KEYINPUT28), .Z(n714) );
  XNOR2_X1 U812 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U813 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U814 ( .A(KEYINPUT29), .B(KEYINPUT102), .ZN(n718) );
  XNOR2_X1 U815 ( .A(n719), .B(n718), .ZN(n722) );
  AND2_X1 U816 ( .A1(G171), .A2(n720), .ZN(n721) );
  NOR2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n726) );
  INV_X1 U819 ( .A(KEYINPUT103), .ZN(n725) );
  XNOR2_X1 U820 ( .A(n726), .B(n725), .ZN(n739) );
  INV_X1 U821 ( .A(n739), .ZN(n727) );
  NAND2_X1 U822 ( .A1(n727), .A2(G286), .ZN(n736) );
  INV_X1 U823 ( .A(G8), .ZN(n734) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n728), .ZN(n729) );
  XNOR2_X1 U825 ( .A(n729), .B(KEYINPUT104), .ZN(n731) );
  NOR2_X1 U826 ( .A1(n764), .A2(G1971), .ZN(n730) );
  NOR2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U828 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U829 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U830 ( .A1(G8), .A2(n738), .ZN(n742) );
  NOR2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n756) );
  AND2_X1 U833 ( .A1(n756), .A2(n764), .ZN(n743) );
  AND2_X1 U834 ( .A1(n755), .A2(n743), .ZN(n748) );
  INV_X1 U835 ( .A(n764), .ZN(n746) );
  NOR2_X1 U836 ( .A1(G2090), .A2(G303), .ZN(n744) );
  NAND2_X1 U837 ( .A1(G8), .A2(n744), .ZN(n745) );
  NOR2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U839 ( .A(n750), .B(n749), .ZN(n754) );
  NOR2_X1 U840 ( .A1(G1981), .A2(G305), .ZN(n751) );
  XOR2_X1 U841 ( .A(n751), .B(KEYINPUT24), .Z(n752) );
  OR2_X1 U842 ( .A1(n764), .A2(n752), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n769) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n760) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n762) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U847 ( .A1(n762), .A2(n757), .ZN(n978) );
  INV_X1 U848 ( .A(KEYINPUT33), .ZN(n758) );
  AND2_X1 U849 ( .A1(n978), .A2(n758), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n766) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n968) );
  INV_X1 U852 ( .A(n968), .ZN(n761) );
  OR2_X1 U853 ( .A1(KEYINPUT33), .A2(n516), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n762), .A2(KEYINPUT33), .ZN(n763) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n957) );
  AND2_X1 U856 ( .A1(n767), .A2(n957), .ZN(n768) );
  NOR2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n806) );
  NAND2_X1 U858 ( .A1(G119), .A2(n878), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G107), .A2(n879), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U861 ( .A(KEYINPUT92), .B(n772), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G95), .A2(n886), .ZN(n773) );
  XNOR2_X1 U863 ( .A(KEYINPUT93), .B(n773), .ZN(n774) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n883), .A2(G131), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n890) );
  NAND2_X1 U867 ( .A1(G1991), .A2(n890), .ZN(n778) );
  XNOR2_X1 U868 ( .A(n778), .B(KEYINPUT94), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G129), .A2(n878), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G117), .A2(n879), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n886), .A2(G105), .ZN(n781) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n883), .A2(G141), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n864) );
  NAND2_X1 U877 ( .A1(G1996), .A2(n864), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U879 ( .A(KEYINPUT95), .B(n788), .ZN(n921) );
  AND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n818) );
  XOR2_X1 U881 ( .A(KEYINPUT96), .B(n818), .Z(n791) );
  NOR2_X1 U882 ( .A1(n921), .A2(n791), .ZN(n810) );
  XOR2_X1 U883 ( .A(KEYINPUT97), .B(n810), .Z(n805) );
  XOR2_X1 U884 ( .A(G1986), .B(G290), .Z(n969) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  XNOR2_X1 U886 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G128), .A2(n878), .ZN(n793) );
  NAND2_X1 U888 ( .A1(G116), .A2(n879), .ZN(n792) );
  NAND2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U890 ( .A(n794), .B(KEYINPUT35), .ZN(n795) );
  XNOR2_X1 U891 ( .A(n796), .B(n795), .ZN(n802) );
  NAND2_X1 U892 ( .A1(G104), .A2(n886), .ZN(n798) );
  NAND2_X1 U893 ( .A1(G140), .A2(n883), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U895 ( .A(KEYINPUT34), .B(n799), .ZN(n800) );
  XOR2_X1 U896 ( .A(KEYINPUT89), .B(n800), .Z(n801) );
  NOR2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U898 ( .A(KEYINPUT36), .B(n803), .ZN(n891) );
  NOR2_X1 U899 ( .A1(n816), .A2(n891), .ZN(n814) );
  INV_X1 U900 ( .A(n814), .ZN(n908) );
  NAND2_X1 U901 ( .A1(n969), .A2(n908), .ZN(n804) );
  OR2_X1 U902 ( .A1(n806), .A2(n514), .ZN(n821) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n864), .ZN(n916) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n890), .ZN(n926) );
  NOR2_X1 U906 ( .A1(n807), .A2(n926), .ZN(n808) );
  XNOR2_X1 U907 ( .A(n808), .B(KEYINPUT106), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n916), .A2(n811), .ZN(n812) );
  XOR2_X1 U910 ( .A(KEYINPUT39), .B(n812), .Z(n813) );
  NOR2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U912 ( .A(n815), .B(KEYINPUT107), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n816), .A2(n891), .ZN(n909) );
  NAND2_X1 U914 ( .A1(n817), .A2(n909), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(KEYINPUT40), .B(n822), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n823), .ZN(G217) );
  INV_X1 U919 ( .A(n823), .ZN(G223) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U921 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U923 ( .A1(n826), .A2(n825), .ZN(G188) );
  NOR2_X1 U925 ( .A1(G860), .A2(n827), .ZN(n828) );
  XOR2_X1 U926 ( .A(n829), .B(n828), .Z(G145) );
  INV_X1 U927 ( .A(G108), .ZN(G238) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  NOR2_X1 U929 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  XOR2_X1 U931 ( .A(KEYINPUT108), .B(n832), .Z(G319) );
  XOR2_X1 U932 ( .A(KEYINPUT42), .B(G2090), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2084), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n835), .B(G2100), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2072), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U939 ( .A(G2678), .B(KEYINPUT109), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n841), .B(n840), .Z(G227) );
  XOR2_X1 U942 ( .A(KEYINPUT110), .B(G1981), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U945 ( .A(n844), .B(G2474), .Z(n847) );
  XOR2_X1 U946 ( .A(G1971), .B(n845), .Z(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(G1956), .B(G1966), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1976), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U952 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U954 ( .A1(n878), .A2(G124), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G112), .A2(n879), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G100), .A2(n886), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G136), .A2(n883), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U961 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U962 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n862) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U965 ( .A(G164), .B(G162), .Z(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n877) );
  NAND2_X1 U968 ( .A1(G130), .A2(n878), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G118), .A2(n879), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U971 ( .A1(n886), .A2(G106), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT112), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G142), .A2(n883), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(KEYINPUT45), .B(n872), .Z(n873) );
  NOR2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n924), .B(n875), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n895) );
  NAND2_X1 U979 ( .A1(G127), .A2(n878), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G115), .A2(n879), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n882), .B(KEYINPUT47), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G139), .A2(n883), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n889) );
  NAND2_X1 U985 ( .A1(G103), .A2(n886), .ZN(n887) );
  XNOR2_X1 U986 ( .A(KEYINPUT113), .B(n887), .ZN(n888) );
  NOR2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n910) );
  XNOR2_X1 U988 ( .A(n890), .B(n910), .ZN(n893) );
  XOR2_X1 U989 ( .A(G160), .B(n891), .Z(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U991 ( .A(n895), .B(n894), .Z(n896) );
  NOR2_X1 U992 ( .A1(G37), .A2(n896), .ZN(G395) );
  INV_X1 U993 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U994 ( .A(n960), .B(n897), .ZN(n899) );
  XOR2_X1 U995 ( .A(G301), .B(n964), .Z(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(G286), .B(n900), .Z(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n902), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n903), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n904) );
  AND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n906), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(KEYINPUT116), .B(n907), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  INV_X1 U1008 ( .A(KEYINPUT55), .ZN(n934) );
  NAND2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n923) );
  XNOR2_X1 U1010 ( .A(G164), .B(G2078), .ZN(n913) );
  XOR2_X1 U1011 ( .A(G2072), .B(n910), .Z(n911) );
  XNOR2_X1 U1012 ( .A(KEYINPUT117), .B(n911), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n914), .B(KEYINPUT50), .ZN(n919) );
  XOR2_X1 U1015 ( .A(G2090), .B(G162), .Z(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n917), .B(KEYINPUT51), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n929) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT52), .B(n930), .ZN(n931) );
  XOR2_X1 U1026 ( .A(KEYINPUT118), .B(n931), .Z(n932) );
  NAND2_X1 U1027 ( .A1(n934), .A2(n932), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n933), .A2(G29), .ZN(n1014) );
  XNOR2_X1 U1029 ( .A(n934), .B(KEYINPUT121), .ZN(n954) );
  XNOR2_X1 U1030 ( .A(G2090), .B(G35), .ZN(n948) );
  XNOR2_X1 U1031 ( .A(G1996), .B(G32), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G1991), .B(G25), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1034 ( .A(G2072), .B(G33), .Z(n937) );
  NAND2_X1 U1035 ( .A1(n937), .A2(G28), .ZN(n940) );
  XOR2_X1 U1036 ( .A(KEYINPUT119), .B(G2067), .Z(n938) );
  XNOR2_X1 U1037 ( .A(G26), .B(n938), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1040 ( .A(G27), .B(n943), .Z(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT53), .B(n946), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n952) );
  XOR2_X1 U1044 ( .A(KEYINPUT120), .B(G34), .Z(n950) );
  XNOR2_X1 U1045 ( .A(G2084), .B(KEYINPUT54), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(n950), .B(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n954), .B(n953), .ZN(n955) );
  OR2_X1 U1049 ( .A1(G29), .A2(n955), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(G11), .A2(n956), .ZN(n1012) );
  INV_X1 U1051 ( .A(G16), .ZN(n1008) );
  XOR2_X1 U1052 ( .A(n1008), .B(KEYINPUT56), .Z(n983) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G168), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT57), .B(n959), .ZN(n981) );
  XNOR2_X1 U1056 ( .A(G1341), .B(KEYINPUT123), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(n960), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n976) );
  XOR2_X1 U1060 ( .A(G1348), .B(n964), .Z(n966) );
  XNOR2_X1 U1061 ( .A(G301), .B(G1961), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(KEYINPUT122), .B(n967), .ZN(n974) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1065 ( .A(G1956), .B(n970), .Z(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1070 ( .A(KEYINPUT124), .B(n979), .Z(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n1010) );
  XOR2_X1 U1073 ( .A(KEYINPUT126), .B(G4), .Z(n985) );
  XNOR2_X1 U1074 ( .A(G1348), .B(KEYINPUT59), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n985), .B(n984), .ZN(n992) );
  XOR2_X1 U1076 ( .A(G1341), .B(G19), .Z(n989) );
  XNOR2_X1 U1077 ( .A(G1981), .B(G6), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(G20), .B(G1956), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1081 ( .A(KEYINPUT125), .B(n990), .Z(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n993), .ZN(n995) );
  XOR2_X1 U1084 ( .A(G1961), .B(G5), .Z(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1005) );
  XOR2_X1 U1086 ( .A(G1966), .B(G21), .Z(n1003) );
  XNOR2_X1 U1087 ( .A(G1986), .B(G24), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G1976), .B(G23), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(G22), .B(G1971), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT127), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT58), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1015), .ZN(G150) );
  INV_X1 U1102 ( .A(G150), .ZN(G311) );
endmodule

