

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U318 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U319 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n429) );
  XNOR2_X1 U320 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U321 ( .A(n304), .B(n303), .ZN(n308) );
  XNOR2_X1 U322 ( .A(n432), .B(KEYINPUT55), .ZN(n449) );
  INV_X1 U323 ( .A(G190GAT), .ZN(n450) );
  XNOR2_X1 U324 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U325 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U326 ( .A(KEYINPUT10), .B(G92GAT), .Z(n287) );
  XNOR2_X1 U327 ( .A(G162GAT), .B(G218GAT), .ZN(n286) );
  XNOR2_X1 U328 ( .A(n287), .B(n286), .ZN(n290) );
  INV_X1 U329 ( .A(n290), .ZN(n288) );
  XOR2_X1 U330 ( .A(G29GAT), .B(G134GAT), .Z(n335) );
  NAND2_X1 U331 ( .A1(n288), .A2(n335), .ZN(n292) );
  INV_X1 U332 ( .A(n335), .ZN(n289) );
  NAND2_X1 U333 ( .A1(n290), .A2(n289), .ZN(n291) );
  NAND2_X1 U334 ( .A1(n292), .A2(n291), .ZN(n294) );
  NAND2_X1 U335 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n296) );
  INV_X1 U337 ( .A(KEYINPUT9), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n304) );
  XOR2_X1 U339 ( .A(G43GAT), .B(G50GAT), .Z(n298) );
  XNOR2_X1 U340 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n392) );
  XNOR2_X1 U342 ( .A(n392), .B(KEYINPUT11), .ZN(n302) );
  XOR2_X1 U343 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n300) );
  XNOR2_X1 U344 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n299) );
  XOR2_X1 U345 ( .A(n300), .B(n299), .Z(n301) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(G85GAT), .ZN(n305) );
  XNOR2_X1 U347 ( .A(n305), .B(KEYINPUT72), .ZN(n367) );
  XNOR2_X1 U348 ( .A(G36GAT), .B(G190GAT), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n306), .B(KEYINPUT77), .ZN(n421) );
  XNOR2_X1 U350 ( .A(n367), .B(n421), .ZN(n307) );
  XOR2_X1 U351 ( .A(n308), .B(n307), .Z(n538) );
  INV_X1 U352 ( .A(n538), .ZN(n552) );
  XOR2_X1 U353 ( .A(G204GAT), .B(KEYINPUT23), .Z(n310) );
  XNOR2_X1 U354 ( .A(G50GAT), .B(KEYINPUT24), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U356 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n312) );
  XNOR2_X1 U357 ( .A(G22GAT), .B(KEYINPUT85), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U359 ( .A(n314), .B(n313), .Z(n324) );
  XNOR2_X1 U360 ( .A(G211GAT), .B(KEYINPUT86), .ZN(n315) );
  XNOR2_X1 U361 ( .A(n315), .B(KEYINPUT21), .ZN(n316) );
  XOR2_X1 U362 ( .A(n316), .B(KEYINPUT87), .Z(n318) );
  XNOR2_X1 U363 ( .A(G197GAT), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n318), .B(n317), .ZN(n418) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(G78GAT), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n319), .B(KEYINPUT71), .ZN(n368) );
  XOR2_X1 U367 ( .A(n368), .B(G148GAT), .Z(n321) );
  NAND2_X1 U368 ( .A1(G228GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n418), .B(n322), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U372 ( .A(KEYINPUT3), .B(G162GAT), .Z(n326) );
  XNOR2_X1 U373 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U375 ( .A(G141GAT), .B(n327), .ZN(n345) );
  XNOR2_X1 U376 ( .A(n328), .B(n345), .ZN(n462) );
  XOR2_X1 U377 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n330) );
  XNOR2_X1 U378 ( .A(G85GAT), .B(KEYINPUT91), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U380 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n332) );
  XNOR2_X1 U381 ( .A(KEYINPUT6), .B(KEYINPUT88), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U383 ( .A(n334), .B(n333), .Z(n340) );
  XOR2_X1 U384 ( .A(G113GAT), .B(KEYINPUT0), .Z(n436) );
  XOR2_X1 U385 ( .A(G1GAT), .B(G127GAT), .Z(n351) );
  XOR2_X1 U386 ( .A(n351), .B(n335), .Z(n337) );
  NAND2_X1 U387 ( .A1(G225GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n436), .B(n338), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(n341), .B(KEYINPUT92), .Z(n344) );
  XNOR2_X1 U392 ( .A(G120GAT), .B(G148GAT), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n342), .B(G57GAT), .ZN(n374) );
  XNOR2_X1 U394 ( .A(n374), .B(KEYINPUT4), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n346), .B(n345), .ZN(n461) );
  XNOR2_X1 U397 ( .A(KEYINPUT93), .B(n461), .ZN(n513) );
  XOR2_X1 U398 ( .A(KEYINPUT116), .B(KEYINPUT48), .Z(n413) );
  XOR2_X1 U399 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n348) );
  XNOR2_X1 U400 ( .A(G211GAT), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n365) );
  XOR2_X1 U402 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n350) );
  XNOR2_X1 U403 ( .A(G64GAT), .B(G57GAT), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n355) );
  XOR2_X1 U405 ( .A(G71GAT), .B(KEYINPUT13), .Z(n378) );
  XOR2_X1 U406 ( .A(n351), .B(n378), .Z(n353) );
  XNOR2_X1 U407 ( .A(G183GAT), .B(G155GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U409 ( .A(n355), .B(n354), .Z(n357) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n359) );
  INV_X1 U412 ( .A(KEYINPUT15), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U414 ( .A(G8GAT), .B(KEYINPUT68), .Z(n361) );
  XNOR2_X1 U415 ( .A(G15GAT), .B(G22GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n391) );
  XNOR2_X1 U417 ( .A(n391), .B(KEYINPUT78), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n535) );
  INV_X1 U420 ( .A(n535), .ZN(n573) );
  XOR2_X1 U421 ( .A(KEYINPUT36), .B(n538), .Z(n576) );
  NOR2_X1 U422 ( .A1(n573), .A2(n576), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n366), .B(KEYINPUT45), .ZN(n383) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n382) );
  XOR2_X1 U425 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n370) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U428 ( .A(n371), .B(KEYINPUT31), .Z(n376) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G92GAT), .Z(n373) );
  XNOR2_X1 U430 ( .A(G176GAT), .B(G204GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n423) );
  XNOR2_X1 U432 ( .A(n423), .B(n374), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U434 ( .A(n377), .B(KEYINPUT73), .Z(n380) );
  XNOR2_X1 U435 ( .A(n378), .B(KEYINPUT32), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n569) );
  NAND2_X1 U438 ( .A1(n383), .A2(n569), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n384), .B(KEYINPUT115), .ZN(n403) );
  XOR2_X1 U440 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n386) );
  XNOR2_X1 U441 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n402) );
  XOR2_X1 U443 ( .A(G197GAT), .B(G141GAT), .Z(n388) );
  XNOR2_X1 U444 ( .A(G169GAT), .B(G113GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n390) );
  XOR2_X1 U446 ( .A(G29GAT), .B(G36GAT), .Z(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n398) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U449 ( .A(KEYINPUT29), .B(KEYINPUT64), .Z(n394) );
  XNOR2_X1 U450 ( .A(KEYINPUT65), .B(KEYINPUT30), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n400) );
  NAND2_X1 U454 ( .A1(G229GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n529) );
  INV_X1 U457 ( .A(n529), .ZN(n564) );
  NAND2_X1 U458 ( .A1(n403), .A2(n564), .ZN(n411) );
  XOR2_X1 U459 ( .A(KEYINPUT47), .B(KEYINPUT114), .Z(n409) );
  XNOR2_X1 U460 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n405) );
  XOR2_X1 U461 ( .A(n569), .B(KEYINPUT41), .Z(n555) );
  INV_X1 U462 ( .A(n555), .ZN(n531) );
  NAND2_X1 U463 ( .A1(n529), .A2(n531), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  NOR2_X1 U465 ( .A1(n535), .A2(n406), .ZN(n407) );
  NAND2_X1 U466 ( .A1(n407), .A2(n552), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n410) );
  NAND2_X1 U468 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n524) );
  XNOR2_X1 U470 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n414), .B(KEYINPUT17), .ZN(n415) );
  XOR2_X1 U472 ( .A(n415), .B(KEYINPUT83), .Z(n417) );
  XNOR2_X1 U473 ( .A(G169GAT), .B(G183GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n446) );
  XNOR2_X1 U475 ( .A(n446), .B(n418), .ZN(n427) );
  XOR2_X1 U476 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n420) );
  NAND2_X1 U477 ( .A1(G226GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n425) );
  XNOR2_X1 U480 ( .A(G8GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U482 ( .A(n427), .B(n426), .Z(n516) );
  XOR2_X1 U483 ( .A(n516), .B(KEYINPUT122), .Z(n428) );
  NOR2_X1 U484 ( .A1(n524), .A2(n428), .ZN(n430) );
  NOR2_X1 U485 ( .A1(n513), .A2(n431), .ZN(n562) );
  NAND2_X1 U486 ( .A1(n462), .A2(n562), .ZN(n432) );
  XOR2_X1 U487 ( .A(G190GAT), .B(G134GAT), .Z(n434) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(G99GAT), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U493 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n440) );
  XNOR2_X1 U494 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n448) );
  XOR2_X1 U497 ( .A(G176GAT), .B(G127GAT), .Z(n444) );
  XNOR2_X1 U498 ( .A(G15GAT), .B(G120GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U501 ( .A(n448), .B(n447), .Z(n464) );
  INV_X1 U502 ( .A(n464), .ZN(n525) );
  NAND2_X1 U503 ( .A1(n449), .A2(n525), .ZN(n559) );
  NOR2_X1 U504 ( .A1(n552), .A2(n559), .ZN(n453) );
  XNOR2_X1 U505 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n451) );
  XOR2_X1 U506 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n470) );
  NAND2_X1 U507 ( .A1(n569), .A2(n529), .ZN(n485) );
  NOR2_X1 U508 ( .A1(n573), .A2(n538), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n454), .B(KEYINPUT16), .ZN(n468) );
  NAND2_X1 U510 ( .A1(n525), .A2(n516), .ZN(n455) );
  NAND2_X1 U511 ( .A1(n462), .A2(n455), .ZN(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT25), .B(n456), .Z(n459) );
  XNOR2_X1 U513 ( .A(n516), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U514 ( .A1(n462), .A2(n525), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n457), .B(KEYINPUT26), .ZN(n561) );
  NAND2_X1 U516 ( .A1(n463), .A2(n561), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n461), .A2(n460), .ZN(n467) );
  XOR2_X1 U519 ( .A(n462), .B(KEYINPUT28), .Z(n527) );
  NAND2_X1 U520 ( .A1(n463), .A2(n513), .ZN(n523) );
  NOR2_X1 U521 ( .A1(n527), .A2(n523), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n481) );
  NAND2_X1 U524 ( .A1(n468), .A2(n481), .ZN(n499) );
  NOR2_X1 U525 ( .A1(n485), .A2(n499), .ZN(n477) );
  NAND2_X1 U526 ( .A1(n477), .A2(n513), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U528 ( .A(G1GAT), .B(n471), .Z(G1324GAT) );
  NAND2_X1 U529 ( .A1(n516), .A2(n477), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n474) );
  NAND2_X1 U532 ( .A1(n477), .A2(n525), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n476) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT97), .Z(n475) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(G1326GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n479) );
  NAND2_X1 U537 ( .A1(n477), .A2(n527), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n480), .ZN(G1327GAT) );
  NAND2_X1 U540 ( .A1(n573), .A2(n481), .ZN(n482) );
  NOR2_X1 U541 ( .A1(n576), .A2(n482), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n512) );
  NOR2_X1 U544 ( .A1(n485), .A2(n512), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT38), .ZN(n495) );
  NAND2_X1 U546 ( .A1(n495), .A2(n513), .ZN(n490) );
  XOR2_X1 U547 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n488) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n495), .A2(n516), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U553 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n495), .A2(n525), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  XOR2_X1 U557 ( .A(G50GAT), .B(KEYINPUT105), .Z(n497) );
  NAND2_X1 U558 ( .A1(n527), .A2(n495), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n502) );
  NAND2_X1 U561 ( .A1(n531), .A2(n564), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT106), .ZN(n511) );
  NOR2_X1 U563 ( .A1(n511), .A2(n499), .ZN(n500) );
  XOR2_X1 U564 ( .A(KEYINPUT107), .B(n500), .Z(n507) );
  NAND2_X1 U565 ( .A1(n507), .A2(n513), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  NAND2_X1 U568 ( .A1(n516), .A2(n507), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U570 ( .A(G71GAT), .B(KEYINPUT109), .Z(n506) );
  NAND2_X1 U571 ( .A1(n507), .A2(n525), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U574 ( .A1(n507), .A2(n527), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  XOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT111), .Z(n515) );
  NOR2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n520), .A2(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n520), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(KEYINPUT112), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(n518), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n525), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n527), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n543) );
  NAND2_X1 U590 ( .A1(n525), .A2(n543), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(KEYINPUT117), .B(n528), .Z(n539) );
  NAND2_X1 U593 ( .A1(n539), .A2(n529), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U596 ( .A1(n539), .A2(n531), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n535), .A2(n539), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  NAND2_X1 U606 ( .A1(n543), .A2(n561), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n564), .A2(n551), .ZN(n544) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n548) );
  NOR2_X1 U612 ( .A1(n555), .A2(n551), .ZN(n547) );
  XOR2_X1 U613 ( .A(n548), .B(n547), .Z(G1345GAT) );
  NOR2_X1 U614 ( .A1(n573), .A2(n551), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NOR2_X1 U619 ( .A1(n564), .A2(n559), .ZN(n554) );
  XOR2_X1 U620 ( .A(G169GAT), .B(n554), .Z(G1348GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n559), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n573), .A2(n559), .ZN(n560) );
  XOR2_X1 U626 ( .A(G183GAT), .B(n560), .Z(G1350GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT125), .B(n563), .Z(n575) );
  NOR2_X1 U629 ( .A1(n564), .A2(n575), .ZN(n568) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT126), .B(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n575), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XOR2_X1 U639 ( .A(G211GAT), .B(n574), .Z(G1354GAT) );
  INV_X1 U640 ( .A(KEYINPUT62), .ZN(n578) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

