//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014;
  INV_X1    g000(.A(G134gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(G127gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G134gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G113gat), .B(G120gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(G113gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G120gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G127gat), .B(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n208), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(KEYINPUT2), .ZN(new_n224));
  XNOR2_X1  g023(.A(G141gat), .B(G148gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT74), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G141gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G148gat), .ZN(new_n229));
  INV_X1    g028(.A(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G141gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n231), .A3(new_n226), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n223), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT75), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n231), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n221), .B1(new_n220), .B2(KEYINPUT2), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n217), .B1(new_n241), .B2(KEYINPUT3), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n229), .A2(new_n231), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT74), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n232), .A3(new_n224), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n246), .A2(new_n223), .B1(new_n238), .B2(new_n239), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n243), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AND4_X1   g048(.A1(new_n243), .A2(new_n234), .A3(new_n248), .A4(new_n240), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n242), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n217), .A2(new_n234), .A3(new_n240), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT4), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(new_n255), .A3(new_n217), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT77), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT77), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n253), .B2(KEYINPUT4), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n251), .B(new_n252), .C1(new_n257), .C2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n208), .A2(new_n216), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(G155gat), .B2(G162gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n244), .B2(KEYINPUT74), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n222), .B1(new_n265), .B2(new_n232), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n238), .A2(new_n239), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n252), .B1(new_n268), .B2(new_n253), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n261), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n252), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n266), .A2(new_n267), .A3(new_n262), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n234), .A2(new_n240), .B1(new_n216), .B2(new_n208), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT5), .B1(new_n254), .B2(new_n256), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n251), .A2(new_n278), .A3(new_n252), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G1gat), .B(G29gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT0), .ZN(new_n283));
  XNOR2_X1  g082(.A(G57gat), .B(G85gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(KEYINPUT6), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT78), .B1(new_n275), .B2(KEYINPUT5), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n269), .A2(new_n261), .A3(new_n270), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n279), .B1(new_n291), .B2(new_n260), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n288), .B1(new_n292), .B2(new_n285), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n277), .A2(new_n285), .A3(new_n280), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n287), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G211gat), .A2(G218gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT22), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G197gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G204gat), .ZN(new_n303));
  INV_X1    g102(.A(G204gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G197gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n299), .B1(new_n298), .B2(new_n300), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n297), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n309), .A2(new_n296), .A3(new_n310), .A4(new_n301), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(KEYINPUT23), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n319), .A2(G169gat), .A3(G176gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT64), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(KEYINPUT23), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT64), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n319), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n316), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n327), .B(new_n328), .C1(G183gat), .C2(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n321), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n318), .A2(new_n331), .A3(new_n320), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n326), .B(KEYINPUT65), .ZN(new_n334));
  OR3_X1    g133(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n328), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n333), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  NOR3_X1   g139(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n317), .ZN(new_n344));
  NOR4_X1   g143(.A1(KEYINPUT69), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(KEYINPUT70), .B(new_n340), .C1(new_n344), .C2(new_n345), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT27), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n352));
  INV_X1    g151(.A(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(KEYINPUT67), .B2(G183gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT27), .B(G183gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT28), .A3(new_n353), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(new_n349), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n339), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n315), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n314), .B1(new_n339), .B2(new_n360), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n313), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n315), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n339), .B2(new_n360), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n366), .B(new_n312), .C1(new_n315), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n365), .A2(new_n372), .A3(new_n368), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n376));
  OR3_X1    g175(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n373), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n295), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT31), .B(G50gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n234), .A2(new_n248), .A3(new_n240), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT76), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n234), .A2(new_n243), .A3(new_n248), .A4(new_n240), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n388), .B2(new_n312), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n362), .B1(new_n249), .B2(new_n250), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT80), .A3(new_n313), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n312), .B2(new_n362), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT79), .B1(new_n392), .B2(new_n247), .ZN(new_n393));
  INV_X1    g192(.A(G228gat), .ZN(new_n394));
  INV_X1    g193(.A(G233gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n308), .B2(new_n311), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n241), .B(new_n397), .C1(new_n398), .C2(KEYINPUT3), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n393), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n389), .A2(new_n391), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G22gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n312), .B1(new_n403), .B2(new_n362), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n392), .A2(new_n247), .ZN(new_n405));
  OAI22_X1  g204(.A1(new_n404), .A2(new_n405), .B1(new_n394), .B2(new_n395), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n401), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n402), .B1(new_n401), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n383), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n401), .A2(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G22gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n401), .A2(new_n406), .A3(new_n402), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n382), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n379), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G15gat), .B(G43gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n339), .A2(new_n360), .A3(new_n217), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n217), .B1(new_n339), .B2(new_n360), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n418), .B1(new_n423), .B2(KEYINPUT32), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT32), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n348), .A2(new_n349), .A3(new_n359), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n334), .A2(new_n337), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n429), .A2(new_n333), .B1(new_n330), .B2(new_n331), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n262), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n339), .A2(new_n360), .A3(new_n217), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n433), .B2(new_n420), .ZN(new_n434));
  INV_X1    g233(.A(new_n418), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT33), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n424), .A2(new_n426), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n431), .A2(new_n419), .A3(new_n432), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT34), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n423), .A2(KEYINPUT32), .A3(new_n436), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n419), .B1(new_n431), .B2(new_n432), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n435), .B1(new_n443), .B2(new_n427), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(KEYINPUT33), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n438), .B(KEYINPUT34), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT36), .B1(new_n441), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n437), .B2(new_n440), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n446), .A2(KEYINPUT72), .A3(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT71), .B1(new_n446), .B2(new_n447), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n456), .A3(new_n440), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n453), .A2(new_n454), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n415), .A2(new_n449), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n287), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n285), .B1(new_n277), .B2(new_n280), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(KEYINPUT84), .A3(KEYINPUT6), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n375), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n365), .A2(new_n466), .A3(new_n368), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT37), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT37), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n365), .A2(new_n466), .A3(new_n368), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n373), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n465), .B1(new_n471), .B2(KEYINPUT38), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n281), .A2(new_n286), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n292), .A2(new_n285), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n288), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n468), .A2(new_n476), .A3(new_n373), .A4(new_n470), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n464), .A2(new_n472), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n409), .A2(new_n413), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n376), .A2(new_n377), .A3(new_n473), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n254), .A2(new_n256), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n251), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT81), .B1(new_n482), .B2(new_n272), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  AOI211_X1 g283(.A(new_n484), .B(new_n252), .C1(new_n251), .C2(new_n481), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT39), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n273), .A2(new_n274), .A3(new_n272), .ZN(new_n487));
  NOR4_X1   g286(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n403), .A2(new_n242), .B1(new_n254), .B2(new_n256), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n484), .B1(new_n490), .B2(new_n252), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(KEYINPUT81), .A3(new_n272), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT39), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n493), .B2(new_n286), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n486), .B1(new_n483), .B2(new_n485), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT82), .A3(new_n285), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n488), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n480), .B1(new_n497), .B2(KEYINPUT40), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  AOI211_X1 g298(.A(new_n499), .B(new_n488), .C1(new_n494), .C2(new_n496), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n478), .B(new_n479), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n441), .A2(new_n448), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n479), .A2(new_n502), .A3(new_n295), .A4(new_n378), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT35), .B1(new_n376), .B2(new_n377), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n479), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n437), .A2(new_n450), .A3(new_n440), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT72), .B1(new_n446), .B2(new_n447), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n455), .A2(new_n457), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n464), .A2(new_n475), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n459), .A2(new_n501), .B1(new_n504), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G230gat), .A2(G233gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  INV_X1    g315(.A(G85gat), .ZN(new_n517));
  INV_X1    g316(.A(G92gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(KEYINPUT91), .A2(G85gat), .A3(G92gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n519), .B(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT92), .B1(G99gat), .B2(G106gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(KEYINPUT92), .A2(G99gat), .A3(G106gat), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n525), .A2(new_n526), .B1(new_n517), .B2(new_n518), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G99gat), .B(G106gat), .Z(new_n529));
  OR2_X1    g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  OR2_X1    g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G64gat), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT89), .B1(new_n537), .B2(G57gat), .ZN(new_n538));
  INV_X1    g337(.A(G57gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(G64gat), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n537), .A2(KEYINPUT89), .A3(G57gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n537), .A2(G57gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n539), .A2(G64gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT9), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n545), .A2(new_n533), .A3(new_n534), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n547), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n549), .A3(new_n531), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n515), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n530), .A2(KEYINPUT10), .A3(new_n549), .A4(new_n531), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT95), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT10), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n555), .A3(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(KEYINPUT95), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT97), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n560), .A3(new_n515), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n559), .B2(new_n515), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n552), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G120gat), .B(G148gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT96), .ZN(new_n566));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(KEYINPUT98), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571));
  INV_X1    g370(.A(new_n554), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n548), .A2(new_n555), .A3(new_n550), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n515), .B(new_n572), .C1(new_n573), .C2(new_n557), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT97), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n551), .B1(new_n575), .B2(new_n561), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n571), .B1(new_n576), .B2(new_n568), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n568), .A3(new_n552), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT21), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n547), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G127gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G15gat), .B(G22gat), .ZN(new_n586));
  INV_X1    g385(.A(G1gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT16), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(G1gat), .B2(new_n586), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(G8gat), .Z(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT87), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(G8gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT87), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n581), .B2(new_n547), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n585), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n218), .ZN(new_n600));
  XOR2_X1   g399(.A(G183gat), .B(G211gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n532), .ZN(new_n607));
  XNOR2_X1  g406(.A(G43gat), .B(G50gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(KEYINPUT15), .ZN(new_n609));
  NOR2_X1   g408(.A1(G29gat), .A2(G36gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT14), .ZN(new_n611));
  INV_X1    g410(.A(G29gat), .ZN(new_n612));
  INV_X1    g411(.A(G36gat), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT86), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n609), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(KEYINPUT15), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n607), .A2(new_n619), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n617), .A2(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT17), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT17), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n532), .B(KEYINPUT93), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n626), .A2(KEYINPUT94), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT94), .B1(new_n626), .B2(new_n627), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n621), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G190gat), .B(G218gat), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n633), .B(new_n621), .C1(new_n628), .C2(new_n629), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT90), .ZN(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n632), .A2(new_n639), .A3(new_n634), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n580), .A2(new_n606), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n619), .B1(new_n592), .B2(new_n595), .ZN(new_n645));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n625), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n593), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT18), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n596), .A2(new_n622), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n645), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n646), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n648), .A2(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G113gat), .B(G141gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G169gat), .B(G197gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT12), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n650), .A2(new_n655), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n514), .A2(new_n644), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n295), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  INV_X1    g470(.A(new_n378), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT99), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(G8gat), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND3_X1  g478(.A1(new_n674), .A2(KEYINPUT42), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(KEYINPUT100), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n675), .B2(new_n677), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n683), .A2(KEYINPUT101), .A3(KEYINPUT42), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n678), .B(new_n680), .C1(new_n686), .C2(new_n687), .ZN(G1325gat));
  INV_X1    g487(.A(G15gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n668), .A2(new_n689), .A3(new_n511), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n458), .A2(new_n449), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n668), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n692), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g492(.A1(new_n668), .A2(new_n414), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT102), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n514), .B2(new_n643), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n641), .A2(new_n642), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n415), .A2(new_n449), .A3(new_n458), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT84), .B1(new_n462), .B2(KEYINPUT6), .ZN(new_n702));
  NOR4_X1   g501(.A1(new_n292), .A2(new_n460), .A3(new_n288), .A4(new_n285), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n475), .B(new_n477), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n414), .B1(new_n705), .B2(new_n472), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n497), .A2(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n497), .A2(KEYINPUT40), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n480), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n701), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n479), .A2(new_n505), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n475), .B2(new_n464), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n712), .A2(new_n511), .B1(KEYINPUT35), .B2(new_n503), .ZN(new_n713));
  OAI211_X1 g512(.A(KEYINPUT44), .B(new_n700), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n606), .B(KEYINPUT103), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n578), .A2(new_n579), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n716), .A2(new_n667), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n699), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n699), .A2(new_n714), .A3(KEYINPUT104), .A4(new_n718), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n669), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n612), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n724), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n514), .A2(new_n667), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n643), .A2(new_n717), .A3(new_n606), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(G29gat), .A3(new_n295), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT45), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n726), .A2(new_n731), .ZN(G1328gat));
  NOR3_X1   g531(.A1(new_n729), .A2(G36gat), .A3(new_n378), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n721), .A2(new_n672), .A3(new_n722), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n613), .B2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n691), .ZN(new_n737));
  OAI21_X1  g536(.A(G43gat), .B1(new_n719), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n511), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(G43gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n738), .B(KEYINPUT47), .C1(new_n729), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n729), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n721), .A2(new_n691), .A3(new_n722), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(G43gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT107), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n749), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1330gat));
  INV_X1    g550(.A(G50gat), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n727), .A2(new_n752), .A3(new_n414), .A4(new_n728), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT48), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n699), .A2(new_n714), .A3(new_n414), .A4(new_n718), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n755), .B2(KEYINPUT108), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  INV_X1    g560(.A(new_n753), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n721), .A2(new_n414), .A3(new_n722), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(G50gat), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n760), .A2(new_n761), .B1(KEYINPUT48), .B2(new_n764), .ZN(G1331gat));
  INV_X1    g564(.A(new_n606), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n700), .A2(new_n766), .A3(new_n666), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n717), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT110), .ZN(new_n769));
  INV_X1    g568(.A(new_n514), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n295), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n539), .ZN(G1332gat));
  NOR2_X1   g572(.A1(new_n771), .A2(new_n378), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  AND2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(G1333gat));
  NOR3_X1   g577(.A1(new_n771), .A2(G71gat), .A3(new_n739), .ZN(new_n779));
  INV_X1    g578(.A(new_n771), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n691), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(G71gat), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n414), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g584(.A(KEYINPUT112), .B1(new_n514), .B2(new_n643), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n787), .B(new_n700), .C1(new_n710), .C2(new_n713), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n667), .A2(new_n766), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT111), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n580), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n517), .A3(new_n669), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n699), .A2(new_n714), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n790), .A2(new_n717), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n797), .A2(new_n669), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n517), .B2(new_n799), .ZN(G1336gat));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n791), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n792), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n791), .A2(new_n801), .A3(KEYINPUT51), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n378), .A2(G92gat), .ZN(new_n805));
  AND4_X1   g604(.A1(new_n717), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n797), .A2(new_n672), .A3(new_n798), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n795), .A2(new_n805), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n808), .A2(KEYINPUT52), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(G1337gat));
  NOR2_X1   g611(.A1(new_n580), .A2(new_n739), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(G99gat), .ZN(new_n815));
  INV_X1    g614(.A(new_n794), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n791), .A2(new_n792), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n691), .A3(new_n798), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G99gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT114), .ZN(G1338gat));
  AND3_X1   g621(.A1(new_n791), .A2(new_n801), .A3(KEYINPUT51), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT51), .B1(new_n791), .B2(new_n801), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n580), .A2(G106gat), .A3(new_n479), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT115), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n798), .A2(new_n699), .A3(new_n414), .A4(new_n714), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G106gat), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT53), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n826), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n816), .B2(new_n817), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n829), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(KEYINPUT116), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n803), .A2(new_n804), .A3(new_n832), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n834), .B1(new_n838), .B2(new_n829), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n829), .A2(new_n834), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n793), .A2(new_n794), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n832), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n837), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n836), .A2(new_n843), .ZN(G1339gat));
  NOR2_X1   g643(.A1(new_n672), .A2(new_n295), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n626), .A2(new_n591), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n646), .B1(new_n847), .B2(new_n645), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n652), .A2(new_n654), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n661), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n665), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n717), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n559), .A2(new_n515), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n559), .B2(new_n515), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n568), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n575), .A2(new_n561), .A3(new_n855), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT55), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n579), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT55), .B1(new_n857), .B2(new_n858), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n666), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n700), .B1(new_n853), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n700), .A2(new_n861), .A3(new_n852), .A4(new_n863), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n715), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n767), .A2(new_n580), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(KEYINPUT117), .A3(new_n479), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872));
  INV_X1    g671(.A(new_n869), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n667), .A2(new_n860), .A3(new_n862), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n851), .B1(new_n578), .B2(new_n579), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n643), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n866), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n873), .B1(new_n877), .B2(new_n715), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n872), .B1(new_n878), .B2(new_n414), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n846), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n511), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n211), .A3(new_n667), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n878), .A2(new_n295), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n479), .A2(new_n502), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n672), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(G113gat), .B1(new_n886), .B2(new_n666), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n882), .A2(new_n887), .ZN(G1340gat));
  AOI21_X1  g687(.A(G120gat), .B1(new_n886), .B2(new_n717), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n814), .A2(new_n209), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n880), .B2(new_n890), .ZN(G1341gat));
  OAI21_X1  g690(.A(G127gat), .B1(new_n881), .B2(new_n715), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n204), .A3(new_n606), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1342gat));
  NAND4_X1  g693(.A1(new_n883), .A2(new_n202), .A3(new_n700), .A4(new_n885), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT56), .Z(new_n896));
  OAI21_X1  g695(.A(G134gat), .B1(new_n881), .B2(new_n643), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1343gat));
  NOR3_X1   g697(.A1(new_n691), .A2(new_n672), .A3(new_n479), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n666), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n900), .A2(new_n228), .B1(KEYINPUT119), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n691), .A2(new_n846), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n667), .A2(new_n228), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n479), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n766), .B1(new_n865), .B2(new_n867), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n873), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n606), .B1(new_n876), .B2(new_n866), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT118), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n907), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n479), .B1(new_n868), .B2(new_n869), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n903), .B(new_n904), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT119), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n902), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n902), .B2(new_n916), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1344gat));
  OAI211_X1 g719(.A(new_n717), .B(new_n903), .C1(new_n913), .C2(new_n915), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n922), .A3(G148gat), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n905), .B(new_n414), .C1(new_n911), .C2(new_n873), .ZN(new_n925));
  INV_X1    g724(.A(new_n903), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n580), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n925), .B(new_n927), .C1(new_n914), .C2(new_n905), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G148gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n924), .B1(new_n929), .B2(KEYINPUT59), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT120), .B(new_n922), .C1(new_n928), .C2(G148gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n883), .A2(new_n899), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n230), .A3(new_n717), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1345gat));
  NAND3_X1  g734(.A1(new_n933), .A2(new_n218), .A3(new_n606), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n913), .A2(new_n915), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n715), .A3(new_n926), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n938), .B2(new_n218), .ZN(G1346gat));
  AOI21_X1  g738(.A(G162gat), .B1(new_n933), .B2(new_n700), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n937), .A2(new_n926), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n643), .A2(new_n219), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n884), .A2(new_n378), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n870), .B2(new_n295), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n878), .A2(KEYINPUT121), .A3(new_n669), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT122), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n870), .A2(new_n945), .A3(new_n295), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT121), .B1(new_n878), .B2(new_n669), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n944), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n949), .A2(new_n666), .A3(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(G169gat), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n669), .A2(new_n378), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n511), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n958), .B1(new_n871), .B2(new_n879), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n667), .A2(new_n956), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n955), .A2(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1348gat));
  NAND3_X1  g760(.A1(new_n949), .A2(new_n717), .A3(new_n954), .ZN(new_n962));
  INV_X1    g761(.A(G176gat), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n580), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g763(.A1(new_n962), .A2(new_n963), .B1(new_n959), .B2(new_n964), .ZN(G1349gat));
  INV_X1    g764(.A(KEYINPUT60), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n952), .A2(new_n357), .A3(new_n606), .A4(new_n944), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n959), .A2(new_n716), .ZN(new_n968));
  INV_X1    g767(.A(G183gat), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n966), .B(new_n967), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n959), .B2(new_n716), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n606), .A2(new_n357), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n948), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT60), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n970), .A2(new_n974), .ZN(G1350gat));
  NAND4_X1  g774(.A1(new_n949), .A2(new_n353), .A3(new_n700), .A4(new_n954), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n700), .ZN(new_n977));
  XNOR2_X1  g776(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n977), .A2(G190gat), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n977), .B2(G190gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(G1351gat));
  OAI21_X1  g780(.A(KEYINPUT57), .B1(new_n878), .B2(new_n479), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(new_n925), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n982), .A2(KEYINPUT125), .A3(new_n925), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n737), .A2(new_n957), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n988), .A2(new_n302), .A3(new_n667), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n691), .A2(new_n378), .A3(new_n479), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n952), .A2(new_n666), .A3(new_n991), .ZN(new_n992));
  AOI22_X1  g791(.A1(new_n987), .A2(new_n989), .B1(new_n302), .B2(new_n992), .ZN(G1352gat));
  NAND4_X1  g792(.A1(new_n952), .A2(new_n304), .A3(new_n717), .A4(new_n991), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n996));
  INV_X1    g795(.A(new_n988), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(new_n717), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n998), .B1(new_n985), .B2(new_n986), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n995), .B(new_n996), .C1(new_n304), .C2(new_n999), .ZN(G1353gat));
  NAND4_X1  g799(.A1(new_n982), .A2(new_n606), .A3(new_n925), .A4(new_n997), .ZN(new_n1001));
  AND3_X1   g800(.A1(new_n1001), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(KEYINPUT63), .B1(new_n1001), .B2(G211gat), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n952), .A2(new_n991), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n766), .A2(G211gat), .ZN(new_n1005));
  OAI22_X1  g804(.A1(new_n1002), .A2(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(G1354gat));
  NAND3_X1  g805(.A1(new_n952), .A2(new_n700), .A3(new_n991), .ZN(new_n1007));
  INV_X1    g806(.A(G218gat), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n1007), .A2(KEYINPUT126), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g808(.A(KEYINPUT126), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n700), .A2(G218gat), .ZN(new_n1011));
  XOR2_X1   g810(.A(new_n1011), .B(KEYINPUT127), .Z(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(new_n997), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1013), .B1(new_n985), .B2(new_n986), .ZN(new_n1014));
  NOR3_X1   g813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1014), .ZN(G1355gat));
endmodule


