//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n203), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n207), .A2(KEYINPUT89), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT89), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n215), .A2(new_n204), .A3(new_n205), .A4(new_n206), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n208), .A3(new_n216), .ZN(new_n217));
  AOI211_X1 g016(.A(new_n213), .B(new_n210), .C1(new_n217), .C2(new_n211), .ZN(new_n218));
  NOR3_X1   g017(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n208), .B1(new_n219), .B2(new_n215), .ZN(new_n220));
  INV_X1    g019(.A(new_n216), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n211), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n210), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT90), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n212), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(G1gat), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n230), .B1(new_n229), .B2(new_n232), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(KEYINPUT17), .B(new_n212), .C1(new_n218), .C2(new_n224), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n227), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n235), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n225), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT92), .B1(new_n225), .B2(new_n239), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n218), .A2(new_n224), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT92), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n212), .A4(new_n235), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n247), .A3(new_n240), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n238), .B(KEYINPUT91), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT13), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n238), .A4(new_n240), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n243), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G197gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT11), .ZN(new_n256));
  INV_X1    g055(.A(G169gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n259), .A2(new_n243), .A3(new_n251), .A4(new_n252), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n269), .B2(new_n270), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n267), .B(new_n268), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT25), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  INV_X1    g075(.A(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n278), .B2(KEYINPUT26), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(KEYINPUT26), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n265), .A2(KEYINPUT67), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n279), .A2(new_n268), .A3(new_n280), .A4(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT27), .B(G183gat), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT28), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n289), .A3(new_n285), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n283), .A2(new_n287), .A3(new_n288), .A4(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n266), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT25), .B1(new_n294), .B2(new_n257), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n266), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT64), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n288), .B2(new_n270), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n288), .A2(new_n270), .ZN(new_n299));
  NAND4_X1  g098(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n298), .A2(new_n272), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n295), .A2(new_n268), .A3(new_n296), .A4(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n275), .A2(new_n291), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT68), .B(G120gat), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n305), .B1(G113gat), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n306), .B2(G113gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(G113gat), .B2(G120gat), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n307), .A2(new_n310), .B1(new_n305), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G227gat), .ZN(new_n315));
  INV_X1    g114(.A(G233gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n305), .A2(new_n312), .ZN(new_n318));
  INV_X1    g117(.A(new_n306), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n304), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n321), .B2(new_n309), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n275), .A2(new_n322), .A3(new_n291), .A4(new_n302), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n314), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n314), .A2(new_n326), .A3(new_n317), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT32), .ZN(new_n329));
  XNOR2_X1  g128(.A(G15gat), .B(G43gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G71gat), .ZN(new_n331));
  INV_X1    g130(.A(G99gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT33), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT70), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT70), .ZN(new_n336));
  AOI211_X1 g135(.A(new_n336), .B(KEYINPUT33), .C1(new_n325), .C2(new_n327), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n329), .B(new_n333), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(KEYINPUT33), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n328), .A2(KEYINPUT32), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n314), .A2(new_n323), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n315), .B2(new_n316), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT71), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT34), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(KEYINPUT72), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT34), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n351), .A3(new_n340), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G228gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(new_n316), .ZN(new_n357));
  INV_X1    g156(.A(G218gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT22), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT73), .B(G218gat), .ZN(new_n360));
  INV_X1    g159(.A(G211gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n362), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n358), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G211gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n362), .A2(new_n361), .A3(new_n363), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(G218gat), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT3), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G155gat), .B(G162gat), .Z(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT80), .B(G155gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT81), .B(G162gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n374), .B1(new_n377), .B2(KEYINPUT2), .ZN(new_n378));
  XNOR2_X1  g177(.A(G141gat), .B(G148gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT79), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n378), .A2(new_n380), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n373), .A2(new_n383), .B1(new_n371), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n357), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n357), .ZN(new_n389));
  INV_X1    g188(.A(new_n383), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n364), .A2(new_n365), .A3(new_n358), .ZN(new_n392));
  AOI21_X1  g191(.A(G218gat), .B1(new_n368), .B2(new_n369), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n391), .B(new_n372), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n384), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n366), .B2(new_n370), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n391), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n385), .A2(KEYINPUT85), .ZN(new_n399));
  INV_X1    g198(.A(new_n371), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT85), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n389), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n372), .B1(new_n392), .B2(new_n393), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n383), .B1(new_n404), .B2(new_n384), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n371), .A2(new_n385), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT83), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n388), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  OAI21_X1  g208(.A(G22gat), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G78gat), .B(G106gat), .Z(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT31), .B(G50gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(new_n408), .B2(new_n409), .ZN(new_n415));
  INV_X1    g214(.A(new_n402), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT3), .B1(new_n396), .B2(new_n391), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n404), .A2(KEYINPUT84), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n383), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n407), .B(new_n357), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n388), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G22gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(KEYINPUT86), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n410), .A2(new_n415), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n413), .B1(new_n422), .B2(KEYINPUT86), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n422), .B2(KEYINPUT86), .ZN(new_n427));
  AOI211_X1 g226(.A(new_n409), .B(G22gat), .C1(new_n420), .C2(new_n421), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AND4_X1   g228(.A1(KEYINPUT35), .A2(new_n355), .A3(new_n425), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT74), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n303), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G226gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n316), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n275), .A2(new_n291), .A3(new_n302), .A4(KEYINPUT74), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n434), .A2(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n303), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n400), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT75), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n432), .A2(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n437), .ZN(new_n442));
  INV_X1    g241(.A(new_n434), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n442), .B(new_n400), .C1(new_n443), .C2(new_n303), .ZN(new_n444));
  XOR2_X1   g243(.A(G64gat), .B(G92gat), .Z(new_n445));
  XNOR2_X1  g244(.A(G8gat), .B(G36gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n440), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n438), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n371), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT75), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT75), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n444), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n449), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n451), .A2(new_n458), .A3(KEYINPUT30), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n457), .A2(KEYINPUT30), .A3(new_n449), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT0), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(G57gat), .ZN(new_n464));
  INV_X1    g263(.A(G85gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n383), .A2(new_n313), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT4), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT4), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n383), .A2(new_n470), .A3(new_n313), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n313), .B1(new_n383), .B2(new_n384), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n390), .A2(new_n322), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n473), .B1(new_n478), .B2(new_n468), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n467), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n469), .A2(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT5), .B1(new_n482), .B2(new_n473), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n466), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n477), .A2(new_n467), .ZN(new_n485));
  INV_X1    g284(.A(new_n466), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n479), .B1(new_n482), .B2(new_n473), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n467), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n484), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n481), .A2(new_n483), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(new_n486), .C1(KEYINPUT82), .C2(KEYINPUT6), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n461), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n484), .A2(new_n488), .A3(new_n490), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n486), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n459), .A2(new_n460), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n355), .A2(new_n500), .A3(new_n429), .A4(new_n425), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n430), .A2(new_n496), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  INV_X1    g302(.A(new_n354), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n351), .B1(new_n338), .B2(new_n340), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n353), .A2(KEYINPUT36), .A3(new_n354), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n429), .A2(new_n425), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n495), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n449), .B1(new_n457), .B2(KEYINPUT37), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n440), .B2(new_n444), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT38), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n442), .B1(new_n443), .B2(new_n303), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n371), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n452), .B2(new_n371), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n436), .A2(KEYINPUT88), .A3(new_n400), .A4(new_n438), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT38), .B1(new_n520), .B2(KEYINPUT37), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n440), .A2(new_n512), .A3(new_n444), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n449), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n498), .A2(new_n499), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n514), .A2(new_n523), .A3(new_n524), .A4(new_n451), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n478), .A2(new_n473), .A3(new_n468), .ZN(new_n526));
  OAI211_X1 g325(.A(KEYINPUT39), .B(new_n526), .C1(new_n482), .C2(new_n473), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n472), .A2(new_n476), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT39), .ZN(new_n529));
  INV_X1    g328(.A(new_n473), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n531), .A2(new_n532), .A3(new_n466), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n531), .B2(new_n466), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT40), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n535), .A2(new_n536), .B1(new_n486), .B2(new_n492), .ZN(new_n537));
  OAI211_X1 g336(.A(KEYINPUT40), .B(new_n527), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n537), .A2(new_n459), .A3(new_n460), .A4(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n525), .A2(new_n539), .A3(new_n425), .A4(new_n429), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n508), .A2(new_n510), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n264), .B1(new_n502), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  OR2_X1    g342(.A1(G57gat), .A2(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(G57gat), .A2(G64gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G71gat), .B(G78gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n544), .B(new_n545), .C1(new_n552), .C2(KEYINPUT9), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n543), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G183gat), .B(G211gat), .Z(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n558), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n235), .B1(new_n557), .B2(new_n556), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT94), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT19), .ZN(new_n566));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT20), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n566), .A2(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n563), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n571), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n569), .A3(new_n562), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT7), .B1(new_n465), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(G85gat), .A3(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G99gat), .B(G106gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n465), .B2(new_n577), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n581), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n225), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n227), .A2(new_n236), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n587), .ZN(new_n591));
  XOR2_X1   g390(.A(G190gat), .B(G218gat), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G134gat), .B(G162gat), .Z(new_n595));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n594), .A2(KEYINPUT95), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n591), .A2(new_n593), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n591), .A2(new_n593), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n600), .A2(new_n601), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n581), .A2(new_n584), .ZN(new_n609));
  INV_X1    g408(.A(new_n582), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n553), .A2(new_n543), .A3(new_n549), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n549), .B1(new_n553), .B2(new_n543), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n551), .B(new_n554), .C1(new_n585), .C2(new_n586), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n587), .A2(new_n555), .A3(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT98), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT99), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n615), .A2(new_n616), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(G230gat), .A3(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n627));
  INV_X1    g426(.A(new_n622), .ZN(new_n628));
  AOI211_X1 g427(.A(new_n627), .B(new_n628), .C1(new_n618), .C2(new_n619), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n624), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n277), .ZN(new_n634));
  INV_X1    g433(.A(G204gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n631), .A2(new_n636), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n618), .A2(new_n619), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n639), .B1(new_n618), .B2(new_n619), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n621), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n636), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n626), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n637), .B1(new_n638), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n576), .A2(new_n608), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n542), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n494), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  INV_X1    g451(.A(new_n461), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n231), .A2(new_n230), .ZN(new_n654));
  NAND2_X1  g453(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n655));
  AND4_X1   g454(.A1(new_n653), .A2(new_n649), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n230), .B1(new_n649), .B2(new_n653), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT42), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(KEYINPUT42), .B2(new_n656), .ZN(G1325gat));
  AOI21_X1  g458(.A(G15gat), .B1(new_n649), .B2(new_n355), .ZN(new_n660));
  INV_X1    g459(.A(G15gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n508), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n660), .B1(new_n649), .B2(new_n663), .ZN(G1326gat));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n509), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NOR2_X1   g466(.A1(new_n576), .A2(new_n608), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n542), .A2(new_n646), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n205), .A3(new_n650), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  AOI211_X1 g471(.A(new_n672), .B(new_n608), .C1(new_n502), .C2(new_n541), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n510), .A2(KEYINPUT104), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n509), .A2(new_n675), .A3(new_n495), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n674), .A2(new_n508), .A3(new_n540), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n502), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n600), .A2(new_n601), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n607), .A2(new_n604), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n673), .B1(new_n672), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n261), .A2(KEYINPUT102), .A3(new_n262), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n261), .B2(new_n262), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n646), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n572), .A2(new_n574), .A3(KEYINPUT103), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT103), .B1(new_n572), .B2(new_n574), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n683), .A2(new_n688), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n494), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n671), .A2(new_n694), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n542), .A2(new_n653), .A3(new_n646), .A4(new_n668), .ZN(new_n697));
  OR3_X1    g496(.A1(new_n697), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT105), .B1(new_n697), .B2(G36gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n696), .B1(new_n700), .B2(KEYINPUT46), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n698), .A2(KEYINPUT106), .A3(new_n702), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(KEYINPUT46), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n693), .B2(new_n461), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n693), .B2(new_n508), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n709));
  INV_X1    g508(.A(G43gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n669), .A2(new_n710), .A3(new_n355), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n709), .B1(new_n708), .B2(new_n711), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(G1330gat));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n429), .A2(new_n425), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n717), .A2(KEYINPUT35), .A3(new_n496), .A4(new_n355), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n501), .A2(new_n497), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n508), .A2(new_n540), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n509), .A2(new_n675), .A3(new_n495), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n675), .B1(new_n509), .B2(new_n495), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n720), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n672), .B1(new_n725), .B2(new_n608), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n508), .A2(new_n510), .A3(new_n540), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT44), .B(new_n681), .C1(new_n727), .C2(new_n720), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n728), .A3(new_n692), .ZN(new_n729));
  INV_X1    g528(.A(new_n688), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n729), .A2(new_n717), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n716), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n669), .A2(new_n732), .A3(new_n509), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI221_X1 g536(.A(new_n734), .B1(new_n716), .B2(KEYINPUT48), .C1(new_n731), .C2(new_n732), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1331gat));
  AOI211_X1 g538(.A(new_n575), .B(new_n681), .C1(new_n677), .C2(new_n502), .ZN(new_n740));
  INV_X1    g539(.A(new_n686), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n646), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n650), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n461), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n743), .B2(new_n508), .ZN(new_n752));
  INV_X1    g551(.A(new_n355), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n753), .A2(G71gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n743), .B2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g555(.A1(new_n743), .A2(new_n717), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT109), .B(G78gat), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n576), .A2(new_n741), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n678), .A2(new_n681), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT51), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n608), .B1(new_n677), .B2(new_n502), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n764), .A3(new_n760), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n762), .A2(new_n687), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n465), .A3(new_n650), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n728), .B(new_n760), .C1(new_n763), .C2(KEYINPUT44), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n650), .A2(new_n687), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(G1336gat));
  NOR2_X1   g570(.A1(new_n461), .A2(G92gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n726), .A2(new_n687), .A3(new_n728), .A4(new_n760), .ZN(new_n775));
  OAI21_X1  g574(.A(G92gat), .B1(new_n775), .B2(new_n461), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n761), .B1(new_n779), .B2(KEYINPUT51), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n763), .A2(KEYINPUT110), .A3(new_n764), .A4(new_n760), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n780), .A2(new_n687), .A3(new_n772), .A4(new_n781), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n778), .B(new_n774), .C1(new_n776), .C2(new_n782), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n461), .A3(new_n646), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n784), .B2(new_n577), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT111), .B1(new_n785), .B2(KEYINPUT52), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n777), .B1(new_n783), .B2(new_n786), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n332), .A3(new_n355), .ZN(new_n788));
  OAI21_X1  g587(.A(G99gat), .B1(new_n775), .B2(new_n508), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  NOR2_X1   g589(.A1(new_n717), .A2(G106gat), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n780), .A2(new_n687), .A3(new_n781), .A4(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n768), .A2(new_n717), .A3(new_n646), .ZN(new_n793));
  INV_X1    g592(.A(G106gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT53), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n683), .A2(new_n509), .A3(new_n687), .A4(new_n760), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT53), .B1(new_n798), .B2(G106gat), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n762), .A2(new_n687), .A3(new_n765), .A4(new_n791), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n802), .B(new_n800), .C1(new_n793), .C2(new_n794), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(KEYINPUT112), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n796), .B1(new_n801), .B2(new_n804), .ZN(G1339gat));
  NOR2_X1   g604(.A1(new_n509), .A2(new_n753), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n618), .A2(new_n619), .A3(new_n628), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n623), .B2(new_n629), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n636), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n644), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n809), .A2(new_n636), .A3(new_n811), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n813), .A2(KEYINPUT113), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(new_n817), .A3(new_n644), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n816), .B(new_n818), .C1(new_n684), .C2(new_n685), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n248), .A2(new_n250), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n238), .B1(new_n237), .B2(new_n240), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n258), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n262), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n687), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n819), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n820), .B1(new_n819), .B2(new_n825), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n826), .A2(new_n827), .A3(new_n681), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n812), .A2(new_n817), .A3(new_n644), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n817), .B1(new_n812), .B2(new_n644), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n815), .A2(new_n814), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n824), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT114), .B1(new_n833), .B2(new_n608), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n681), .A2(new_n832), .A3(new_n835), .A4(new_n824), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n692), .B1(new_n828), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n647), .A2(new_n741), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n807), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n653), .A2(new_n494), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n264), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n741), .A2(new_n320), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(G1340gat));
  INV_X1    g645(.A(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n687), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(G120gat), .ZN(G1341gat));
  INV_X1    g648(.A(G127gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n843), .A2(new_n850), .A3(new_n692), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n576), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(G1342gat));
  AOI211_X1 g652(.A(new_n608), .B(new_n843), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n854));
  NOR2_X1   g653(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1343gat));
  NAND2_X1  g655(.A1(new_n508), .A2(new_n842), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n836), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n859));
  AND2_X1   g658(.A1(new_n815), .A2(new_n859), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n860), .A2(new_n813), .A3(KEYINPUT117), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT117), .B1(new_n860), .B2(new_n813), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n263), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n825), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n608), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n576), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n509), .B1(new_n866), .B2(new_n839), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n857), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n815), .A2(new_n814), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n818), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n825), .B1(new_n686), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT115), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n819), .A2(new_n820), .A3(new_n825), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n608), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n691), .B1(new_n876), .B2(new_n858), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n869), .B(new_n509), .C1(new_n877), .C2(new_n839), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n264), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n509), .B1(new_n877), .B2(new_n839), .ZN(new_n882));
  OR4_X1    g681(.A1(G141gat), .A2(new_n882), .A3(new_n264), .A4(new_n857), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n741), .A3(new_n878), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G141gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n883), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT118), .B1(new_n887), .B2(KEYINPUT58), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n889), .B(new_n881), .C1(new_n886), .C2(new_n883), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n884), .B1(new_n888), .B2(new_n890), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n838), .A2(new_n840), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n717), .A2(G148gat), .A3(new_n646), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n892), .A2(new_n508), .A3(new_n842), .A4(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n882), .A2(KEYINPUT57), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n681), .B1(new_n863), .B2(new_n825), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n833), .A2(new_n608), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n575), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n263), .B2(new_n647), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n869), .A3(new_n509), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n857), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n687), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n895), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n868), .A2(new_n687), .A3(new_n878), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(new_n895), .A3(G148gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n894), .B1(new_n905), .B2(new_n907), .ZN(G1345gat));
  AND2_X1   g707(.A1(new_n868), .A2(new_n878), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n691), .A2(new_n375), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT119), .Z(new_n911));
  INV_X1    g710(.A(new_n375), .ZN(new_n912));
  INV_X1    g711(.A(new_n882), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n576), .A3(new_n903), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n909), .A2(new_n911), .B1(new_n912), .B2(new_n914), .ZN(G1346gat));
  INV_X1    g714(.A(new_n376), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n879), .A2(new_n916), .A3(new_n608), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n681), .A3(new_n903), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n461), .A2(new_n650), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT121), .Z(new_n921));
  OAI211_X1 g720(.A(new_n806), .B(new_n921), .C1(new_n877), .C2(new_n839), .ZN(new_n922));
  OAI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n264), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n841), .A2(new_n920), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(G169gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n926), .B2(new_n741), .ZN(new_n927));
  NOR4_X1   g726(.A1(new_n925), .A2(KEYINPUT120), .A3(G169gat), .A4(new_n686), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n841), .A2(new_n687), .A3(new_n920), .ZN(new_n930));
  INV_X1    g729(.A(new_n922), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n687), .A2(new_n292), .A3(new_n293), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n930), .A2(new_n277), .B1(new_n931), .B2(new_n932), .ZN(G1349gat));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n841), .A2(KEYINPUT122), .A3(new_n691), .A4(new_n921), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n936), .B1(new_n922), .B2(new_n692), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n937), .A3(G183gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n841), .A2(new_n284), .A3(new_n576), .A4(new_n920), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n934), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n938), .A2(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT123), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(KEYINPUT60), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n947), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n922), .B2(new_n608), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT61), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n925), .A2(G190gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n681), .ZN(new_n953));
  NOR4_X1   g752(.A1(new_n925), .A2(KEYINPUT124), .A3(G190gat), .A4(new_n608), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1351gat));
  AND2_X1   g754(.A1(new_n508), .A2(new_n920), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n509), .B(new_n956), .C1(new_n877), .C2(new_n839), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n957), .A2(KEYINPUT125), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(G197gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n961), .A3(new_n741), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n921), .A2(new_n508), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n902), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n964), .A2(new_n263), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n965), .B2(new_n961), .ZN(G1352gat));
  NOR3_X1   g765(.A1(new_n957), .A2(G204gat), .A3(new_n646), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT62), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n902), .A2(new_n687), .A3(new_n963), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n635), .ZN(G1353gat));
  NAND4_X1  g769(.A1(new_n896), .A2(new_n576), .A3(new_n901), .A4(new_n963), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G211gat), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT63), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n973), .A2(KEYINPUT63), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(KEYINPUT63), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n971), .A2(G211gat), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(G211gat), .B1(new_n958), .B2(new_n959), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT126), .A3(new_n576), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT126), .B1(new_n978), .B2(new_n576), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n974), .B(new_n977), .C1(new_n979), .C2(new_n980), .ZN(G1354gat));
  AOI21_X1  g780(.A(G218gat), .B1(new_n960), .B2(new_n681), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n608), .A2(new_n360), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n964), .B2(new_n983), .ZN(G1355gat));
endmodule


