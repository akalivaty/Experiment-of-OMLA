//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT69), .A2(G237), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT69), .A2(G237), .ZN(new_n189));
  AOI21_X1  g003(.A(G953), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT27), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n191), .B(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(new_n193), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n187), .B1(new_n195), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n193), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n194), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT70), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n208), .A3(new_n212), .A4(new_n209), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(G131), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n210), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(G131), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G143), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  OR2_X1    g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT64), .B1(new_n221), .B2(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n219), .A3(G143), .ZN(new_n229));
  INV_X1    g043(.A(new_n224), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .A4(new_n222), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n218), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT2), .B(G113), .Z(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n236), .A2(new_n237), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT67), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(KEYINPUT1), .ZN(new_n249));
  AND4_X1   g063(.A1(new_n227), .A2(new_n229), .A3(new_n222), .A4(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n251), .A2(G128), .B1(new_n220), .B2(new_n222), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n205), .A2(G137), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n207), .A2(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(G131), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n216), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n210), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n251), .A2(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n223), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n227), .A2(new_n229), .A3(new_n222), .A4(new_n249), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n217), .A2(new_n263), .A3(new_n264), .A4(new_n256), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n233), .A2(new_n247), .A3(new_n259), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n247), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n226), .A2(new_n231), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n214), .B2(new_n217), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n253), .A2(new_n258), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n267), .B(new_n268), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n213), .A2(G131), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n274), .A2(new_n211), .B1(new_n216), .B2(new_n215), .ZN(new_n275));
  OAI22_X1  g089(.A1(new_n275), .A2(new_n269), .B1(new_n253), .B2(new_n258), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n268), .B1(new_n276), .B2(new_n267), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT28), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n276), .A2(new_n267), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n203), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n200), .A2(new_n201), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT30), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n233), .A2(new_n259), .A3(new_n265), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n284), .B1(KEYINPUT30), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n266), .B(new_n283), .C1(new_n286), .C2(new_n247), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n266), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n259), .A2(new_n265), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT30), .B1(new_n291), .B2(new_n270), .ZN(new_n292));
  OR3_X1    g106(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT30), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(new_n294), .B2(new_n267), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT31), .A3(new_n283), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n281), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT32), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n278), .A2(new_n280), .ZN(new_n301));
  INV_X1    g115(.A(new_n203), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT31), .B1(new_n295), .B2(new_n283), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n247), .B1(new_n292), .B2(new_n293), .ZN(new_n305));
  NOR4_X1   g119(.A1(new_n305), .A2(new_n288), .A3(new_n290), .A4(new_n282), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n298), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT72), .B1(new_n295), .B2(new_n283), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n278), .A2(new_n280), .A3(new_n203), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n314), .B(new_n282), .C1(new_n305), .C2(new_n290), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n285), .A2(new_n267), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n266), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n319), .B2(KEYINPUT28), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n282), .A2(new_n312), .ZN(new_n321));
  AOI21_X1  g135(.A(G902), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G472), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n310), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G234), .ZN(new_n326));
  OAI21_X1  g140(.A(G217), .B1(new_n326), .B2(G902), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n248), .A2(KEYINPUT23), .A3(G119), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT74), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n330));
  AOI22_X1  g144(.A1(KEYINPUT75), .A2(new_n330), .B1(new_n248), .B2(G119), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(KEYINPUT75), .B2(new_n330), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n238), .A2(G128), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n248), .A2(G119), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n333), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n337), .ZN(new_n340));
  INV_X1    g154(.A(new_n338), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT73), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n334), .A2(G110), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT16), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(G125), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n346), .B1(new_n350), .B2(new_n344), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT76), .A3(new_n219), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n219), .ZN(new_n353));
  OAI211_X1 g167(.A(G146), .B(new_n346), .C1(new_n350), .C2(new_n344), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n343), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n334), .A2(G110), .B1(new_n340), .B2(new_n341), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G125), .B(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT77), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n362), .A3(new_n219), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n363), .A3(new_n354), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT22), .B(G137), .ZN(new_n366));
  INV_X1    g180(.A(G221), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n367), .A2(new_n326), .A3(G953), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n366), .B(new_n368), .Z(new_n369));
  XNOR2_X1  g183(.A(new_n365), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT25), .ZN(new_n371));
  AOI21_X1  g185(.A(G902), .B1(new_n371), .B2(KEYINPUT78), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n371), .A2(KEYINPUT78), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n327), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n370), .B(new_n372), .C1(KEYINPUT78), .C2(new_n371), .ZN(new_n376));
  INV_X1    g190(.A(G902), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n327), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n375), .A2(new_n376), .B1(new_n370), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n325), .A2(KEYINPUT79), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n300), .A2(new_n309), .B1(new_n323), .B2(G472), .ZN(new_n383));
  INV_X1    g197(.A(new_n380), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(G107), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n392), .A2(KEYINPUT81), .A3(KEYINPUT3), .A4(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  OAI22_X1  g208(.A1(new_n392), .A2(G104), .B1(KEYINPUT81), .B2(KEYINPUT3), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n388), .B1(new_n397), .B2(G101), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  AND4_X1   g213(.A1(KEYINPUT82), .A2(new_n394), .A3(new_n399), .A4(new_n396), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n395), .B1(new_n391), .B2(new_n393), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT82), .B1(new_n401), .B2(new_n399), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n398), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n397), .A2(new_n388), .A3(G101), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n267), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n242), .A2(new_n243), .ZN(new_n406));
  INV_X1    g220(.A(G113), .ZN(new_n407));
  AND2_X1   g221(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n408));
  NOR2_X1   g222(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n239), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n235), .B1(new_n409), .B2(new_n408), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n392), .A2(G104), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n392), .A2(G104), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n399), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n414), .B(new_n419), .C1(new_n400), .C2(new_n402), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n387), .B1(new_n405), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT6), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT4), .B1(new_n401), .B2(new_n399), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n397), .B2(G101), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n401), .A2(KEYINPUT82), .A3(new_n399), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n404), .A2(new_n245), .A3(new_n246), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n420), .B(new_n387), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n405), .A2(KEYINPUT86), .A3(new_n420), .A4(new_n387), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n423), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n422), .B1(new_n434), .B2(new_n421), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n263), .A2(G125), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n348), .B1(new_n226), .B2(new_n231), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT87), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n437), .A2(KEYINPUT87), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G953), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G224), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n440), .B(new_n442), .Z(new_n443));
  NAND2_X1  g257(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT5), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(new_n242), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n235), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n448), .B(new_n449), .C1(new_n412), .C2(new_n450), .ZN(new_n451));
  AOI211_X1 g265(.A(KEYINPUT89), .B(new_n407), .C1(new_n410), .C2(new_n411), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n236), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n418), .B1(new_n426), .B2(new_n427), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n419), .B1(new_n400), .B2(new_n402), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n414), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n387), .B(KEYINPUT8), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n438), .A2(KEYINPUT7), .A3(new_n442), .A4(new_n439), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT7), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n442), .B1(new_n463), .B2(KEYINPUT7), .ZN(new_n464));
  OAI22_X1  g278(.A1(new_n436), .A2(new_n437), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n459), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n432), .A2(new_n433), .ZN(new_n467));
  AOI21_X1  g281(.A(G902), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI211_X1 g284(.A(KEYINPUT91), .B(G902), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n444), .B(new_n445), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n444), .B1(new_n470), .B2(new_n471), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT92), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n445), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n444), .B(KEYINPUT92), .C1(new_n470), .C2(new_n471), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT97), .ZN(new_n479));
  AOI21_X1  g293(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n480));
  AND2_X1   g294(.A1(KEYINPUT69), .A2(G237), .ZN(new_n481));
  NOR2_X1   g295(.A1(KEYINPUT69), .A2(G237), .ZN(new_n482));
  OAI211_X1 g296(.A(G214), .B(new_n441), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n221), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n257), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n221), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n216), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT96), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT96), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n485), .A2(new_n492), .A3(new_n486), .A4(new_n489), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n216), .B1(new_n487), .B2(new_n488), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n356), .A2(new_n352), .B1(new_n494), .B2(KEYINPUT17), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G113), .B(G122), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n390), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n350), .A2(G146), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n363), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT18), .ZN(new_n502));
  INV_X1    g316(.A(G131), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT93), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n487), .A2(new_n488), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n487), .B2(new_n488), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(KEYINPUT94), .A3(new_n501), .A4(new_n506), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n496), .A2(new_n498), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n485), .A2(new_n489), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT19), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n360), .A2(new_n362), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n350), .A2(KEYINPUT95), .A3(KEYINPUT19), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n361), .B2(new_n515), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n514), .B(new_n354), .C1(new_n520), .C2(G146), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n498), .B1(new_n512), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n479), .B1(new_n513), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(G475), .A2(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n512), .A2(new_n521), .ZN(new_n525));
  INV_X1    g339(.A(new_n498), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n496), .A2(new_n498), .A3(new_n512), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(KEYINPUT97), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n528), .ZN(new_n531));
  NOR3_X1   g345(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n530), .A2(KEYINPUT20), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G475), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n498), .B1(new_n496), .B2(new_n512), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n513), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n536), .B2(new_n377), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT9), .B(G234), .Z(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT80), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n367), .B1(new_n540), .B2(new_n377), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n227), .A2(new_n229), .A3(new_n222), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n260), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n262), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n419), .B(new_n544), .C1(new_n400), .C2(new_n402), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT10), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n403), .A2(new_n232), .A3(new_n404), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n253), .A2(new_n546), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n454), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n218), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n547), .A2(new_n548), .A3(new_n550), .A4(new_n275), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G140), .ZN(new_n555));
  INV_X1    g369(.A(G227), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G953), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n555), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n545), .B1(new_n454), .B2(new_n263), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n218), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT12), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(KEYINPUT12), .A3(new_n218), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n558), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n553), .A2(KEYINPUT83), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT83), .B1(new_n553), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n559), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n377), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n560), .A2(KEYINPUT12), .A3(new_n218), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT12), .B1(new_n560), .B2(new_n218), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n553), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n553), .A2(new_n566), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n575), .A2(new_n558), .B1(new_n576), .B2(new_n552), .ZN(new_n577));
  OAI21_X1  g391(.A(G469), .B1(new_n577), .B2(G902), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n541), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(G234), .A2(G237), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n580), .A2(G952), .A3(new_n441), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n580), .A2(G902), .A3(G953), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT21), .B(G898), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT15), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G478), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n221), .A2(G128), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n248), .A2(G143), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G134), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n588), .A3(new_n205), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G122), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G116), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n392), .B1(new_n596), .B2(KEYINPUT14), .ZN(new_n597));
  XNOR2_X1  g411(.A(G116), .B(G122), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n590), .A2(KEYINPUT98), .A3(new_n591), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n594), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT13), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n587), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n588), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n587), .A2(new_n602), .ZN(new_n605));
  OAI21_X1  g419(.A(G134), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n598), .A2(G107), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n598), .A2(G107), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n591), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n441), .A2(G217), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n540), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n601), .A2(new_n540), .A3(new_n611), .A4(new_n609), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(KEYINPUT99), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n610), .A2(new_n616), .A3(new_n612), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n377), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n586), .B1(new_n619), .B2(KEYINPUT100), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n615), .A2(KEYINPUT100), .A3(new_n377), .A4(new_n617), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n584), .B(new_n620), .C1(new_n624), .C2(new_n586), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n538), .A2(new_n579), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(G214), .B1(G237), .B2(G902), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT84), .Z(new_n628));
  NOR3_X1   g442(.A1(new_n478), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n386), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n399), .ZN(G3));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n432), .A2(new_n433), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n459), .A2(new_n460), .A3(new_n465), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n377), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT91), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n468), .A2(new_n469), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n636), .A2(new_n637), .B1(new_n443), .B2(new_n435), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n632), .B1(new_n638), .B2(new_n445), .ZN(new_n639));
  INV_X1    g453(.A(new_n445), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n474), .A2(KEYINPUT101), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n472), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n628), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n579), .A2(new_n380), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n297), .B2(G902), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n299), .B2(new_n297), .ZN(new_n647));
  INV_X1    g461(.A(new_n584), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n615), .A2(new_n649), .A3(new_n617), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n613), .A2(KEYINPUT33), .A3(new_n614), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(G478), .A3(new_n377), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n619), .A2(G478), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n648), .B(new_n655), .C1(new_n533), .C2(new_n537), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n645), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n644), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  NOR2_X1   g474(.A1(new_n645), .A2(new_n647), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n530), .A2(KEYINPUT20), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT20), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n523), .A2(new_n529), .A3(new_n663), .A4(new_n524), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n537), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n620), .B1(new_n624), .B2(new_n586), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n667), .A2(new_n584), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n644), .A2(new_n661), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NAND2_X1  g486(.A1(new_n375), .A2(new_n376), .ZN(new_n673));
  INV_X1    g487(.A(new_n369), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n365), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n379), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n647), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n629), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  INV_X1    g495(.A(new_n668), .ZN(new_n682));
  INV_X1    g496(.A(new_n581), .ZN(new_n683));
  INV_X1    g497(.A(new_n582), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n683), .B1(new_n684), .B2(G900), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n666), .A2(new_n682), .A3(new_n665), .A4(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n642), .A3(new_n643), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n673), .A2(new_n677), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n325), .A2(new_n579), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n248), .ZN(G30));
  XNOR2_X1  g505(.A(new_n478), .B(KEYINPUT38), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n538), .A2(new_n668), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n295), .A2(new_n283), .B1(new_n302), .B2(new_n319), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n310), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n628), .A3(new_n688), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n685), .B(KEYINPUT39), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n579), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  NAND4_X1  g516(.A1(new_n693), .A2(new_n694), .A3(new_n699), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  INV_X1    g518(.A(new_n689), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n531), .A2(new_n532), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n662), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n666), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n655), .A3(new_n685), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n705), .A2(new_n644), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NOR2_X1   g526(.A1(new_n383), .A2(new_n384), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n707), .A2(new_n666), .B1(new_n654), .B2(new_n653), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n648), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n553), .A2(new_n566), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT83), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n565), .A3(new_n567), .ZN(new_n719));
  AOI21_X1  g533(.A(G902), .B1(new_n719), .B2(new_n559), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n541), .B1(new_n720), .B2(new_n571), .ZN(new_n721));
  OAI21_X1  g535(.A(G469), .B1(new_n720), .B2(KEYINPUT102), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n570), .A2(KEYINPUT102), .A3(new_n377), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT103), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n726), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n725), .A2(new_n642), .A3(new_n643), .A4(new_n727), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n715), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT104), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT41), .B(G113), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND4_X1  g546(.A1(new_n713), .A2(new_n669), .A3(new_n643), .A4(new_n642), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n725), .A2(new_n727), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  AND2_X1   g550(.A1(new_n538), .A2(new_n625), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n325), .A3(new_n688), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n728), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n238), .ZN(G21));
  OAI22_X1  g554(.A1(new_n304), .A2(new_n306), .B1(new_n203), .B2(new_n320), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n298), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n648), .A2(new_n380), .A3(new_n646), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n725), .A2(new_n743), .A3(new_n727), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n642), .A2(new_n694), .A3(new_n643), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n595), .ZN(G24));
  AND2_X1   g561(.A1(new_n646), .A2(new_n742), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n688), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n710), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n728), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n348), .ZN(G27));
  NAND2_X1  g566(.A1(new_n472), .A2(new_n643), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n476), .B2(new_n477), .ZN(new_n754));
  NAND2_X1  g568(.A1(G469), .A2(G902), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT105), .Z(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n577), .B2(G469), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n541), .B1(new_n572), .B2(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n754), .A2(KEYINPUT106), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT106), .B1(new_n754), .B2(new_n759), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n713), .B(new_n710), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n754), .A2(new_n759), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n754), .A2(KEYINPUT106), .A3(new_n759), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(KEYINPUT42), .A3(new_n713), .A4(new_n710), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  OAI211_X1 g586(.A(new_n713), .B(new_n686), .C1(new_n760), .C2(new_n761), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n769), .A2(KEYINPUT107), .A3(new_n713), .A4(new_n686), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n538), .A2(new_n655), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT43), .Z(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n647), .A3(new_n688), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n577), .A2(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n577), .A2(KEYINPUT45), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(G469), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n756), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n572), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n541), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n792), .A2(new_n700), .A3(new_n754), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n781), .A2(new_n782), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n783), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(KEYINPUT47), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n799));
  MUX2_X1   g613(.A(new_n798), .B(new_n799), .S(new_n792), .Z(new_n800));
  INV_X1    g614(.A(new_n754), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(new_n325), .A3(new_n380), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n710), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NOR4_X1   g618(.A1(new_n779), .A2(new_n628), .A3(new_n541), .A4(new_n384), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n722), .A2(new_n723), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n571), .B2(new_n720), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT109), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n697), .B1(new_n808), .B2(new_n806), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n692), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n640), .B1(new_n638), .B2(KEYINPUT92), .ZN(new_n814));
  INV_X1    g628(.A(new_n477), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n472), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n533), .A2(new_n668), .A3(new_n537), .A4(new_n584), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n643), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT111), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n816), .A2(new_n820), .A3(new_n643), .A4(new_n817), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n661), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n478), .A2(new_n628), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n386), .A2(new_n629), .B1(new_n823), .B2(new_n657), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n822), .B(new_n679), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI221_X4 g640(.A(KEYINPUT110), .B1(new_n823), .B2(new_n657), .C1(new_n386), .C2(new_n629), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n813), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n823), .A2(new_n657), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT110), .B1(new_n630), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n661), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n818), .B2(KEYINPUT111), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n832), .A2(new_n821), .B1(new_n629), .B2(new_n678), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n824), .A2(new_n825), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n830), .A2(new_n833), .A3(KEYINPUT112), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n728), .A2(new_n738), .B1(new_n744), .B2(new_n745), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT114), .A3(new_n735), .A4(new_n729), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  OAI22_X1  g654(.A1(new_n733), .A2(new_n734), .B1(new_n715), .B2(new_n728), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(new_n837), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n728), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n714), .A2(new_n748), .A3(new_n688), .A4(new_n685), .ZN(new_n845));
  INV_X1    g659(.A(new_n687), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n844), .A2(new_n845), .B1(new_n846), .B2(new_n705), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n642), .A2(new_n714), .A3(new_n643), .A4(new_n685), .ZN(new_n848));
  INV_X1    g662(.A(new_n685), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n688), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n697), .A2(new_n759), .A3(new_n850), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n848), .A2(new_n689), .B1(new_n745), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n853), .A3(KEYINPUT52), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n750), .A2(new_n728), .B1(new_n687), .B2(new_n689), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n856), .B2(new_n852), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n845), .B1(new_n760), .B2(new_n761), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n667), .A2(new_n682), .A3(new_n849), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n705), .A2(new_n754), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n775), .B2(new_n776), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n764), .B2(new_n770), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n843), .A2(new_n858), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT115), .B1(new_n836), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n828), .A2(new_n835), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n863), .A2(new_n865), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n839), .A2(new_n842), .B1(new_n854), .B2(new_n857), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT113), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT52), .B1(new_n847), .B2(new_n853), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n856), .A2(new_n852), .A3(new_n855), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n854), .A2(KEYINPUT113), .A3(new_n857), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n863), .A2(new_n771), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n841), .A2(new_n837), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(new_n868), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n864), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n873), .A2(new_n874), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(KEYINPUT53), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT53), .B1(new_n854), .B2(new_n857), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n868), .A2(new_n881), .A3(new_n882), .A4(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(KEYINPUT54), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n885), .A2(KEYINPUT116), .A3(new_n889), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n748), .A2(new_n581), .A3(new_n380), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n780), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n808), .A2(new_n541), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n754), .B(new_n897), .C1(new_n800), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n734), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT118), .B1(new_n901), .B2(new_n754), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n734), .A2(new_n903), .A3(new_n801), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n904), .A3(new_n683), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n749), .A3(new_n780), .ZN(new_n906));
  NOR4_X1   g720(.A1(new_n896), .A2(new_n693), .A3(new_n643), .A4(new_n734), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT50), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n900), .A2(new_n906), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n905), .A2(new_n380), .A3(new_n698), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n912), .A2(new_n708), .A3(new_n655), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n894), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT51), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n894), .B(new_n916), .C1(new_n911), .C2(new_n913), .ZN(new_n917));
  INV_X1    g731(.A(G952), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n918), .B(G953), .C1(new_n897), .C2(new_n844), .ZN(new_n919));
  INV_X1    g733(.A(new_n714), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n905), .A2(new_n713), .A3(new_n780), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(KEYINPUT48), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(KEYINPUT48), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n915), .A2(new_n917), .A3(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n892), .A2(new_n893), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(G952), .A2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n812), .B1(new_n927), .B2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n441), .A2(G952), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT119), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI22_X1  g746(.A1(new_n867), .A2(new_n872), .B1(new_n883), .B2(new_n864), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n377), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT56), .B1(new_n934), .B2(G210), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n435), .B(new_n443), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n937), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(G51));
  AOI21_X1  g754(.A(KEYINPUT120), .B1(new_n933), .B2(new_n874), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n873), .A2(new_n884), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT54), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n756), .B(KEYINPUT57), .Z(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n570), .B(KEYINPUT121), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n786), .B(KEYINPUT122), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n934), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n930), .B1(new_n949), .B2(new_n951), .ZN(G54));
  NAND3_X1  g766(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n523), .A2(new_n529), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n930), .ZN(G60));
  NAND2_X1  g771(.A1(new_n892), .A2(new_n893), .ZN(new_n958));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n652), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n652), .A2(new_n961), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n944), .A2(new_n945), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n931), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n962), .A2(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT123), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT60), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n942), .A2(new_n676), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n931), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n942), .A2(new_n970), .ZN(new_n975));
  INV_X1    g789(.A(new_n370), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n967), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  AND4_X1   g792(.A1(new_n967), .A2(new_n977), .A3(new_n971), .A4(new_n973), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G66));
  NAND2_X1  g794(.A1(new_n868), .A2(new_n882), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n441), .ZN(new_n982));
  INV_X1    g796(.A(G224), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n583), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(KEYINPUT125), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(KEYINPUT125), .B2(new_n982), .ZN(new_n986));
  INV_X1    g800(.A(new_n435), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(G898), .B2(new_n441), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n986), .B(new_n988), .Z(G69));
  NOR2_X1   g803(.A1(new_n801), .A2(new_n701), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n920), .B1(new_n708), .B2(new_n668), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n386), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n803), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n847), .A2(new_n711), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n703), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n993), .A2(new_n795), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n441), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n294), .B(new_n520), .ZN(new_n1000));
  INV_X1    g814(.A(new_n745), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n792), .A2(new_n713), .A3(new_n700), .A4(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n803), .A2(new_n795), .A3(new_n994), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n771), .A2(new_n777), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n441), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1000), .B1(G900), .B2(G953), .ZN(new_n1007));
  AOI22_X1  g821(.A1(new_n999), .A2(new_n1000), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n441), .B1(G227), .B2(G900), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(G72));
  NAND3_X1  g824(.A1(new_n1005), .A2(new_n868), .A3(new_n882), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n305), .A2(new_n290), .A3(new_n283), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n930), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n311), .A2(new_n315), .ZN(new_n1017));
  AOI22_X1  g831(.A1(new_n1017), .A2(KEYINPUT126), .B1(new_n283), .B2(new_n295), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(KEYINPUT126), .B2(new_n1017), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n1013), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT127), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n886), .A2(new_n888), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1013), .B1(new_n998), .B2(new_n981), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1023), .B(new_n283), .C1(new_n290), .C2(new_n305), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1016), .A2(new_n1022), .A3(new_n1024), .ZN(G57));
endmodule


