//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT67), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT70), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(new_n462), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n464), .A2(G137), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n460), .A2(new_n463), .B1(KEYINPUT3), .B2(new_n459), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(KEYINPUT71), .A3(G137), .A4(new_n465), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n459), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n469), .A2(new_n471), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(KEYINPUT69), .B1(new_n475), .B2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n462), .A2(G2104), .ZN(new_n477));
  AND4_X1   g052(.A1(KEYINPUT69), .A2(new_n466), .A3(new_n477), .A4(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND3_X1  g057(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n464), .A2(G2105), .A3(new_n466), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(G124), .B2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT72), .Z(G162));
  NAND4_X1  g066(.A1(new_n464), .A2(G126), .A3(G2105), .A4(new_n466), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n493));
  OR3_X1    g068(.A1(new_n465), .A2(KEYINPUT73), .A3(G114), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT73), .B1(new_n465), .B2(G114), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n494), .A2(G2104), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n492), .B2(new_n497), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT4), .A2(G138), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n466), .A2(new_n477), .A3(G138), .A4(new_n465), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n498), .A2(new_n499), .A3(new_n505), .ZN(G164));
  NAND2_X1  g081(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n510), .ZN(new_n515));
  AOI21_X1  g090(.A(G543), .B1(KEYINPUT75), .B2(KEYINPUT5), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI21_X1  g096(.A(G543), .B1(new_n517), .B2(new_n518), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n514), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI221_X1 g103(.A(new_n526), .B1(new_n527), .B2(new_n522), .C1(new_n519), .C2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  OR3_X1    g105(.A1(new_n515), .A2(KEYINPUT76), .A3(new_n516), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n511), .A2(KEYINPUT76), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n533), .A2(G63), .A3(G651), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  INV_X1    g110(.A(new_n519), .ZN(new_n536));
  INV_X1    g111(.A(new_n522), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n536), .A2(G90), .B1(G52), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n533), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n513), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n533), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n513), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n519), .A2(new_n544), .B1(new_n545), .B2(new_n522), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT77), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n537), .A2(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n536), .A2(G91), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n513), .C2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G168), .ZN(G286));
  INV_X1    g135(.A(G166), .ZN(G303));
  OAI21_X1  g136(.A(G651), .B1(new_n533), .B2(G74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n536), .A2(G87), .B1(G49), .B2(new_n537), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(G288));
  OAI21_X1  g139(.A(G61), .B1(new_n515), .B2(new_n516), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT78), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n511), .A2(new_n568), .A3(G61), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  INV_X1    g147(.A(G48), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n519), .A2(new_n572), .B1(new_n573), .B2(new_n522), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G305));
  XNOR2_X1  g151(.A(KEYINPUT79), .B(G85), .ZN(new_n577));
  INV_X1    g152(.A(G47), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n519), .A2(new_n577), .B1(new_n578), .B2(new_n522), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n533), .A2(G60), .ZN(new_n580));
  INV_X1    g155(.A(G72), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n508), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n579), .B1(new_n582), .B2(G651), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT80), .Z(new_n586));
  NAND2_X1  g161(.A1(new_n536), .A2(G92), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n511), .A2(G66), .ZN(new_n590));
  INV_X1    g165(.A(G79), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n508), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n537), .B2(G54), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT81), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n586), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n586), .B1(new_n596), .B2(G868), .ZN(G321));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  XNOR2_X1  g174(.A(G299), .B(KEYINPUT82), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G297));
  XOR2_X1   g176(.A(G297), .B(KEYINPUT83), .Z(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  OR2_X1    g179(.A1(new_n543), .A2(new_n546), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n595), .A2(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n475), .A2(new_n472), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n489), .A2(G123), .ZN(new_n615));
  INV_X1    g190(.A(new_n483), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G135), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n465), .A2(G111), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT84), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n615), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n614), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2435), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2438), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(G14), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2072), .B(G2078), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(KEYINPUT85), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT17), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n639), .B2(new_n641), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n640), .A2(new_n641), .ZN(new_n647));
  MUX2_X1   g222(.A(new_n647), .B(new_n641), .S(new_n639), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n643), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2100), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n655), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n659), .A3(new_n661), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n665), .C1(new_n663), .C2(new_n662), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(G1986), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1991), .B(G1996), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT22), .B(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G29), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G27), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G164), .B2(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(G2078), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT30), .B(G28), .ZN(new_n679));
  OR2_X1    g254(.A1(KEYINPUT31), .A2(G11), .ZN(new_n680));
  NAND2_X1  g255(.A1(KEYINPUT31), .A2(G11), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n679), .A2(new_n674), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n621), .B2(new_n674), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT97), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(KEYINPUT97), .ZN(new_n685));
  NOR2_X1   g260(.A1(G5), .A2(G16), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G171), .B2(G16), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n684), .A2(new_n685), .B1(new_n687), .B2(G1961), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT96), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G168), .B2(G16), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G16), .B2(G21), .ZN(new_n691));
  NAND3_X1  g266(.A1(G168), .A2(new_n689), .A3(G16), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n691), .A2(G1966), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(G1966), .B1(new_n691), .B2(new_n692), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n688), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(KEYINPUT98), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT98), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(new_n688), .C1(new_n693), .C2(new_n694), .ZN(new_n698));
  INV_X1    g273(.A(G1956), .ZN(new_n699));
  NAND2_X1  g274(.A1(G299), .A2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n701), .A2(KEYINPUT23), .A3(G20), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n703));
  INV_X1    g278(.A(G20), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G16), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT100), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n696), .A2(new_n698), .B1(new_n699), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(G6), .A2(G16), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G305), .B2(new_n701), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT32), .B(G1981), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n715), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n713), .B(new_n717), .C1(G305), .C2(new_n701), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n562), .A2(G16), .A3(new_n563), .ZN(new_n720));
  OR2_X1    g295(.A1(G16), .A2(G23), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT33), .B(G1976), .Z(new_n722));
  AND3_X1   g297(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n720), .B2(new_n721), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(G16), .B1(new_n514), .B2(new_n523), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n701), .A2(G22), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G1971), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n726), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT34), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n719), .A2(new_n725), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(G95), .A2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n736), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n737));
  INV_X1    g312(.A(G131), .ZN(new_n738));
  INV_X1    g313(.A(G119), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n737), .B1(new_n483), .B2(new_n738), .C1(new_n739), .C2(new_n488), .ZN(new_n740));
  MUX2_X1   g315(.A(G25), .B(new_n740), .S(G29), .Z(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT35), .B(G1991), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n741), .B(new_n742), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n701), .A2(G24), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n583), .B2(new_n701), .ZN(new_n745));
  INV_X1    g320(.A(G1986), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(G1986), .B(new_n744), .C1(new_n583), .C2(new_n701), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n735), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n735), .A2(new_n743), .A3(new_n749), .A4(KEYINPUT87), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n732), .A2(new_n723), .A3(new_n724), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n734), .B1(new_n755), .B2(new_n719), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n712), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n756), .B(new_n711), .C1(new_n752), .C2(new_n753), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n678), .B(new_n708), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT99), .A2(G2084), .ZN(new_n761));
  OR2_X1    g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT24), .A2(G34), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n762), .A2(new_n674), .A3(new_n763), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n761), .B(new_n764), .C1(G160), .C2(new_n674), .ZN(new_n765));
  NOR2_X1   g340(.A1(KEYINPUT99), .A2(G2084), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G29), .A2(G35), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G162), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT29), .Z(new_n771));
  INV_X1    g346(.A(G2090), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n771), .A2(new_n772), .B1(new_n699), .B2(new_n707), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n760), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n547), .A2(new_n701), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n701), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT90), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(KEYINPUT90), .B2(new_n776), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G1341), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n771), .A2(new_n772), .ZN(new_n780));
  OR2_X1    g355(.A1(G29), .A2(G32), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n616), .A2(G141), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n489), .A2(G129), .B1(G105), .B2(new_n472), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT95), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT26), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n783), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n781), .B1(new_n788), .B2(new_n674), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT27), .B(G1996), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n674), .A2(G26), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(G128), .A2(new_n489), .B1(new_n616), .B2(G140), .ZN(new_n795));
  OR3_X1    g370(.A1(KEYINPUT91), .A2(G104), .A3(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G116), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n459), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT91), .B1(G104), .B2(G2105), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT92), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n794), .B1(new_n802), .B2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2067), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n687), .A2(G1961), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n789), .A2(new_n790), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n791), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n774), .A2(new_n779), .A3(new_n780), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n596), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G4), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT89), .B(G1348), .Z(new_n812));
  XOR2_X1   g387(.A(new_n811), .B(new_n812), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n616), .A2(G139), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n472), .A2(G103), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT25), .Z(new_n816));
  AOI22_X1  g391(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n814), .B(new_n816), .C1(new_n465), .C2(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G33), .B(new_n818), .S(G29), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2072), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n809), .A2(new_n813), .A3(new_n820), .ZN(G311));
  AOI21_X1  g396(.A(new_n756), .B1(new_n752), .B2(new_n753), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n712), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n823), .A2(new_n678), .A3(new_n708), .A4(new_n767), .ZN(new_n824));
  INV_X1    g399(.A(new_n780), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n824), .A2(new_n825), .A3(new_n807), .A4(new_n773), .ZN(new_n826));
  INV_X1    g401(.A(new_n813), .ZN(new_n827));
  INV_X1    g402(.A(new_n820), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n826), .A2(new_n827), .A3(new_n779), .A4(new_n828), .ZN(G150));
  AOI22_X1  g404(.A1(new_n533), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n513), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n519), .A2(new_n832), .B1(new_n833), .B2(new_n522), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT101), .Z(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n547), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n605), .A2(new_n835), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n595), .A2(new_n603), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n839), .B1(new_n846), .B2(G860), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT102), .ZN(G145));
  XNOR2_X1  g423(.A(new_n481), .B(new_n621), .ZN(new_n849));
  XNOR2_X1  g424(.A(G162), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n788), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n818), .B(new_n612), .Z(new_n852));
  NAND4_X1  g427(.A1(new_n501), .A2(new_n492), .A3(new_n504), .A4(new_n497), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n802), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(G142), .ZN(new_n856));
  NOR2_X1   g431(.A1(G106), .A2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n483), .A2(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G130), .B2(new_n489), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n740), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n855), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n851), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g441(.A(new_n608), .B(new_n842), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n594), .B(G299), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT103), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n868), .B(KEYINPUT41), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT42), .ZN(new_n876));
  XNOR2_X1  g451(.A(G303), .B(G288), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G305), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G290), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n870), .A2(new_n872), .A3(new_n880), .A4(new_n874), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n876), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n879), .B1(new_n876), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(G868), .B2(new_n835), .ZN(G295));
  OAI21_X1  g460(.A(new_n884), .B1(G868), .B2(new_n835), .ZN(G331));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  XNOR2_X1  g462(.A(G168), .B(G301), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n842), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n842), .B(new_n888), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(new_n887), .ZN(new_n891));
  INV_X1    g466(.A(new_n871), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n891), .A2(new_n868), .B1(new_n892), .B2(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n879), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n864), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n891), .A2(new_n871), .ZN(new_n896));
  INV_X1    g471(.A(new_n868), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n879), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n895), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n893), .A2(new_n879), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n893), .B2(new_n879), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT43), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT44), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n895), .A2(new_n899), .A3(KEYINPUT43), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n905), .B1(new_n908), .B2(KEYINPUT44), .ZN(G397));
  NAND3_X1  g484(.A1(new_n473), .A2(G40), .A3(new_n480), .ZN(new_n910));
  INV_X1    g485(.A(G1384), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n853), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G1996), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n788), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n802), .A2(G2067), .ZN(new_n918));
  INV_X1    g493(.A(G2067), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n795), .A2(new_n919), .A3(new_n801), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n742), .B2(new_n740), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n740), .A2(new_n742), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G290), .A2(G1986), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT106), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n583), .A2(new_n746), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT105), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n915), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G8), .ZN(new_n932));
  NOR2_X1   g507(.A1(G168), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n492), .A2(new_n497), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT74), .ZN(new_n935));
  INV_X1    g510(.A(new_n505), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(KEYINPUT45), .A3(new_n911), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n473), .A2(G40), .A3(new_n480), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n940), .A3(new_n914), .ZN(new_n941));
  INV_X1    g516(.A(G1966), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n944));
  XOR2_X1   g519(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n945));
  NOR2_X1   g520(.A1(new_n912), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT117), .B(G2084), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n944), .A2(new_n940), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n943), .A2(KEYINPUT121), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT121), .B1(new_n943), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n933), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n953));
  OAI21_X1  g528(.A(G8), .B1(new_n950), .B2(new_n951), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n933), .B(KEYINPUT122), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n943), .A2(new_n949), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(G8), .A3(G168), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n953), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(new_n933), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n952), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n963));
  NAND4_X1  g538(.A1(G303), .A2(KEYINPUT111), .A3(new_n963), .A4(G8), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(G166), .B2(new_n932), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n853), .A2(KEYINPUT45), .A3(new_n911), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n853), .A2(KEYINPUT108), .A3(KEYINPUT45), .A4(new_n911), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT45), .B1(new_n938), .B2(new_n911), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n974), .B(new_n913), .C1(G164), .C2(G1384), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n940), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT109), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n910), .B1(new_n973), .B2(new_n974), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n913), .B1(G164), .B2(G1384), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT107), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n979), .A2(new_n981), .A3(new_n982), .A4(new_n972), .ZN(new_n983));
  AOI21_X1  g558(.A(G1971), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n944), .A2(new_n940), .A3(new_n947), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(G2090), .ZN(new_n986));
  OAI211_X1 g561(.A(G8), .B(new_n967), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n562), .A2(new_n563), .A3(new_n989), .A4(G1976), .ZN(new_n990));
  OAI211_X1 g565(.A(G8), .B(new_n990), .C1(new_n910), .C2(new_n912), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G288), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n989), .B1(new_n993), .B2(G1976), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n988), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n988), .B1(new_n993), .B2(G1976), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n991), .A2(new_n997), .A3(new_n994), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n571), .B2(new_n575), .ZN(new_n1001));
  AOI211_X1 g576(.A(G1981), .B(new_n574), .C1(new_n570), .C2(G651), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT49), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n910), .A2(new_n912), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(new_n932), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n999), .B(new_n1007), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1004), .A2(new_n1006), .A3(KEYINPUT114), .A4(new_n1008), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n996), .B(new_n998), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n987), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n983), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n980), .A2(KEYINPUT107), .B1(new_n970), .B2(new_n971), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n982), .B1(new_n1016), .B2(new_n979), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n730), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n938), .A2(new_n1020), .A3(new_n911), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n912), .A2(new_n945), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n940), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(G2090), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1019), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT116), .B1(new_n984), .B2(new_n1024), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  INV_X1    g603(.A(new_n967), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1014), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1020), .B1(new_n938), .B2(new_n911), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1031), .A2(new_n910), .A3(new_n946), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G1961), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n978), .A2(new_n677), .A3(new_n983), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n941), .A2(new_n1035), .A3(G2078), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G301), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT62), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n952), .B(new_n1040), .C1(new_n956), .C2(new_n960), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n962), .A2(new_n1030), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n986), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n932), .B1(new_n1018), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(new_n967), .A3(new_n1013), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1006), .B(KEYINPUT115), .ZN(new_n1046));
  AOI211_X1 g621(.A(G1976), .B(G288), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n1002), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n473), .B(KEYINPUT123), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n479), .B(KEYINPUT124), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1051), .B(G40), .C1(new_n465), .C2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n972), .A2(KEYINPUT53), .A3(new_n677), .A4(new_n914), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1033), .B(new_n1055), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT125), .B1(new_n1056), .B2(G301), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1037), .B(new_n1033), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(G301), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1055), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1036), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT125), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(G171), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1057), .A2(new_n1060), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1030), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1036), .A2(G301), .A3(new_n1061), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1058), .B1(new_n1067), .B2(new_n1039), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1023), .A2(new_n699), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n979), .A2(new_n981), .A3(new_n972), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT56), .B(G2072), .Z(new_n1071));
  OAI21_X1  g646(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(G299), .B(KEYINPUT57), .Z(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1073), .B(new_n1069), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1076));
  INV_X1    g651(.A(new_n594), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1005), .A2(new_n1078), .A3(new_n919), .ZN(new_n1079));
  INV_X1    g654(.A(new_n912), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1080), .A2(G40), .A3(new_n480), .A4(new_n473), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT120), .B1(new_n1081), .B2(G2067), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1079), .B(new_n1082), .C1(new_n1032), .C2(G1348), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1076), .A2(new_n1077), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT58), .B(G1341), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1005), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n975), .A2(new_n977), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n916), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1089), .B2(new_n605), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1083), .A2(new_n594), .ZN(new_n1091));
  INV_X1    g666(.A(G1348), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n985), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(new_n1077), .A3(new_n1079), .A4(new_n1082), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(KEYINPUT60), .A3(new_n1094), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1070), .A2(G1996), .B1(new_n1005), .B2(new_n1086), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(KEYINPUT59), .A3(new_n547), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1078), .B1(new_n1005), .B2(new_n919), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1092), .B2(new_n985), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1090), .A2(new_n1095), .A3(new_n1097), .A4(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1076), .B(KEYINPUT61), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1075), .B(new_n1084), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1068), .A2(new_n1104), .A3(new_n961), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1042), .B(new_n1050), .C1(new_n1066), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1014), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n1109));
  OAI21_X1  g684(.A(G8), .B1(new_n984), .B2(new_n986), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n1029), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n958), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n957), .A2(KEYINPUT118), .A3(G8), .A4(G168), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1107), .A2(new_n1108), .A3(new_n1111), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT63), .B1(new_n1044), .B2(new_n967), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n987), .A2(new_n1013), .A3(new_n1115), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT119), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT63), .B1(new_n1030), .B2(new_n1115), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n931), .B1(new_n1106), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1124), .A2(new_n915), .ZN(new_n1125));
  INV_X1    g700(.A(new_n921), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n915), .B1(new_n1126), .B2(new_n788), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT46), .ZN(new_n1128));
  INV_X1    g703(.A(new_n915), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(G1996), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n915), .A2(KEYINPUT46), .A3(new_n916), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT47), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n925), .A2(new_n915), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n929), .A2(new_n1129), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT48), .Z(new_n1136));
  AOI211_X1 g711(.A(new_n1125), .B(new_n1133), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1123), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g713(.A1(new_n637), .A2(G319), .A3(new_n652), .ZN(new_n1140));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n1141));
  XNOR2_X1  g715(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  NAND2_X1  g716(.A1(new_n1142), .A2(new_n865), .ZN(new_n1143));
  NOR3_X1   g717(.A1(new_n908), .A2(G229), .A3(new_n1143), .ZN(G308));
  AND2_X1   g718(.A1(new_n1142), .A2(new_n865), .ZN(new_n1145));
  INV_X1    g719(.A(G229), .ZN(new_n1146));
  OAI211_X1 g720(.A(new_n1145), .B(new_n1146), .C1(new_n906), .C2(new_n907), .ZN(G225));
endmodule


