//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT2), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT81), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(new_n204), .B2(new_n205), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n206), .A2(new_n209), .B1(new_n204), .B2(new_n205), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  XNOR2_X1  g014(.A(G197gat), .B(G204gat), .ZN(new_n216));
  INV_X1    g015(.A(G211gat), .ZN(new_n217));
  INV_X1    g016(.A(G218gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(KEYINPUT22), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G211gat), .B(G218gat), .Z(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n214), .B1(new_n215), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n211), .A2(new_n215), .A3(new_n212), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n226), .B2(new_n223), .ZN(new_n227));
  INV_X1    g026(.A(G228gat), .ZN(new_n228));
  INV_X1    g027(.A(G233gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n225), .A2(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n215), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n213), .ZN(new_n232));
  INV_X1    g031(.A(new_n227), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n228), .A2(new_n229), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G22gat), .ZN(new_n237));
  INV_X1    g036(.A(G22gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(new_n230), .B2(new_n235), .ZN(new_n239));
  XOR2_X1   g038(.A(G78gat), .B(G106gat), .Z(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT31), .B(G50gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n237), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n236), .A2(G22gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT84), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(KEYINPUT84), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT83), .B1(new_n236), .B2(G22gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT83), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n230), .A2(new_n235), .A3(new_n249), .A4(new_n238), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n246), .A2(new_n247), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n243), .B1(new_n251), .B2(new_n242), .ZN(new_n252));
  NAND2_X1  g051(.A1(G226gat), .A2(G233gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT23), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(KEYINPUT65), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(new_n254), .B2(KEYINPUT23), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n257), .A2(new_n259), .B1(KEYINPUT23), .B2(new_n254), .ZN(new_n260));
  NAND3_X1  g059(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(G183gat), .B2(G190gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G169gat), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n274), .A2(new_n261), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT25), .B1(new_n267), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n278), .B2(new_n267), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n280), .A3(new_n260), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n271), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT28), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n267), .B1(KEYINPUT26), .B2(new_n255), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n255), .A2(KEYINPUT26), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n288), .A2(new_n289), .B1(G183gat), .B2(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n253), .B1(new_n292), .B2(KEYINPUT29), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT77), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n287), .A2(KEYINPUT69), .A3(new_n290), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n282), .ZN(new_n299));
  INV_X1    g098(.A(new_n253), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n253), .C1(new_n292), .C2(KEYINPUT29), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n294), .A2(new_n301), .A3(new_n222), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n296), .A2(new_n297), .ZN(new_n305));
  INV_X1    g104(.A(new_n282), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n223), .B(new_n253), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n222), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n300), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G8gat), .B(G36gat), .Z(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT78), .ZN(new_n312));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n312), .B(new_n313), .Z(new_n314));
  NAND4_X1  g113(.A1(new_n304), .A2(KEYINPUT30), .A3(new_n310), .A4(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT79), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n304), .A2(new_n310), .A3(new_n314), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n304), .B2(new_n310), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G127gat), .B(G134gat), .Z(new_n325));
  XOR2_X1   g124(.A(KEYINPUT70), .B(G120gat), .Z(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G113gat), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT71), .B(G113gat), .Z(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G120gat), .ZN(new_n329));
  AOI211_X1 g128(.A(KEYINPUT1), .B(new_n325), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(G113gat), .A2(G120gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(G113gat), .A2(G120gat), .ZN(new_n332));
  OR3_X1    g131(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT1), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n333), .A2(new_n325), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n214), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n330), .A2(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n226), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n335), .A2(new_n214), .A3(KEYINPUT4), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n338), .A2(new_n341), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n213), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n347), .B2(new_n336), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n344), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT0), .ZN(new_n352));
  XNOR2_X1  g151(.A(G57gat), .B(G85gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT6), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n346), .A2(new_n354), .A3(new_n349), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(KEYINPUT82), .A3(new_n357), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n252), .B1(new_n324), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n354), .B(KEYINPUT85), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n346), .A2(KEYINPUT86), .A3(new_n349), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT86), .B1(new_n346), .B2(new_n349), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n363), .B1(new_n370), .B2(new_n356), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT37), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n314), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n320), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n304), .B2(new_n310), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT38), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n307), .A2(new_n309), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n372), .B1(new_n377), .B2(new_n222), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n294), .A2(new_n301), .A3(new_n308), .A4(new_n303), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT38), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n320), .B2(new_n373), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n371), .A2(new_n376), .A3(new_n381), .A4(new_n317), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n251), .A2(new_n242), .ZN(new_n383));
  INV_X1    g182(.A(new_n243), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n367), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n338), .A2(new_n341), .A3(new_n343), .ZN(new_n387));
  INV_X1    g186(.A(new_n342), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n389), .B2(KEYINPUT39), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n347), .A2(new_n342), .A3(new_n336), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT39), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n392), .B1(new_n387), .B2(new_n388), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT40), .ZN(new_n394));
  OR3_X1    g193(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n390), .B2(new_n393), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n370), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n382), .B(new_n385), .C1(new_n323), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT36), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n335), .A2(KEYINPUT72), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT72), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n330), .B2(new_n334), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n305), .B2(new_n306), .ZN(new_n404));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n298), .A2(new_n282), .A3(new_n402), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT74), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n408), .A2(KEYINPUT34), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(KEYINPUT34), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n410), .B(KEYINPUT75), .Z(new_n411));
  AND3_X1   g210(.A1(new_n407), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n407), .B2(new_n409), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n405), .B1(new_n404), .B2(new_n406), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT73), .B(KEYINPUT33), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n417), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT32), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n406), .ZN(new_n425));
  INV_X1    g224(.A(new_n405), .ZN(new_n426));
  AOI221_X4 g225(.A(new_n422), .B1(new_n420), .B2(new_n417), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n414), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n409), .ZN(new_n429));
  INV_X1    g228(.A(new_n411), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n409), .A3(new_n411), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n298), .A2(new_n282), .B1(new_n400), .B2(new_n402), .ZN(new_n434));
  AND4_X1   g233(.A1(new_n282), .A2(new_n402), .A3(new_n296), .A4(new_n297), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n426), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n419), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n417), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n423), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n399), .B1(new_n428), .B2(new_n441), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n441), .A3(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(new_n399), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n366), .A2(new_n398), .A3(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n371), .A2(KEYINPUT35), .A3(new_n252), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n445), .A2(new_n448), .A3(new_n323), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n441), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n252), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n385), .A2(KEYINPUT87), .A3(new_n441), .A4(new_n428), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n323), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(KEYINPUT88), .A3(KEYINPUT35), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n447), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G43gat), .B(G50gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT15), .ZN(new_n462));
  NOR3_X1   g261(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(KEYINPUT90), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(KEYINPUT90), .B2(new_n464), .ZN(new_n466));
  NAND2_X1  g265(.A1(G29gat), .A2(G36gat), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n467), .B(KEYINPUT91), .Z(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n462), .ZN(new_n471));
  INV_X1    g270(.A(new_n464), .ZN(new_n472));
  OAI22_X1  g271(.A1(new_n461), .A2(KEYINPUT15), .B1(new_n472), .B2(new_n463), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n475), .A3(KEYINPUT17), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT16), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(G1gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(G1gat), .B2(new_n477), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n480), .B(G8gat), .Z(new_n481));
  INV_X1    g280(.A(KEYINPUT17), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n468), .B2(new_n474), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n476), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n468), .A2(new_n474), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n480), .B(G8gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT18), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n484), .A2(KEYINPUT18), .A3(new_n489), .A4(new_n485), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n485), .B(KEYINPUT13), .Z(new_n494));
  INV_X1    g293(.A(new_n489), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n487), .A2(new_n488), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G169gat), .B(G197gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT12), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n492), .A2(new_n493), .A3(new_n497), .A4(new_n504), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n460), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G57gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G64gat), .ZN(new_n512));
  INV_X1    g311(.A(G64gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(G57gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT9), .ZN(new_n516));
  INV_X1    g315(.A(G71gat), .ZN(new_n517));
  INV_X1    g316(.A(G78gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G71gat), .B(G78gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n515), .A2(new_n521), .A3(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G127gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n532));
  INV_X1    g331(.A(new_n524), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n521), .B1(new_n519), .B2(new_n515), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n523), .A2(KEYINPUT93), .A3(new_n524), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n481), .B1(new_n537), .B2(new_n526), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n531), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT92), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G155gat), .ZN(new_n542));
  XOR2_X1   g341(.A(G183gat), .B(G211gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n539), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G99gat), .ZN(new_n553));
  INV_X1    g352(.A(G106gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(KEYINPUT95), .A3(new_n549), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT96), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n549), .A2(KEYINPUT8), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  INV_X1    g359(.A(G92gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n557), .A2(new_n558), .A3(new_n563), .A4(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n550), .A2(new_n551), .A3(new_n548), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT95), .B1(new_n555), .B2(new_n549), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n563), .B(new_n567), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n559), .A2(new_n574), .A3(new_n562), .A4(new_n564), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(new_n552), .A3(new_n556), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(KEYINPUT96), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n476), .A2(new_n483), .A3(new_n568), .A4(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n568), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n487), .B2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G190gat), .B(G218gat), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n578), .B2(new_n581), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT94), .ZN(new_n589));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT97), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(KEYINPUT97), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n587), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n585), .B2(new_n586), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n547), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n577), .A2(new_n525), .A3(new_n568), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n571), .A2(new_n523), .A3(new_n576), .A4(new_n524), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n535), .B2(new_n536), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n580), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT99), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n607), .B1(new_n600), .B2(new_n602), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(KEYINPUT98), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n608), .B(new_n615), .C1(KEYINPUT98), .C2(new_n614), .ZN(new_n616));
  INV_X1    g415(.A(new_n607), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n603), .B2(new_n605), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n613), .B1(new_n618), .B2(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n599), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n202), .B1(new_n510), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n510), .A2(new_n202), .A3(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n365), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g426(.A1(new_n623), .A2(new_n624), .ZN(new_n628));
  OAI21_X1  g427(.A(G8gat), .B1(new_n628), .B2(new_n323), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT42), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n323), .B1(new_n623), .B2(new_n624), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT16), .B(G8gat), .Z(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(KEYINPUT101), .B2(new_n630), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n635), .B1(KEYINPUT101), .B2(new_n634), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n629), .A2(new_n633), .B1(new_n631), .B2(new_n636), .ZN(G1325gat));
  INV_X1    g436(.A(new_n445), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n628), .A2(G15gat), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(G15gat), .B1(new_n628), .B2(new_n446), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(G1326gat));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n252), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT43), .B(G22gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1327gat));
  NOR3_X1   g443(.A1(new_n547), .A2(new_n598), .A3(new_n620), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT102), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n460), .A2(new_n509), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(G29gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n648), .A3(new_n365), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT45), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n460), .B2(new_n598), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n455), .A2(KEYINPUT88), .A3(KEYINPUT35), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT88), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n653), .A2(new_n654), .A3(new_n449), .ZN(new_n655));
  OAI211_X1 g454(.A(KEYINPUT44), .B(new_n597), .C1(new_n655), .C2(new_n447), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n620), .B(KEYINPUT103), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n547), .A2(new_n659), .A3(new_n509), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n657), .A2(new_n365), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n650), .B1(new_n648), .B2(new_n661), .ZN(G1328gat));
  XOR2_X1   g461(.A(KEYINPUT104), .B(KEYINPUT46), .Z(new_n663));
  NOR2_X1   g462(.A1(new_n323), .A2(G36gat), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n647), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n647), .B2(new_n664), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n652), .A2(new_n656), .A3(new_n324), .A4(new_n660), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(G36gat), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT106), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n667), .B(new_n675), .C1(new_n671), .C2(new_n672), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(G1329gat));
  INV_X1    g476(.A(new_n446), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n652), .A2(new_n656), .A3(new_n678), .A4(new_n660), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G43gat), .ZN(new_n680));
  INV_X1    g479(.A(G43gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n647), .A2(new_n681), .A3(new_n445), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT47), .Z(G1330gat));
  NAND4_X1  g483(.A1(new_n652), .A2(new_n656), .A3(new_n252), .A4(new_n660), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G50gat), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT48), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(G50gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n647), .A2(new_n689), .A3(new_n252), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n688), .B(new_n691), .ZN(G1331gat));
  NOR4_X1   g491(.A1(new_n460), .A2(new_n508), .A3(new_n599), .A4(new_n658), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n365), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g494(.A(new_n323), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT108), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1333gat));
  AOI21_X1  g499(.A(new_n517), .B1(new_n693), .B2(new_n678), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n638), .A2(G71gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n693), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g503(.A1(new_n693), .A2(new_n252), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g505(.A1(new_n547), .A2(new_n508), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n620), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT109), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n657), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710), .B2(new_n453), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n597), .B(new_n707), .C1(new_n655), .C2(new_n447), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n460), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n715), .A2(KEYINPUT51), .A3(new_n597), .A4(new_n707), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n717), .A2(new_n560), .A3(new_n365), .A4(new_n620), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n718), .ZN(G1336gat));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n712), .A2(new_n720), .A3(new_n713), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n323), .A2(G92gat), .A3(new_n658), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n721), .B(new_n722), .C1(new_n717), .C2(new_n720), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n652), .A2(new_n656), .A3(new_n324), .A4(new_n709), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G92gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT52), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT52), .B1(new_n717), .B2(new_n722), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G92gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n724), .A2(new_n729), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n733), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n710), .B2(new_n446), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n553), .A3(new_n445), .A4(new_n620), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1338gat));
  NAND3_X1  g536(.A1(new_n657), .A2(new_n252), .A3(new_n709), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G106gat), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n385), .A2(new_n658), .A3(G106gat), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n721), .B(new_n740), .C1(new_n717), .C2(new_n720), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT53), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n717), .A2(new_n740), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n739), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1339gat));
  NAND2_X1  g546(.A1(new_n621), .A2(new_n509), .ZN(new_n748));
  INV_X1    g547(.A(new_n547), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n607), .B1(new_n604), .B2(new_n580), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n603), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n608), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n612), .B1(new_n618), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759));
  AND4_X1   g558(.A1(new_n759), .A2(new_n753), .A3(new_n755), .A4(KEYINPUT55), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n757), .B1(new_n608), .B2(new_n752), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(new_n761), .B2(new_n755), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n616), .B(new_n758), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT115), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n495), .A2(new_n496), .A3(new_n494), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n485), .B1(new_n484), .B2(new_n489), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n503), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n507), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n595), .B2(new_n596), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n603), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT54), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT55), .B1(new_n771), .B2(new_n618), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n618), .A2(new_n754), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n613), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT114), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n761), .A2(new_n759), .A3(new_n755), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n777), .A2(new_n778), .A3(new_n616), .A4(new_n758), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n764), .A2(new_n769), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n508), .A3(new_n779), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n507), .A2(new_n767), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n620), .ZN(new_n784));
  INV_X1    g583(.A(new_n620), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n768), .A2(new_n785), .A3(KEYINPUT116), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n780), .B1(new_n788), .B2(new_n598), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n749), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI211_X1 g590(.A(KEYINPUT117), .B(new_n780), .C1(new_n788), .C2(new_n598), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n748), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(KEYINPUT118), .B(new_n748), .C1(new_n791), .C2(new_n792), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n324), .A2(new_n453), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n638), .A2(new_n252), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n800), .B2(new_n509), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n797), .A2(new_n365), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(new_n323), .A3(new_n452), .A4(new_n454), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n508), .A2(new_n328), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(G1340gat));
  OAI21_X1  g604(.A(G120gat), .B1(new_n800), .B2(new_n658), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n620), .A2(new_n326), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT119), .Z(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n803), .B2(new_n808), .ZN(G1341gat));
  OAI21_X1  g608(.A(G127gat), .B1(new_n800), .B2(new_n749), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n547), .A2(new_n530), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n803), .B2(new_n811), .ZN(G1342gat));
  NOR2_X1   g611(.A1(new_n598), .A2(G134gat), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n803), .A2(KEYINPUT56), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G134gat), .B1(new_n800), .B2(new_n598), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT56), .B1(new_n803), .B2(new_n814), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(G1343gat));
  NAND3_X1  g617(.A1(new_n795), .A2(new_n252), .A3(new_n796), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n783), .A2(new_n620), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT120), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT55), .B1(new_n756), .B2(KEYINPUT121), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(KEYINPUT121), .B2(new_n756), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n508), .A3(new_n616), .A4(new_n777), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n597), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(KEYINPUT122), .ZN(new_n827));
  INV_X1    g626(.A(new_n780), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n826), .B2(KEYINPUT122), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n749), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n748), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n385), .A2(new_n820), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n819), .A2(new_n820), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n446), .A2(new_n798), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(new_n509), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(G141gat), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n678), .A2(new_n385), .A3(new_n324), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n802), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n508), .A2(new_n836), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT58), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843));
  OAI221_X1 g642(.A(new_n843), .B1(new_n839), .B2(new_n840), .C1(new_n835), .C2(new_n836), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1344gat));
  INV_X1    g644(.A(new_n839), .ZN(new_n846));
  INV_X1    g645(.A(G148gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n620), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n785), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n598), .A2(new_n763), .A3(new_n768), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n749), .B1(new_n826), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n748), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT57), .B1(new_n854), .B2(new_n252), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n795), .A2(new_n796), .A3(new_n832), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(KEYINPUT123), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n795), .A2(new_n858), .A3(new_n796), .A4(new_n832), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n851), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n847), .B1(new_n860), .B2(KEYINPUT124), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n856), .A2(KEYINPUT123), .ZN(new_n862));
  INV_X1    g661(.A(new_n855), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n850), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n849), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n833), .A2(new_n834), .ZN(new_n869));
  AOI211_X1 g668(.A(KEYINPUT59), .B(new_n847), .C1(new_n869), .C2(new_n620), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n848), .B1(new_n868), .B2(new_n870), .ZN(G1345gat));
  NAND3_X1  g670(.A1(new_n846), .A2(new_n204), .A3(new_n547), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n833), .A2(new_n749), .A3(new_n834), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n204), .B2(new_n873), .ZN(G1346gat));
  AOI21_X1  g673(.A(G162gat), .B1(new_n846), .B2(new_n597), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n598), .A2(new_n205), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n869), .B2(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n365), .A2(new_n323), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n795), .A2(new_n796), .A3(new_n799), .A4(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n265), .A3(new_n509), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n452), .A2(new_n324), .A3(new_n454), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n797), .A2(new_n453), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n508), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n880), .B1(new_n884), .B2(new_n265), .ZN(G1348gat));
  OAI21_X1  g684(.A(G176gat), .B1(new_n879), .B2(new_n658), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n620), .A2(new_n266), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n882), .B2(new_n887), .ZN(G1349gat));
  OAI21_X1  g687(.A(G183gat), .B1(new_n879), .B2(new_n749), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n547), .A2(new_n283), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g691(.A1(new_n883), .A2(new_n284), .A3(new_n597), .ZN(new_n893));
  OAI21_X1  g692(.A(G190gat), .B1(new_n879), .B2(new_n598), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT125), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(KEYINPUT125), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n893), .B1(new_n898), .B2(new_n899), .ZN(G1351gat));
  NAND2_X1  g699(.A1(new_n797), .A2(new_n453), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n446), .A2(new_n252), .A3(new_n324), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(G197gat), .B1(new_n903), .B2(new_n508), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n446), .A2(new_n878), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n905), .B1(new_n857), .B2(new_n859), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n508), .A2(G197gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1352gat));
  INV_X1    g707(.A(new_n903), .ZN(new_n909));
  INV_X1    g708(.A(G204gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n620), .A2(new_n910), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n909), .A2(KEYINPUT62), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT62), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n906), .A2(new_n659), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n912), .B(new_n913), .C1(new_n910), .C2(new_n914), .ZN(G1353gat));
  NAND3_X1  g714(.A1(new_n903), .A2(new_n217), .A3(new_n547), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n906), .A2(new_n547), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT63), .B1(new_n917), .B2(G211gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n919), .B(new_n217), .C1(new_n906), .C2(new_n547), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n916), .B1(new_n918), .B2(new_n920), .ZN(G1354gat));
  OAI21_X1  g720(.A(new_n218), .B1(new_n909), .B2(new_n598), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n924), .B(new_n218), .C1(new_n909), .C2(new_n598), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n597), .A2(G218gat), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT127), .Z(new_n927));
  AOI22_X1  g726(.A1(new_n923), .A2(new_n925), .B1(new_n906), .B2(new_n927), .ZN(G1355gat));
endmodule


