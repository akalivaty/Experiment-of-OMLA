//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n457), .A2(KEYINPUT68), .A3(G567), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n456), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n468), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(new_n473), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n472), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n467), .A2(G2105), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n476), .A2(new_n480), .A3(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT70), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n468), .A2(new_n471), .A3(G2105), .A4(new_n473), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n474), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(G136), .B2(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n468), .A2(new_n495), .A3(new_n471), .A4(new_n473), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n468), .A2(new_n471), .A3(G126), .A4(new_n473), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n472), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n477), .A2(new_n473), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n494), .A2(G2105), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT4), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n498), .A2(new_n501), .A3(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(G543), .B1(new_n516), .B2(new_n517), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n513), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n527), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT71), .B(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n515), .A2(new_n514), .ZN(new_n532));
  OAI21_X1  g107(.A(G89), .B1(new_n516), .B2(new_n517), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n518), .A2(new_n537), .B1(new_n520), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(G64), .B1(new_n515), .B2(new_n514), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n512), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AND2_X1   g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n510), .B2(G56), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n512), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n518), .A2(new_n547), .B1(new_n520), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n520), .B2(new_n556), .ZN(new_n557));
  OR2_X1    g132(.A1(KEYINPUT6), .A2(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(KEYINPUT6), .A2(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  INV_X1    g139(.A(G78), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n532), .A2(new_n564), .B1(new_n565), .B2(new_n507), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n558), .A2(new_n559), .B1(new_n508), .B2(new_n509), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G91), .ZN(new_n569));
  AND4_X1   g144(.A1(KEYINPUT72), .A2(new_n563), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n566), .A2(G651), .B1(new_n568), .B2(G91), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT72), .B1(new_n571), .B2(new_n563), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n570), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  OR2_X1    g149(.A1(new_n531), .A2(new_n535), .ZN(G286));
  NAND2_X1  g150(.A1(new_n568), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n507), .B1(new_n558), .B2(new_n559), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n568), .A2(G86), .B1(new_n578), .B2(G48), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n508), .B2(new_n509), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n586), .B(G61), .C1(new_n515), .C2(new_n514), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G61), .B1(new_n515), .B2(new_n514), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT73), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n594), .A2(new_n588), .A3(new_n583), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n595), .A2(KEYINPUT74), .A3(G651), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n582), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n593), .A2(KEYINPUT73), .B1(G73), .B2(G543), .ZN(new_n600));
  AOI211_X1 g175(.A(new_n591), .B(new_n512), .C1(new_n600), .C2(new_n588), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT74), .B1(new_n595), .B2(G651), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n598), .B(new_n581), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n599), .A2(new_n604), .ZN(G305));
  AOI22_X1  g180(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n512), .ZN(new_n607));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  INV_X1    g183(.A(G47), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n518), .A2(new_n608), .B1(new_n520), .B2(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n607), .A2(new_n610), .ZN(G290));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(G171), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT76), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n568), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n518), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n532), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n622), .A2(G651), .B1(G54), .B2(new_n578), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(KEYINPUT77), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(KEYINPUT77), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n614), .B1(new_n628), .B2(G868), .ZN(G284));
  OAI21_X1  g204(.A(new_n614), .B1(new_n628), .B2(G868), .ZN(G321));
  NAND2_X1  g205(.A1(G299), .A2(new_n612), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g207(.A(new_n631), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n628), .B1(new_n634), .B2(G860), .ZN(G148));
  INV_X1    g210(.A(new_n550), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(new_n612), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n627), .A2(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n502), .A2(new_n481), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n488), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(G135), .B2(new_n491), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(G2096), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n644), .A2(new_n651), .A3(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT78), .ZN(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n655), .B(new_n657), .Z(new_n658));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n658), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT17), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT80), .Z(new_n677));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n674), .B1(new_n671), .B2(new_n675), .ZN(new_n679));
  AOI22_X1  g254(.A1(new_n678), .A2(new_n679), .B1(new_n672), .B2(new_n675), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n678), .B2(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n673), .A2(new_n671), .A3(new_n675), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT18), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n677), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT81), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n688), .A2(new_n689), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n696), .A2(new_n692), .A3(new_n690), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n695), .B(new_n697), .C1(new_n692), .C2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n698), .B(new_n699), .ZN(new_n703));
  INV_X1    g278(.A(new_n701), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n707), .B1(new_n702), .B2(new_n705), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(G229));
  MUX2_X1   g286(.A(G6), .B(G305), .S(G16), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(G23), .ZN(new_n721));
  INV_X1    g296(.A(G288), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n716), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT33), .B(G1976), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n714), .A2(new_n715), .A3(new_n720), .A4(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT34), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(KEYINPUT34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n716), .A2(G24), .ZN(new_n729));
  INV_X1    g304(.A(G290), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n716), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G1986), .Z(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  OR2_X1    g309(.A1(G95), .A2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n736));
  INV_X1    g311(.A(G119), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n488), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G131), .B2(new_n491), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(new_n733), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n732), .B1(KEYINPUT82), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(KEYINPUT82), .B2(new_n743), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n727), .A2(new_n728), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT36), .ZN(new_n747));
  NAND2_X1  g322(.A1(G160), .A2(G29), .ZN(new_n748));
  INV_X1    g323(.A(G34), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT24), .ZN(new_n750));
  AOI21_X1  g325(.A(G29), .B1(new_n749), .B2(KEYINPUT24), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(KEYINPUT84), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT84), .B2(new_n751), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2084), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n491), .A2(G139), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT83), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n502), .A2(G127), .ZN(new_n759));
  INV_X1    g334(.A(G115), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n467), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(G103), .A2(G2104), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G2105), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n761), .A2(G2105), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(new_n733), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n733), .B2(G33), .ZN(new_n769));
  INV_X1    g344(.A(G2072), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n756), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n733), .A2(G32), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT26), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n776), .A2(new_n777), .B1(G105), .B2(new_n481), .ZN(new_n778));
  INV_X1    g353(.A(G129), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n488), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n491), .A2(G141), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT85), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n773), .B1(new_n784), .B2(new_n733), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT86), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n772), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n789), .A2(KEYINPUT87), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(KEYINPUT87), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n733), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n733), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT29), .Z(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G2090), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(G2090), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n785), .A2(new_n787), .ZN(new_n798));
  NAND2_X1  g373(.A1(G299), .A2(G16), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n716), .A2(G20), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT23), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT31), .B(G11), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT30), .B(G28), .Z(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G29), .ZN(new_n808));
  NOR2_X1   g383(.A1(G168), .A2(new_n716), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n716), .B2(G21), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT88), .B(G1966), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n716), .A2(G19), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n550), .B2(new_n716), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G1341), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n812), .B(new_n815), .C1(new_n810), .C2(new_n811), .ZN(new_n816));
  NAND2_X1  g391(.A1(G171), .A2(G16), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G5), .B2(G16), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT89), .B(G1961), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n818), .A2(new_n819), .B1(G29), .B2(new_n649), .ZN(new_n820));
  OAI221_X1 g395(.A(new_n820), .B1(G1341), .B2(new_n814), .C1(new_n818), .C2(new_n819), .ZN(new_n821));
  AOI211_X1 g396(.A(new_n816), .B(new_n821), .C1(new_n755), .C2(new_n754), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n733), .A2(G26), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT28), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n491), .A2(G140), .ZN(new_n825));
  OR2_X1    g400(.A1(G104), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n827));
  INV_X1    g402(.A(G128), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n488), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n830), .B2(new_n733), .ZN(new_n831));
  INV_X1    g406(.A(G2067), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(G27), .A2(G29), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G164), .B2(G29), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT90), .B(G2078), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n716), .A2(G4), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n628), .B2(new_n716), .ZN(new_n839));
  INV_X1    g414(.A(G1348), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n822), .A2(new_n833), .A3(new_n837), .A4(new_n841), .ZN(new_n842));
  NOR4_X1   g417(.A1(new_n790), .A2(new_n791), .A3(new_n805), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n747), .A2(new_n843), .ZN(G150));
  INV_X1    g419(.A(G150), .ZN(G311));
  NOR2_X1   g420(.A1(new_n627), .A2(new_n634), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n510), .A2(G67), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n512), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  INV_X1    g426(.A(G55), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n518), .A2(new_n851), .B1(new_n520), .B2(new_n852), .ZN(new_n853));
  OAI22_X1  g428(.A1(new_n546), .A2(new_n549), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G56), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n532), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(G651), .B1(new_n856), .B2(new_n544), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n568), .A2(G81), .B1(new_n578), .B2(G43), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n568), .A2(G93), .B1(new_n578), .B2(G55), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n849), .B1(new_n532), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G651), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n854), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n847), .B(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n850), .A2(new_n853), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n868), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(G145));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT93), .ZN(new_n876));
  INV_X1    g451(.A(G118), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(G2105), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n876), .B2(new_n875), .ZN(new_n879));
  INV_X1    g454(.A(G130), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n488), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(G142), .B2(new_n491), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n642), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(new_n739), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G164), .B(KEYINPUT91), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n782), .B1(new_n825), .B2(new_n829), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n830), .B1(new_n780), .B2(new_n781), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n889), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n767), .A2(KEYINPUT92), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT92), .B1(new_n767), .B2(new_n783), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n885), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n884), .A3(new_n895), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n649), .B(G160), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(G162), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n902), .B1(new_n898), .B2(new_n900), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g483(.A(new_n638), .B(new_n864), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n624), .B1(new_n570), .B2(new_n572), .ZN(new_n910));
  INV_X1    g485(.A(new_n624), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT72), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n557), .A2(new_n562), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n565), .A2(new_n507), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n510), .B2(G65), .ZN(new_n915));
  INV_X1    g490(.A(G91), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n915), .A2(new_n512), .B1(new_n916), .B2(new_n518), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n912), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n571), .A2(KEYINPUT72), .A3(new_n563), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n910), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n909), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(KEYINPUT94), .B(KEYINPUT41), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n910), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT41), .B1(new_n910), .B2(new_n920), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n909), .A2(new_n926), .ZN(new_n927));
  OR3_X1    g502(.A1(new_n922), .A2(new_n927), .A3(KEYINPUT95), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT95), .B1(new_n922), .B2(new_n927), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G303), .B(G288), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n581), .B1(new_n601), .B2(new_n602), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT75), .ZN(new_n933));
  AOI21_X1  g508(.A(G290), .B1(new_n933), .B2(new_n603), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n603), .A3(G290), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  INV_X1    g513(.A(new_n931), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n938), .A2(new_n934), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n930), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n942), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n928), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n612), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n871), .A2(G868), .ZN(new_n947));
  OR3_X1    g522(.A1(new_n946), .A2(KEYINPUT96), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT96), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(G295));
  INV_X1    g525(.A(KEYINPUT97), .ZN(new_n951));
  INV_X1    g526(.A(new_n946), .ZN(new_n952));
  INV_X1    g527(.A(new_n947), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n946), .A2(KEYINPUT97), .A3(new_n947), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(G331));
  OAI21_X1  g531(.A(KEYINPUT98), .B1(new_n539), .B2(new_n542), .ZN(new_n957));
  INV_X1    g532(.A(G64), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n508), .B2(new_n509), .ZN(new_n959));
  INV_X1    g534(.A(new_n541), .ZN(new_n960));
  OAI21_X1  g535(.A(G651), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT98), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n578), .A2(G52), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n560), .A2(new_n510), .A3(G90), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(G286), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(G171), .A2(new_n962), .A3(G168), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n966), .A2(new_n967), .B1(new_n854), .B2(new_n863), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n966), .A2(new_n854), .A3(new_n967), .A4(new_n863), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n921), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(KEYINPUT99), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT99), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n864), .A2(new_n974), .A3(new_n967), .A4(new_n966), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n968), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT100), .B1(new_n926), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT41), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n570), .A2(new_n572), .A3(new_n624), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n918), .A2(new_n919), .B1(new_n619), .B2(new_n623), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n910), .A2(new_n920), .A3(new_n923), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT100), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n970), .B(new_n974), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n983), .B(new_n984), .C1(new_n985), .C2(new_n968), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n972), .B1(new_n977), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n904), .B1(new_n987), .B2(new_n941), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n941), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n937), .A2(new_n940), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n921), .A2(new_n923), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n969), .A2(new_n970), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n993), .B(new_n994), .C1(KEYINPUT41), .C2(new_n921), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n921), .A2(new_n969), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n985), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G37), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n998), .A2(new_n989), .ZN(new_n999));
  OAI221_X1 g574(.A(KEYINPUT44), .B1(new_n988), .B2(new_n991), .C1(new_n999), .C2(new_n990), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n977), .A2(new_n986), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n1001), .A2(new_n941), .A3(new_n971), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n988), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n989), .A3(new_n990), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT101), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT101), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n1008), .B(KEYINPUT44), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1000), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT102), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT102), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1012), .B(new_n1000), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(G397));
  NAND2_X1  g589(.A1(new_n496), .A2(new_n497), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n472), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n499), .A2(new_n500), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G2105), .ZN(new_n1018));
  INV_X1    g593(.A(new_n504), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT103), .B(G40), .Z(new_n1024));
  NOR4_X1   g599(.A1(new_n476), .A2(new_n480), .A3(new_n482), .A4(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1996), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n784), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n830), .B(G2067), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1029), .B(new_n1030), .C1(new_n1028), .C2(new_n782), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n739), .B(new_n742), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT104), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G290), .B(G1986), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1027), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n501), .A2(new_n504), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n1038), .B2(new_n1016), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1025), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT105), .B(G2090), .Z(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1023), .B1(G164), .B2(G1384), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1020), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1025), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n719), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1037), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(G166), .B2(new_n1037), .ZN(new_n1052));
  NAND3_X1  g627(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1053));
  NAND2_X1  g628(.A1(KEYINPUT110), .A2(G8), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1037), .B(new_n1055), .C1(new_n1045), .C2(new_n1049), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT106), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n1062), .B(new_n1037), .C1(new_n1039), .C2(new_n1025), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1025), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT106), .B1(new_n1064), .B2(G8), .ZN(new_n1065));
  OAI221_X1 g640(.A(new_n1061), .B1(new_n1060), .B2(G288), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1062), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(KEYINPUT106), .A3(G8), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1069), .A2(new_n1070), .B1(G1976), .B2(new_n722), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1073));
  INV_X1    g648(.A(G1981), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n590), .B2(new_n581), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1074), .B(new_n581), .C1(new_n601), .C2(new_n602), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT107), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n592), .A2(new_n596), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(KEYINPUT107), .A3(new_n1074), .A4(new_n581), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1075), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1073), .B1(new_n1081), .B2(KEYINPUT49), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1083), .B(new_n1075), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT108), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1075), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT107), .B1(new_n597), .B2(new_n1074), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1083), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT108), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1081), .A2(KEYINPUT49), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1073), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1072), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1059), .B1(new_n1094), .B2(KEYINPUT111), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1072), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1089), .B2(new_n1083), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1091), .B1(new_n1098), .B2(new_n1092), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1082), .A2(KEYINPUT108), .A3(new_n1084), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1966), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1048), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1025), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1042), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1105), .B1(new_n1109), .B2(G2084), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G8), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G286), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1095), .A2(new_n1103), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1050), .B(new_n1116), .Z(new_n1117));
  NAND4_X1  g692(.A1(new_n1117), .A2(KEYINPUT63), .A3(new_n1094), .A4(new_n1112), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(KEYINPUT111), .B(new_n1096), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1059), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1094), .A2(KEYINPUT111), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT122), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1095), .A2(new_n1103), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G168), .A2(new_n1037), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(KEYINPUT51), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1043), .A2(new_n755), .B1(new_n1104), .B2(new_n1048), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n1037), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1110), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1127), .B(KEYINPUT120), .Z(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n1111), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1127), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n1134), .A2(new_n1137), .B1(new_n1131), .B2(new_n1138), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT62), .ZN(new_n1140));
  INV_X1    g715(.A(G1961), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1109), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1048), .B2(G2078), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(G2078), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1046), .A2(new_n1025), .A3(new_n1047), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G171), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1139), .B2(KEYINPUT62), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1124), .A2(new_n1126), .A3(new_n1140), .A4(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1094), .A2(new_n1050), .A3(new_n1116), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G288), .A2(G1976), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1153), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1097), .B1(new_n1157), .B2(KEYINPUT109), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT109), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1159), .B(new_n1153), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1119), .A2(new_n1151), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1128), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1137), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1163), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(G160), .A2(G40), .A3(new_n1146), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1046), .A2(new_n1047), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1145), .A2(G301), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT54), .B1(new_n1149), .B2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1142), .A2(new_n1144), .A3(G301), .A4(new_n1147), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT54), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1145), .A2(KEYINPUT123), .A3(new_n1169), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1142), .A2(new_n1144), .A3(new_n1169), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n1176));
  AOI21_X1  g751(.A(G301), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1173), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1167), .A2(new_n1171), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1124), .A2(new_n1179), .A3(new_n1126), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n803), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1181));
  OAI211_X1 g756(.A(KEYINPUT112), .B(KEYINPUT57), .C1(new_n913), .C2(new_n917), .ZN(new_n1182));
  NAND2_X1  g757(.A1(KEYINPUT112), .A2(KEYINPUT57), .ZN(new_n1183));
  OR2_X1    g758(.A1(KEYINPUT112), .A2(KEYINPUT57), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n571), .A2(new_n563), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(KEYINPUT56), .B(G2072), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1046), .A2(new_n1025), .A3(new_n1047), .A4(new_n1188), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1181), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1186), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT113), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1187), .B1(new_n1181), .B2(new_n1189), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT113), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n840), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1039), .A2(new_n832), .A3(new_n1025), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n911), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1190), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT60), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT119), .B1(new_n1204), .B2(new_n911), .ZN(new_n1205));
  AOI21_X1  g780(.A(KEYINPUT60), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT119), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1206), .A2(new_n1207), .A3(new_n624), .ZN(new_n1208));
  OAI22_X1  g783(.A1(new_n1205), .A2(new_n1208), .B1(new_n1203), .B2(new_n1200), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1204), .A2(KEYINPUT119), .A3(new_n911), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1207), .B1(new_n1206), .B2(new_n624), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1209), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1046), .A2(new_n1028), .A3(new_n1047), .A4(new_n1025), .ZN(new_n1215));
  XOR2_X1   g790(.A(KEYINPUT58), .B(G1341), .Z(new_n1216));
  NAND2_X1  g791(.A1(new_n1064), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n550), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(KEYINPUT115), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT59), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1221), .A2(KEYINPUT114), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT115), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1218), .A2(new_n1224), .A3(new_n550), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1220), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1224), .B1(new_n1218), .B2(new_n550), .ZN(new_n1227));
  AOI211_X1 g802(.A(KEYINPUT115), .B(new_n636), .C1(new_n1215), .C2(new_n1217), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1222), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1181), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1231));
  NAND4_X1  g806(.A1(new_n1193), .A2(KEYINPUT61), .A3(new_n1196), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1192), .A2(new_n1231), .ZN(new_n1233));
  XOR2_X1   g808(.A(KEYINPUT116), .B(KEYINPUT61), .Z(new_n1234));
  AOI21_X1  g809(.A(KEYINPUT117), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g810(.A(KEYINPUT117), .B(new_n1234), .C1(new_n1190), .C2(new_n1194), .ZN(new_n1236));
  INV_X1    g811(.A(new_n1236), .ZN(new_n1237));
  OAI211_X1 g812(.A(new_n1230), .B(new_n1232), .C1(new_n1235), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1214), .B1(new_n1238), .B2(KEYINPUT118), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1240));
  INV_X1    g815(.A(KEYINPUT117), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1242), .A2(new_n1236), .ZN(new_n1243));
  INV_X1    g818(.A(KEYINPUT118), .ZN(new_n1244));
  NAND4_X1  g819(.A1(new_n1243), .A2(new_n1244), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1245));
  AOI21_X1  g820(.A(new_n1202), .B1(new_n1239), .B2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g821(.A1(new_n1180), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g822(.A(new_n1036), .B1(new_n1162), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g823(.A1(new_n1026), .A2(G1996), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1249), .A2(KEYINPUT46), .ZN(new_n1250));
  XNOR2_X1  g825(.A(new_n1250), .B(KEYINPUT125), .ZN(new_n1251));
  AND2_X1   g826(.A1(new_n1030), .A2(new_n782), .ZN(new_n1252));
  OAI221_X1 g827(.A(new_n1251), .B1(KEYINPUT46), .B2(new_n1249), .C1(new_n1026), .C2(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g828(.A(new_n1253), .B(KEYINPUT126), .ZN(new_n1254));
  OR2_X1    g829(.A1(new_n1254), .A2(KEYINPUT47), .ZN(new_n1255));
  NAND2_X1  g830(.A1(new_n1254), .A2(KEYINPUT47), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n739), .A2(new_n741), .ZN(new_n1257));
  XNOR2_X1  g832(.A(new_n1257), .B(KEYINPUT124), .ZN(new_n1258));
  OR2_X1    g833(.A1(new_n1031), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n830), .A2(new_n832), .ZN(new_n1260));
  AOI21_X1  g835(.A(new_n1026), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1034), .A2(new_n1027), .ZN(new_n1262));
  NOR3_X1   g837(.A1(new_n1026), .A2(G1986), .A3(G290), .ZN(new_n1263));
  XOR2_X1   g838(.A(new_n1263), .B(KEYINPUT48), .Z(new_n1264));
  AOI21_X1  g839(.A(new_n1261), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  AND3_X1   g840(.A1(new_n1255), .A2(new_n1256), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1248), .A2(new_n1266), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g842(.A1(G227), .A2(new_n465), .ZN(new_n1269));
  OAI211_X1 g843(.A(new_n669), .B(new_n1269), .C1(new_n709), .C2(new_n710), .ZN(new_n1270));
  NOR2_X1   g844(.A1(new_n907), .A2(new_n1270), .ZN(new_n1271));
  AND3_X1   g845(.A1(new_n1271), .A2(KEYINPUT127), .A3(new_n1005), .ZN(new_n1272));
  AOI21_X1  g846(.A(KEYINPUT127), .B1(new_n1271), .B2(new_n1005), .ZN(new_n1273));
  NOR2_X1   g847(.A1(new_n1272), .A2(new_n1273), .ZN(G308));
  NAND2_X1  g848(.A1(new_n1271), .A2(new_n1005), .ZN(new_n1275));
  INV_X1    g849(.A(KEYINPUT127), .ZN(new_n1276));
  NAND2_X1  g850(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g851(.A1(new_n1271), .A2(KEYINPUT127), .A3(new_n1005), .ZN(new_n1278));
  NAND2_X1  g852(.A1(new_n1277), .A2(new_n1278), .ZN(G225));
endmodule


