//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1325, new_n1326,
    new_n1327, new_n1329, new_n1330, new_n1331, new_n1332, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421, new_n1422, new_n1423, new_n1424, new_n1425,
    new_n1426;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n209), .B1(new_n203), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n208), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g0021(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n204), .A2(new_n205), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n208), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT0), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n218), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n217), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G97), .B(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  OAI21_X1  g0052(.A(KEYINPUT69), .B1(new_n225), .B2(G1), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n255), .A3(G20), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n228), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n221), .A2(new_n259), .A3(new_n222), .A4(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n259), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n258), .A2(new_n262), .B1(new_n228), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n221), .A2(new_n222), .A3(new_n260), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT8), .B(G58), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n225), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G150), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n265), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n221), .A2(new_n222), .B1(G33), .B2(G41), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G223), .A3(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G77), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n277), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n286), .A2(G222), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n276), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  AND2_X1   g0089(.A1(G1), .A2(G13), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT68), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n255), .C1(G41), .C2(G45), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n296), .B1(new_n301), .B2(G226), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n288), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  AOI211_X1 g0105(.A(new_n275), .B(new_n304), .C1(new_n305), .C2(new_n303), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(G200), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n288), .A2(G190), .A3(new_n302), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT73), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n264), .B2(new_n273), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n264), .A2(new_n312), .A3(new_n273), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n315), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n317), .A2(KEYINPUT9), .A3(new_n313), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n310), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT9), .B1(new_n317), .B2(new_n313), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(new_n311), .A3(new_n315), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(new_n310), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n306), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT75), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n268), .A2(new_n279), .B1(new_n225), .B2(G68), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(KEYINPUT74), .B1(new_n228), .B2(new_n271), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n328), .A2(KEYINPUT74), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n327), .B(new_n265), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(KEYINPUT74), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT74), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n334), .B1(new_n225), .B2(G68), .C1(new_n268), .C2(new_n279), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n335), .C1(new_n228), .C2(new_n271), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n327), .B1(new_n336), .B2(new_n265), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT11), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n265), .B1(new_n329), .B2(new_n330), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT75), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT11), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n331), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n263), .A2(new_n203), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT12), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT76), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n257), .A2(new_n203), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n262), .ZN(new_n347));
  NOR4_X1   g0147(.A1(new_n257), .A2(new_n261), .A3(KEYINPUT76), .A4(new_n203), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n338), .A2(new_n342), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT77), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n340), .A2(new_n331), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n349), .B1(new_n353), .B2(KEYINPUT11), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT77), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n342), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n277), .A2(G232), .A3(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n277), .A2(new_n285), .ZN(new_n359));
  INV_X1    g0159(.A(G226), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n276), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n296), .B1(new_n301), .B2(G238), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT13), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n362), .B2(new_n363), .ZN(new_n366));
  OAI21_X1  g0166(.A(G169), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n363), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n367), .A2(KEYINPUT14), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n371), .B2(G169), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n352), .B(new_n356), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(G200), .B1(new_n365), .B2(new_n366), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n369), .A2(G190), .A3(new_n370), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n351), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT72), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT15), .B(G87), .Z(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  INV_X1    g0184(.A(new_n268), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT15), .B(G87), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT71), .B1(new_n387), .B2(new_n268), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT8), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G58), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n270), .B1(G20), .B2(G77), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT70), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n386), .B(new_n388), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n267), .A2(new_n271), .B1(new_n225), .B2(new_n279), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n396), .A2(KEYINPUT70), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n265), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n253), .A2(new_n256), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G77), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n400), .A2(new_n261), .B1(G77), .B2(new_n259), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G200), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n277), .A2(G232), .A3(new_n285), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n277), .A2(G238), .A3(G1698), .ZN(new_n406));
  INV_X1    g0206(.A(G107), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(new_n277), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n276), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n296), .B1(new_n301), .B2(G244), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n404), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n382), .B1(new_n403), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G200), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(KEYINPUT72), .A3(new_n398), .A4(new_n402), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n409), .A2(new_n410), .A3(G190), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n305), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n409), .A2(new_n410), .A3(new_n372), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n403), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n326), .A2(new_n376), .A3(new_n381), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n399), .A2(new_n392), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n425), .A2(new_n261), .B1(new_n259), .B2(new_n392), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(G20), .B1(G159), .B2(new_n270), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT7), .ZN(new_n430));
  AOI211_X1 g0230(.A(new_n430), .B(G20), .C1(new_n282), .C2(new_n284), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n283), .A2(G33), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT78), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT78), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n282), .A2(new_n284), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n225), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n431), .B1(new_n437), .B2(new_n430), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT16), .B(new_n429), .C1(new_n438), .C2(new_n203), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT16), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n428), .A2(G20), .ZN(new_n442));
  INV_X1    g0242(.A(G159), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(new_n271), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n430), .B1(new_n277), .B2(G20), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n282), .A2(new_n284), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n203), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n441), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n265), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n427), .B1(new_n440), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n297), .A2(G232), .A3(new_n298), .A4(new_n300), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n295), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n282), .A2(new_n284), .A3(G226), .A4(G1698), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n282), .A2(new_n284), .A3(G223), .A4(new_n285), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G87), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n453), .B1(new_n276), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n372), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n458), .A2(G169), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n452), .A2(new_n295), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n457), .A2(new_n276), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n372), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n460), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n451), .A2(new_n466), .A3(KEYINPUT18), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT80), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n451), .A2(new_n466), .A3(new_n469), .A4(KEYINPUT18), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT18), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n459), .B1(new_n458), .B2(new_n372), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n462), .A2(new_n463), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n305), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n221), .A2(new_n222), .A3(new_n260), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT7), .B1(new_n446), .B2(new_n225), .ZN(new_n478));
  OAI21_X1  g0278(.A(G68), .B1(new_n478), .B2(new_n431), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n429), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n480), .B2(new_n441), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n426), .B1(new_n481), .B2(new_n439), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n471), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n468), .A2(new_n470), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n439), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n404), .B1(new_n462), .B2(new_n463), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(G190), .B2(new_n458), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n487), .A3(new_n427), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT17), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n482), .A2(KEYINPUT17), .A3(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT81), .B1(new_n424), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n376), .A2(new_n423), .A3(new_n381), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT81), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT18), .B1(new_n451), .B2(new_n466), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(KEYINPUT80), .B2(new_n467), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n499), .B2(new_n470), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n496), .A2(new_n497), .A3(new_n500), .A4(new_n326), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G41), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n255), .B(G45), .C1(new_n503), .C2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(G41), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n505), .A2(new_n292), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n508), .A2(G41), .ZN(new_n511));
  OAI211_X1 g0311(.A(G264), .B(new_n298), .C1(new_n504), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT91), .ZN(new_n513));
  INV_X1    g0313(.A(G45), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G1), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(G41), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT91), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(G264), .A4(new_n298), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n212), .A2(new_n285), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(G257), .B2(new_n285), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n523), .A2(new_n446), .B1(new_n281), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n276), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n521), .A2(KEYINPUT92), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT92), .B1(new_n521), .B2(new_n526), .ZN(new_n528));
  OAI211_X1 g0328(.A(G179), .B(new_n510), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n512), .A3(new_n510), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n225), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n407), .A2(KEYINPUT23), .A3(G20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n225), .A2(G33), .A3(G116), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n277), .A2(new_n225), .A3(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n277), .A2(new_n541), .A3(new_n225), .A4(G87), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n265), .B1(new_n543), .B2(KEYINPUT24), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n261), .B1(new_n255), .B2(G33), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n259), .A2(G107), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT25), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n547), .A2(KEYINPUT90), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT90), .B1(new_n547), .B2(new_n549), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n544), .A2(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n532), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n552), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n510), .B1(new_n527), .B2(new_n528), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(KEYINPUT93), .A3(new_n404), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n530), .A2(G190), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT93), .B1(new_n555), .B2(new_n404), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n546), .A2(G97), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n259), .A2(G97), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT6), .ZN(new_n566));
  INV_X1    g0366(.A(G97), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(new_n407), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n407), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n225), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n271), .A2(new_n279), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n565), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n478), .B2(new_n431), .ZN(new_n575));
  INV_X1    g0375(.A(new_n573), .ZN(new_n576));
  INV_X1    g0376(.A(new_n571), .ZN(new_n577));
  XNOR2_X1  g0377(.A(G97), .B(G107), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(new_n566), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(KEYINPUT82), .B(new_n576), .C1(new_n579), .C2(new_n225), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n574), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n564), .B1(new_n581), .B2(new_n265), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT83), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n286), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(G244), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n282), .A2(new_n284), .A3(G250), .A4(G1698), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G283), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n286), .A2(G244), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n276), .ZN(new_n595));
  OAI211_X1 g0395(.A(G257), .B(new_n298), .C1(new_n504), .C2(new_n511), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT85), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n518), .A2(KEYINPUT85), .A3(G257), .A4(new_n298), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n510), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(G190), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n276), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n587), .B2(new_n593), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(KEYINPUT86), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT86), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n600), .A2(new_n607), .A3(new_n510), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n582), .B(new_n603), .C1(new_n609), .C2(new_n404), .ZN(new_n610));
  INV_X1    g0410(.A(new_n608), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n607), .B1(new_n600), .B2(new_n510), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n595), .B(new_n372), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n581), .A2(new_n265), .ZN(new_n614));
  INV_X1    g0414(.A(new_n564), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n305), .B1(new_n605), .B2(new_n601), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n255), .A2(G45), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n298), .A2(G250), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n298), .A2(G274), .A3(new_n515), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT87), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT87), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n292), .A2(new_n624), .A3(new_n515), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n621), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n282), .A2(new_n284), .A3(G244), .A4(G1698), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n282), .A2(new_n284), .A3(G238), .A4(new_n285), .ZN(new_n628));
  NAND2_X1  g0428(.A1(G33), .A2(G116), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n276), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n372), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n626), .A2(new_n631), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n211), .A2(KEYINPUT88), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G87), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n637), .A3(new_n569), .ZN(new_n638));
  NAND3_X1  g0438(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n225), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n282), .A2(new_n284), .A3(new_n225), .A4(G68), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT19), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n268), .B2(new_n567), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n645), .A2(new_n265), .B1(new_n263), .B2(new_n387), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n546), .A2(new_n383), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n305), .A2(new_n634), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n404), .B1(new_n626), .B2(new_n631), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n642), .A2(new_n644), .ZN(new_n650));
  XNOR2_X1  g0450(.A(KEYINPUT88), .B(G87), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(new_n569), .B1(new_n225), .B2(new_n639), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n265), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n387), .A2(new_n263), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n255), .A2(G33), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n262), .A2(G87), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n649), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n632), .A2(G190), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n633), .A2(new_n648), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(G270), .B(new_n298), .C1(new_n504), .C2(new_n511), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n510), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(G257), .A2(G1698), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n285), .A2(G264), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n277), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G303), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n446), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n276), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n305), .B1(new_n663), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n477), .A2(G116), .A3(new_n259), .A4(new_n655), .ZN(new_n671));
  INV_X1    g0471(.A(G116), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n263), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(G20), .B1(G33), .B2(G283), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n281), .A2(G97), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(G20), .B2(new_n672), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n676), .A2(new_n265), .A3(KEYINPUT20), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT20), .B1(new_n676), .B2(new_n265), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n671), .B(new_n673), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT21), .B1(new_n670), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n669), .A2(new_n510), .A3(new_n661), .ZN(new_n681));
  AND4_X1   g0481(.A1(KEYINPUT21), .A2(new_n679), .A3(G169), .A4(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  INV_X1    g0484(.A(new_n679), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n669), .A2(G179), .A3(new_n510), .A4(new_n661), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n686), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(KEYINPUT89), .A3(new_n679), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(G200), .ZN(new_n691));
  INV_X1    g0491(.A(G190), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n685), .B(new_n691), .C1(new_n692), .C2(new_n681), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n660), .A2(new_n683), .A3(new_n690), .A4(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n619), .A2(new_n694), .ZN(new_n695));
  AND4_X1   g0495(.A1(new_n502), .A2(new_n553), .A3(new_n560), .A4(new_n695), .ZN(G372));
  AND2_X1   g0496(.A1(new_n483), .A2(new_n467), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n355), .B1(new_n354), .B2(new_n342), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n355), .A2(new_n338), .A3(new_n342), .A4(new_n350), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n371), .A2(new_n374), .A3(G169), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n702), .B(new_n703), .C1(new_n372), .C2(new_n371), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n701), .A2(new_n704), .B1(new_n381), .B2(new_n422), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n698), .B1(new_n705), .B2(new_n492), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n320), .A2(new_n325), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n306), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n502), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n634), .A2(G200), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT94), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT94), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n649), .B2(new_n657), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n659), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n648), .A2(new_n633), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n679), .A2(G169), .A3(new_n681), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT21), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n670), .A2(KEYINPUT21), .A3(new_n679), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n688), .A2(KEYINPUT89), .A3(new_n679), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT89), .B1(new_n688), .B2(new_n679), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n721), .B(new_n722), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n718), .B1(new_n726), .B2(new_n553), .ZN(new_n727));
  INV_X1    g0527(.A(new_n619), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n727), .A2(new_n560), .A3(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n716), .A2(new_n717), .ZN(new_n730));
  INV_X1    g0530(.A(new_n618), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT26), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n660), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT26), .B1(new_n734), .B2(new_n618), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(new_n717), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n709), .B1(new_n710), .B2(new_n737), .ZN(G369));
  NAND3_X1  g0538(.A1(new_n255), .A2(new_n225), .A3(G13), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT95), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n739), .A2(new_n740), .A3(KEYINPUT27), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n740), .B1(new_n739), .B2(KEYINPUT27), .ZN(new_n742));
  OAI221_X1 g0542(.A(G213), .B1(KEYINPUT27), .B2(new_n739), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G343), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n553), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n552), .A2(new_n745), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n560), .A2(new_n553), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n553), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n745), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT96), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n748), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n726), .A2(new_n745), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n746), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n745), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n685), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n726), .A2(new_n693), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n726), .B2(new_n760), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n762), .A2(G330), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n755), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n764), .ZN(G399));
  NOR2_X1   g0565(.A1(new_n638), .A2(G116), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n231), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G41), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n767), .A2(new_n255), .A3(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n770), .A2(KEYINPUT97), .B1(new_n229), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(KEYINPUT97), .B2(new_n770), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT28), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT29), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n737), .B2(new_n745), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n619), .A2(KEYINPUT98), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT98), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n610), .A2(new_n618), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n776), .A2(new_n727), .A3(new_n560), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(KEYINPUT26), .B1(new_n718), .B2(new_n618), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n595), .A2(new_n602), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n582), .B1(new_n305), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n782), .A2(new_n660), .A3(new_n732), .A4(new_n613), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n780), .A2(new_n717), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n745), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(KEYINPUT29), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n775), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT30), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n634), .A2(new_n686), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n527), .B2(new_n528), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n788), .B1(new_n790), .B2(new_n781), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n595), .B1(new_n611), .B2(new_n612), .ZN(new_n792));
  AND3_X1   g0592(.A1(new_n634), .A2(new_n372), .A3(new_n681), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n792), .A2(new_n555), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n528), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n521), .A2(KEYINPUT92), .A3(new_n526), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n605), .A2(new_n601), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT30), .A4(new_n789), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n791), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g0600(.A1(new_n800), .A2(KEYINPUT31), .A3(new_n745), .ZN(new_n801));
  AOI21_X1  g0601(.A(KEYINPUT31), .B1(new_n800), .B2(new_n745), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n695), .A2(new_n553), .A3(new_n560), .A4(new_n758), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G330), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n787), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n773), .B1(new_n809), .B2(G1), .ZN(G364));
  NOR2_X1   g0610(.A1(new_n762), .A2(G330), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT99), .Z(new_n812));
  INV_X1    g0612(.A(new_n763), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n225), .A2(G13), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n255), .B1(new_n814), .B2(G45), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n769), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n812), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n768), .A2(new_n446), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G355), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(G116), .B2(new_n231), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n282), .A2(new_n284), .A3(new_n435), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n435), .B1(new_n282), .B2(new_n284), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n768), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n514), .B2(new_n229), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n247), .A2(new_n514), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n822), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n224), .B1(G20), .B2(new_n305), .ZN(new_n832));
  NOR2_X1   g0632(.A1(G13), .A2(G33), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(G20), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n817), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n832), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n225), .A2(new_n372), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(G190), .A3(new_n404), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT100), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n841), .A2(KEYINPUT100), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT101), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n404), .B2(G179), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n372), .A2(KEYINPUT101), .A3(G200), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n225), .A2(G190), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n846), .A2(G322), .B1(G283), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n840), .A2(G200), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n692), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G326), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n840), .A2(new_n692), .A3(G200), .ZN(new_n858));
  XOR2_X1   g0658(.A(KEYINPUT33), .B(G317), .Z(new_n859));
  OAI22_X1  g0659(.A1(new_n856), .A2(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(G179), .A2(G200), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n225), .B1(new_n861), .B2(G190), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n860), .B1(G294), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n850), .A2(new_n861), .ZN(new_n865));
  INV_X1    g0665(.A(G329), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n840), .A2(new_n692), .A3(new_n404), .ZN(new_n867));
  INV_X1    g0667(.A(G311), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n446), .B1(new_n865), .B2(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n225), .A2(new_n692), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n848), .A2(new_n870), .A3(new_n849), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n869), .B1(G303), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n853), .A2(new_n864), .A3(new_n873), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n856), .A2(new_n228), .B1(new_n203), .B2(new_n858), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n865), .A2(new_n443), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(KEYINPUT32), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n862), .A2(new_n567), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n875), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n846), .A2(G58), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n277), .B1(new_n867), .B2(new_n279), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(KEYINPUT32), .B2(new_n877), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n871), .A2(new_n651), .B1(new_n851), .B2(new_n407), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n880), .A2(new_n881), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n839), .B1(new_n874), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n838), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n835), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n762), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n819), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G396));
  INV_X1    g0692(.A(new_n808), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n421), .A2(KEYINPUT102), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n419), .A2(new_n403), .A3(new_n895), .A4(new_n420), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n418), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n758), .B(new_n898), .C1(new_n729), .C2(new_n736), .ZN(new_n899));
  INV_X1    g0699(.A(new_n736), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n727), .A2(new_n560), .A3(new_n728), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n745), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n403), .A2(new_n745), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n417), .A2(new_n903), .A3(new_n894), .A4(new_n896), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n422), .A2(new_n745), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n899), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n817), .B1(new_n893), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n893), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n839), .A2(new_n834), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n817), .B1(new_n910), .B2(G77), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n846), .A2(G294), .B1(G87), .B2(new_n852), .ZN(new_n912));
  INV_X1    g0712(.A(G283), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n858), .A2(new_n913), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n879), .B(new_n914), .C1(G303), .C2(new_n855), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n446), .B1(new_n865), .B2(new_n868), .C1(new_n867), .C2(new_n672), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(G107), .B2(new_n872), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n867), .ZN(new_n919));
  AOI22_X1  g0719(.A1(G137), .A2(new_n855), .B1(new_n919), .B2(G159), .ZN(new_n920));
  INV_X1    g0720(.A(G143), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n920), .B1(new_n269), .B2(new_n858), .C1(new_n845), .C2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT34), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(G132), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n826), .B1(new_n202), .B2(new_n862), .C1(new_n925), .C2(new_n865), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(G50), .A2(new_n872), .B1(new_n852), .B2(G68), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n922), .A2(new_n923), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n918), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n911), .B1(new_n931), .B2(new_n832), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n906), .B2(new_n834), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n909), .A2(new_n933), .ZN(G384));
  NAND3_X1  g0734(.A1(new_n502), .A2(new_n775), .A3(new_n786), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n935), .A2(new_n709), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT104), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT7), .B1(new_n825), .B2(new_n225), .ZN(new_n939));
  OAI21_X1  g0739(.A(G68), .B1(new_n939), .B2(new_n431), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT16), .B1(new_n940), .B2(new_n429), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n439), .A2(new_n265), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n427), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n743), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n484), .B2(new_n493), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT37), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n943), .A2(new_n466), .B1(new_n482), .B2(new_n487), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n948), .B2(new_n945), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n488), .B1(new_n476), .B2(new_n482), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n482), .A2(new_n743), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n950), .A2(KEYINPUT37), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n938), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n451), .A2(new_n466), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n451), .A2(new_n944), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n955), .A2(new_n956), .A3(new_n947), .A4(new_n488), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n429), .B1(new_n438), .B2(new_n203), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n441), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(new_n439), .A3(new_n265), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n473), .A2(new_n475), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n960), .A2(new_n427), .B1(new_n961), .B2(new_n460), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n743), .B1(new_n960), .B2(new_n427), .ZN(new_n963));
  INV_X1    g0763(.A(new_n488), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n957), .B1(new_n965), .B2(new_n947), .ZN(new_n966));
  OAI211_X1 g0766(.A(KEYINPUT38), .B(new_n966), .C1(new_n500), .C2(new_n945), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT103), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n954), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(KEYINPUT103), .B(new_n938), .C1(new_n946), .C2(new_n953), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT39), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n376), .A2(new_n745), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n951), .B1(new_n697), .B2(new_n492), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT37), .B1(new_n950), .B2(new_n951), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n957), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n938), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT39), .B1(new_n967), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n972), .A2(new_n973), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n352), .A2(new_n356), .A3(new_n745), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n376), .A2(new_n381), .A3(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n701), .B(new_n745), .C1(new_n704), .C2(new_n380), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n897), .A2(new_n758), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n986), .B1(new_n899), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(new_n969), .A3(new_n970), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n697), .A2(new_n743), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n981), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n937), .B(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n906), .ZN(new_n995));
  AOI221_X4 g0795(.A(new_n995), .B1(new_n983), .B2(new_n984), .C1(new_n803), .C2(new_n804), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT40), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n969), .A2(new_n996), .A3(new_n997), .A4(new_n970), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT38), .B1(new_n974), .B2(new_n976), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n946), .A2(new_n953), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(KEYINPUT38), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n805), .A2(new_n906), .A3(new_n985), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT40), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n710), .A2(new_n806), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1007), .A2(new_n1008), .A3(new_n807), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n994), .A2(new_n1009), .B1(new_n255), .B2(new_n814), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n994), .B2(new_n1009), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n579), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT35), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT35), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1013), .A2(G116), .A3(new_n226), .A4(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT36), .Z(new_n1016));
  OAI211_X1 g0816(.A(new_n229), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n228), .A2(G68), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n255), .B(G13), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1011), .A2(new_n1016), .A3(new_n1019), .ZN(G367));
  NOR2_X1   g0820(.A1(new_n828), .A2(new_n243), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n836), .B1(new_n231), .B2(new_n387), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n817), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n846), .A2(G150), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n858), .A2(new_n443), .B1(new_n862), .B2(new_n203), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G143), .B2(new_n855), .ZN(new_n1026));
  INV_X1    g0826(.A(G137), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n277), .B1(new_n865), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G50), .B2(new_n919), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G58), .A2(new_n872), .B1(new_n852), .B2(G77), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1024), .A2(new_n1026), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n856), .A2(new_n868), .B1(new_n862), .B2(new_n407), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n858), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1032), .B1(G294), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(G317), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n867), .A2(new_n913), .B1(new_n865), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n826), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n846), .A2(G303), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n852), .A2(G97), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n871), .A2(new_n672), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT46), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1031), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT47), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1023), .B1(new_n1044), .B2(new_n832), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n745), .A2(new_n657), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n730), .A2(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n717), .A2(new_n1046), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1045), .B1(new_n1049), .B2(new_n889), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT109), .Z(new_n1051));
  INV_X1    g0851(.A(new_n809), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT44), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT106), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n748), .A2(new_n753), .A3(new_n750), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n753), .B1(new_n748), .B2(new_n750), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n756), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n746), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n776), .A2(new_n778), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n616), .A2(new_n745), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n618), .B2(new_n758), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1054), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(KEYINPUT106), .B(new_n1063), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1053), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT108), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n764), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT45), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n757), .A2(KEYINPUT45), .A3(new_n1063), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT106), .B1(new_n757), .B2(new_n1063), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1059), .A2(new_n1054), .A3(new_n1064), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(KEYINPUT44), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1067), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n764), .A2(new_n1068), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1067), .A2(new_n1073), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1057), .A2(KEYINPUT107), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(new_n763), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n755), .A2(new_n756), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1052), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n769), .B(KEYINPUT41), .Z(new_n1090));
  OAI21_X1  g0890(.A(new_n815), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n755), .A2(new_n1063), .A3(new_n763), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT105), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1049), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT43), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n755), .A2(new_n1063), .A3(new_n756), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT42), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1060), .A2(new_n749), .A3(new_n1061), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n745), .B1(new_n1101), .B2(new_n618), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1099), .B2(KEYINPUT42), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1098), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(KEYINPUT43), .B2(new_n1049), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1100), .A2(new_n1103), .A3(new_n1097), .A4(new_n1096), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1095), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1094), .B(new_n1093), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1051), .B1(new_n1091), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G387));
  NAND2_X1  g0913(.A1(new_n1088), .A2(new_n816), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n755), .A2(new_n889), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G303), .A2(new_n919), .B1(new_n1033), .B2(G311), .ZN(new_n1116));
  INV_X1    g0916(.A(G322), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n856), .C1(new_n845), .C2(new_n1035), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT48), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n872), .A2(G294), .B1(G283), .B2(new_n863), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT49), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n825), .B1(new_n672), .B2(new_n851), .C1(new_n857), .C2(new_n865), .ZN(new_n1127));
  OR3_X1    g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n846), .A2(G50), .B1(G77), .B2(new_n872), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n863), .A2(new_n383), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n267), .B2(new_n858), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G159), .B2(new_n855), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n867), .A2(new_n203), .B1(new_n865), .B2(new_n269), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(new_n825), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1129), .A2(new_n1039), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n839), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n828), .B1(new_n240), .B2(G45), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n767), .B2(new_n820), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n267), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT50), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n392), .B2(new_n228), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n514), .B1(new_n203), .B2(new_n279), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n767), .A2(new_n1139), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1138), .A2(new_n1143), .B1(G107), .B2(new_n231), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n818), .B(new_n1136), .C1(new_n836), .C2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT110), .Z(new_n1146));
  NOR2_X1   g0946(.A1(new_n1088), .A2(new_n809), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1087), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n809), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n769), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1114), .B1(new_n1115), .B2(new_n1146), .C1(new_n1147), .C2(new_n1151), .ZN(G393));
  NAND2_X1  g0952(.A1(new_n1082), .A2(new_n816), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n837), .B1(G97), .B2(new_n768), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n827), .A2(new_n251), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n818), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n845), .A2(new_n868), .B1(new_n1035), .B2(new_n856), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT52), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n446), .B1(new_n865), .B2(new_n1117), .C1(new_n867), .C2(new_n524), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n871), .A2(new_n913), .B1(new_n851), .B2(new_n407), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n858), .A2(new_n667), .B1(new_n862), .B2(new_n672), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n845), .A2(new_n443), .B1(new_n269), .B2(new_n856), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT51), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n871), .A2(new_n203), .B1(new_n851), .B2(new_n211), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n867), .A2(new_n267), .B1(new_n865), .B2(new_n921), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n858), .A2(new_n228), .B1(new_n862), .B2(new_n279), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n825), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1158), .A2(new_n1162), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1156), .B1(new_n839), .B2(new_n1169), .C1(new_n1063), .C2(new_n889), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1052), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1082), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n769), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1082), .A2(new_n1171), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1153), .B(new_n1170), .C1(new_n1173), .C2(new_n1174), .ZN(G390));
  NAND2_X1  g0975(.A1(new_n502), .A2(new_n808), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n935), .A2(new_n709), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT114), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT114), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n935), .A2(new_n1176), .A3(new_n1179), .A4(new_n709), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n995), .B1(new_n803), .B2(new_n804), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(G330), .A3(new_n985), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n985), .B1(new_n1181), .B2(G330), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n902), .A2(new_n898), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n987), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n1183), .A2(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1184), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n785), .B2(new_n898), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n1182), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1178), .A2(new_n1180), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT112), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1189), .A2(new_n986), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n967), .A2(new_n978), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n973), .B(KEYINPUT111), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1193), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1196), .B1(new_n967), .B2(new_n978), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1200), .B(KEYINPUT112), .C1(new_n986), .C2(new_n1189), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT39), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n969), .B2(new_n970), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1204), .A2(new_n979), .B1(new_n973), .B2(new_n988), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1182), .A2(KEYINPUT113), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1202), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1206), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1192), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1206), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1202), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1178), .A2(new_n1180), .A3(new_n1191), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1209), .A2(new_n1215), .A3(new_n769), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n979), .B1(new_n971), .B2(KEYINPUT39), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(new_n834), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n867), .A2(new_n567), .B1(new_n865), .B2(new_n524), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n856), .A2(new_n913), .B1(new_n407), .B2(new_n858), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(G77), .C2(new_n863), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n203), .B2(new_n851), .C1(new_n672), .C2(new_n845), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n446), .B1(new_n871), .B2(new_n211), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT117), .Z(new_n1224));
  NOR2_X1   g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT118), .ZN(new_n1226));
  INV_X1    g1026(.A(G128), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n845), .A2(new_n925), .B1(new_n1227), .B2(new_n856), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT115), .Z(new_n1229));
  NOR2_X1   g1029(.A1(new_n871), .A2(new_n269), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT53), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n858), .A2(new_n1027), .B1(new_n862), .B2(new_n443), .ZN(new_n1232));
  INV_X1    g1032(.A(G125), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(KEYINPUT54), .B(G143), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n277), .B1(new_n865), .B2(new_n1233), .C1(new_n867), .C2(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1232), .B(new_n1235), .C1(G50), .C2(new_n852), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1229), .A2(new_n1231), .A3(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT116), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n839), .B1(new_n1226), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n817), .B1(new_n910), .B2(new_n392), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1218), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1242), .B2(new_n816), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1216), .A2(new_n1243), .ZN(G378));
  INV_X1    g1044(.A(KEYINPUT119), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n743), .B1(new_n314), .B2(new_n315), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n707), .B2(new_n306), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1246), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n326), .A2(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1004), .B2(G330), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n807), .B(new_n1253), .C1(new_n998), .C2(new_n1003), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n993), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n991), .B1(new_n973), .B2(new_n1217), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1004), .A2(G330), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1253), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1004), .A2(G330), .A3(new_n1254), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1245), .B1(new_n1257), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1258), .A3(new_n1261), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n993), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(KEYINPUT119), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n816), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1253), .A2(new_n833), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n817), .B1(new_n910), .B2(G50), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n856), .A2(new_n672), .B1(new_n567), .B2(new_n858), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n826), .B(new_n1270), .C1(G68), .C2(new_n863), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n503), .B1(new_n865), .B2(new_n913), .C1(new_n867), .C2(new_n387), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G77), .B2(new_n872), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n852), .A2(G58), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n846), .A2(G107), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1271), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT58), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n503), .B1(new_n825), .B2(new_n281), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1276), .A2(new_n1277), .B1(new_n228), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1234), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n846), .A2(G128), .B1(new_n872), .B2(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(G125), .A2(new_n855), .B1(new_n919), .B2(G137), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1033), .A2(G132), .B1(new_n863), .B2(G150), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(KEYINPUT59), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(KEYINPUT59), .ZN(new_n1286));
  INV_X1    g1086(.A(G124), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n281), .B(new_n503), .C1(new_n865), .C2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G159), .B2(new_n852), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n1279), .B1(new_n1277), .B2(new_n1276), .C1(new_n1285), .C2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1269), .B1(new_n1291), .B2(new_n832), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1268), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1267), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1209), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1263), .A3(new_n1266), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT57), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n769), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1299), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1297), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1294), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(G375));
  NAND2_X1  g1105(.A1(new_n986), .A2(new_n833), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n817), .B1(new_n910), .B2(G68), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n846), .A2(G137), .B1(G159), .B2(new_n872), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n856), .A2(new_n925), .B1(new_n862), .B2(new_n228), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1033), .B2(new_n1280), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n867), .A2(new_n269), .B1(new_n865), .B2(new_n1227), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(new_n825), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1308), .A2(new_n1310), .A3(new_n1274), .A4(new_n1312), .ZN(new_n1313));
  OAI221_X1 g1113(.A(new_n1130), .B1(new_n672), .B2(new_n858), .C1(new_n856), .C2(new_n524), .ZN(new_n1314));
  OAI221_X1 g1114(.A(new_n446), .B1(new_n865), .B2(new_n667), .C1(new_n867), .C2(new_n407), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(G77), .B2(new_n852), .ZN(new_n1316));
  OAI221_X1 g1116(.A(new_n1316), .B1(new_n567), .B2(new_n871), .C1(new_n913), .C2(new_n845), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1313), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1307), .B1(new_n1318), .B2(new_n832), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n1191), .A2(new_n816), .B1(new_n1306), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1090), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1214), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1191), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1320), .B1(new_n1322), .B2(new_n1323), .ZN(G381));
  NOR3_X1   g1124(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(KEYINPUT120), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(G390), .A2(G378), .A3(G381), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(new_n1112), .A3(new_n1304), .A4(new_n1327), .ZN(G407));
  INV_X1    g1128(.A(G378), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n744), .A2(G213), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1304), .A2(new_n1329), .A3(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(G407), .A2(G213), .A3(new_n1332), .ZN(G409));
  NAND4_X1  g1133(.A1(new_n1295), .A2(KEYINPUT60), .A3(new_n1187), .A4(new_n1190), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n769), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1323), .B1(KEYINPUT60), .B2(new_n1214), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1320), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(G384), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  OAI211_X1 g1139(.A(G384), .B(new_n1320), .C1(new_n1335), .C2(new_n1336), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1331), .A2(KEYINPUT121), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(G2897), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1342), .B1(new_n1343), .B2(new_n1330), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1330), .A2(new_n1343), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1339), .A2(new_n1340), .A3(new_n1345), .A4(new_n1341), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1297), .A2(new_n1263), .A3(new_n1321), .A4(new_n1266), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1293), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1349), .B1(new_n1350), .B2(new_n816), .ZN(new_n1351));
  AOI21_X1  g1151(.A(G378), .B1(new_n1348), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1352), .B1(new_n1304), .B2(G378), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1347), .B1(new_n1353), .B2(new_n1331), .ZN(new_n1354));
  AND3_X1   g1154(.A1(new_n1264), .A2(new_n1265), .A3(KEYINPUT119), .ZN(new_n1355));
  AOI21_X1  g1155(.A(KEYINPUT119), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1349), .B1(new_n1357), .B2(new_n816), .ZN(new_n1358));
  AOI21_X1  g1158(.A(KEYINPUT57), .B1(new_n1357), .B2(new_n1297), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1295), .B1(new_n1242), .B2(new_n1192), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1350), .A2(KEYINPUT57), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n769), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1362));
  OAI211_X1 g1162(.A(G378), .B(new_n1358), .C1(new_n1359), .C2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1352), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT62), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1367), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1365), .A2(new_n1366), .A3(new_n1330), .A4(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT61), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1354), .A2(new_n1369), .A3(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1331), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1366), .B1(new_n1372), .B2(new_n1368), .ZN(new_n1373));
  OAI21_X1  g1173(.A(KEYINPUT124), .B1(new_n1371), .B2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1373), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1365), .A2(new_n1330), .ZN(new_n1376));
  AOI21_X1  g1176(.A(KEYINPUT61), .B1(new_n1376), .B2(new_n1347), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT124), .ZN(new_n1378));
  NAND4_X1  g1178(.A1(new_n1375), .A2(new_n1377), .A3(new_n1378), .A4(new_n1369), .ZN(new_n1379));
  XNOR2_X1  g1179(.A(G393), .B(new_n891), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1091), .A2(new_n1111), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1051), .ZN(new_n1382));
  AOI21_X1  g1182(.A(G390), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT122), .ZN(new_n1384));
  OAI21_X1  g1184(.A(new_n1380), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1385));
  INV_X1    g1185(.A(G390), .ZN(new_n1386));
  INV_X1    g1186(.A(new_n1111), .ZN(new_n1387));
  AOI21_X1  g1187(.A(new_n1150), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1321), .B1(new_n1388), .B2(new_n1052), .ZN(new_n1389));
  AOI21_X1  g1189(.A(new_n1387), .B1(new_n1389), .B2(new_n815), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1386), .B1(new_n1390), .B2(new_n1051), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1112), .A2(G390), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1391), .A2(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1385), .A2(new_n1393), .ZN(new_n1394));
  NAND4_X1  g1194(.A1(new_n1391), .A2(new_n1392), .A3(new_n1380), .A4(new_n1384), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1394), .A2(new_n1395), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1374), .A2(new_n1379), .A3(new_n1396), .ZN(new_n1397));
  NAND3_X1  g1197(.A1(new_n1394), .A2(new_n1370), .A3(new_n1395), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1398), .A2(KEYINPUT123), .ZN(new_n1399));
  AND3_X1   g1199(.A1(new_n1372), .A2(KEYINPUT63), .A3(new_n1368), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1372), .A2(new_n1368), .ZN(new_n1401));
  XNOR2_X1  g1201(.A(new_n1342), .B(new_n1345), .ZN(new_n1402));
  OAI21_X1  g1202(.A(KEYINPUT63), .B1(new_n1372), .B2(new_n1402), .ZN(new_n1403));
  AOI21_X1  g1203(.A(new_n1400), .B1(new_n1401), .B2(new_n1403), .ZN(new_n1404));
  INV_X1    g1204(.A(KEYINPUT123), .ZN(new_n1405));
  NAND4_X1  g1205(.A1(new_n1394), .A2(new_n1405), .A3(new_n1370), .A4(new_n1395), .ZN(new_n1406));
  NAND3_X1  g1206(.A1(new_n1399), .A2(new_n1404), .A3(new_n1406), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1397), .A2(new_n1407), .ZN(G405));
  AOI21_X1  g1208(.A(new_n1362), .B1(new_n1299), .B2(new_n1298), .ZN(new_n1409));
  OAI21_X1  g1209(.A(new_n1329), .B1(new_n1409), .B2(new_n1294), .ZN(new_n1410));
  NAND3_X1  g1210(.A1(new_n1410), .A2(new_n1363), .A3(new_n1367), .ZN(new_n1411));
  AND2_X1   g1211(.A1(new_n1411), .A2(KEYINPUT126), .ZN(new_n1412));
  NOR2_X1   g1212(.A1(new_n1411), .A2(KEYINPUT126), .ZN(new_n1413));
  NAND2_X1  g1213(.A1(new_n1410), .A2(new_n1363), .ZN(new_n1414));
  AOI21_X1  g1214(.A(KEYINPUT125), .B1(new_n1414), .B2(new_n1368), .ZN(new_n1415));
  INV_X1    g1215(.A(KEYINPUT125), .ZN(new_n1416));
  AOI211_X1 g1216(.A(new_n1416), .B(new_n1367), .C1(new_n1410), .C2(new_n1363), .ZN(new_n1417));
  OAI22_X1  g1217(.A1(new_n1412), .A2(new_n1413), .B1(new_n1415), .B2(new_n1417), .ZN(new_n1418));
  INV_X1    g1218(.A(KEYINPUT127), .ZN(new_n1419));
  NAND2_X1  g1219(.A1(new_n1396), .A2(new_n1419), .ZN(new_n1420));
  NAND3_X1  g1220(.A1(new_n1394), .A2(KEYINPUT127), .A3(new_n1395), .ZN(new_n1421));
  NAND3_X1  g1221(.A1(new_n1418), .A2(new_n1420), .A3(new_n1421), .ZN(new_n1422));
  OR2_X1    g1222(.A1(new_n1415), .A2(new_n1417), .ZN(new_n1423));
  INV_X1    g1223(.A(new_n1396), .ZN(new_n1424));
  XNOR2_X1  g1224(.A(new_n1411), .B(KEYINPUT126), .ZN(new_n1425));
  NAND4_X1  g1225(.A1(new_n1423), .A2(new_n1424), .A3(KEYINPUT127), .A4(new_n1425), .ZN(new_n1426));
  NAND2_X1  g1226(.A1(new_n1422), .A2(new_n1426), .ZN(G402));
endmodule


