//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT67), .B(G128), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G143), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n191), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n200), .B2(KEYINPUT65), .ZN(new_n201));
  AOI21_X1  g015(.A(G143), .B1(new_n190), .B2(new_n192), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n194), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n189), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n193), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n187), .B1(new_n205), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n213));
  INV_X1    g027(.A(new_n188), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n195), .B1(new_n202), .B2(new_n203), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT64), .B(G146), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n217), .A2(KEYINPUT65), .A3(G143), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n210), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n221), .A2(KEYINPUT81), .A3(KEYINPUT3), .A4(G104), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n221), .A2(KEYINPUT81), .A3(G104), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n221), .B2(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n222), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(G104), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G107), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n227), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n212), .A2(new_n220), .A3(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT0), .B(G128), .Z(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n216), .B2(new_n218), .ZN(new_n239));
  OAI211_X1 g053(.A(G101), .B(new_n222), .C1(new_n223), .C2(new_n225), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n228), .A2(new_n240), .A3(KEYINPUT4), .ZN(new_n241));
  OR3_X1    g055(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n206), .B1(new_n217), .B2(G143), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT0), .A3(G128), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n239), .A2(new_n241), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G134), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(KEYINPUT11), .A3(G134), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G131), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n208), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n210), .B1(new_n243), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT82), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n232), .B1(new_n226), .B2(new_n227), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n235), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n237), .A2(new_n245), .A3(new_n255), .A4(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n219), .A2(new_n210), .A3(new_n234), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n260), .B2(new_n261), .ZN(new_n265));
  INV_X1    g079(.A(new_n255), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n265), .A2(KEYINPUT12), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT12), .B1(new_n265), .B2(new_n266), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OR2_X1    g083(.A1(KEYINPUT70), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT70), .A2(G953), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G227), .ZN(new_n273));
  XOR2_X1   g087(.A(G110), .B(G140), .Z(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n237), .A2(new_n245), .A3(new_n262), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n266), .ZN(new_n278));
  INV_X1    g092(.A(new_n275), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n263), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G469), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT83), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n263), .A2(new_n279), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n278), .A2(new_n285), .B1(new_n269), .B2(new_n275), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n284), .B(G469), .C1(new_n286), .C2(G902), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n267), .B2(new_n268), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n278), .A2(new_n263), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n275), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT84), .B(G469), .Z(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n283), .A2(new_n287), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G221), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n298), .B2(new_n292), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n295), .A2(KEYINPUT85), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT91), .ZN(new_n306));
  INV_X1    g120(.A(G119), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G116), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G119), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT5), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT5), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n307), .A3(G116), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G113), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT86), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT5), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT86), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G113), .A4(new_n313), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n308), .A2(new_n310), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT2), .B(G113), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT87), .B1(new_n324), .B2(new_n234), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n323), .A2(new_n318), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n259), .A4(new_n315), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n322), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n241), .A2(new_n242), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n325), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT6), .ZN(new_n335));
  XNOR2_X1  g149(.A(G110), .B(G122), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n334), .A2(new_n337), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n325), .A2(new_n328), .A3(new_n333), .A4(new_n336), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT6), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT88), .B(new_n338), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n334), .A2(new_n337), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT88), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT6), .A4(new_n340), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n239), .A2(new_n244), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT74), .B(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(KEYINPUT74), .A2(G125), .ZN(new_n350));
  NOR2_X1   g164(.A1(KEYINPUT74), .A2(G125), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n219), .A2(new_n352), .A3(new_n210), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G224), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G953), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n349), .B2(new_n353), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n346), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G210), .B1(G237), .B2(G902), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n349), .A2(KEYINPUT89), .A3(new_n353), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(KEYINPUT7), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n353), .B2(KEYINPUT89), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n340), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n349), .A2(KEYINPUT7), .A3(new_n353), .A4(new_n358), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n323), .B1(new_n311), .B2(new_n314), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n259), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n336), .B(KEYINPUT8), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n371), .B(new_n372), .C1(new_n324), .C2(new_n259), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n292), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n362), .A2(new_n363), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n378));
  INV_X1    g192(.A(new_n363), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n360), .B1(new_n342), .B2(new_n345), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n362), .A2(KEYINPUT90), .A3(new_n363), .A4(new_n376), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G214), .B1(G237), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n306), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(KEYINPUT91), .A3(new_n383), .A4(new_n385), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G475), .ZN(new_n390));
  INV_X1    g204(.A(G237), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n270), .A2(G214), .A3(new_n391), .A4(new_n271), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n392), .A2(new_n197), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n197), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G131), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT17), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n254), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n352), .A2(KEYINPUT16), .A3(G140), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT75), .ZN(new_n402));
  OAI21_X1  g216(.A(G140), .B1(new_n350), .B2(new_n351), .ZN(new_n403));
  NOR2_X1   g217(.A1(G125), .A2(G140), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n402), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT16), .ZN(new_n408));
  AOI211_X1 g222(.A(KEYINPUT75), .B(new_n408), .C1(new_n403), .C2(new_n405), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n401), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n189), .ZN(new_n411));
  OAI211_X1 g225(.A(G146), .B(new_n401), .C1(new_n407), .C2(new_n409), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n395), .A2(KEYINPUT17), .A3(G131), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n399), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT18), .A2(G131), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT93), .B1(new_n395), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n393), .A2(new_n418), .A3(new_n394), .A4(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G125), .B(G140), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n217), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n404), .B1(new_n348), .B2(G140), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G146), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n395), .A2(new_n416), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n414), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(new_n230), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n414), .A2(new_n429), .A3(new_n426), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n390), .B1(new_n433), .B2(new_n292), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n421), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(KEYINPUT19), .B2(new_n423), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n396), .A2(new_n398), .B1(new_n217), .B2(new_n439), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n412), .A2(new_n440), .B1(new_n420), .B2(new_n425), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n429), .B1(new_n441), .B2(KEYINPUT94), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n412), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n426), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT94), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n427), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n442), .A2(new_n446), .B1(new_n447), .B2(new_n429), .ZN(new_n448));
  NOR2_X1   g262(.A1(G475), .A2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n436), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n430), .B1(new_n444), .B2(new_n445), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n441), .A2(KEYINPUT94), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n432), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n449), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n434), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT95), .B1(new_n458), .B2(G116), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT95), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n309), .A3(G122), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n309), .B2(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(G107), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n197), .A2(G128), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT96), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n188), .A2(G143), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n251), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n466), .A2(new_n470), .B1(G143), .B2(new_n188), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n251), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G217), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n297), .A2(new_n476), .A3(G953), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n462), .A2(KEYINPUT14), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n462), .A2(KEYINPUT14), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n309), .B2(G122), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n480), .B2(KEYINPUT97), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(KEYINPUT97), .B2(new_n480), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n482), .A2(G107), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n466), .A2(new_n467), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G134), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n251), .B1(new_n466), .B2(new_n467), .ZN(new_n486));
  OAI22_X1  g300(.A1(new_n485), .A2(new_n486), .B1(G107), .B2(new_n463), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n475), .B(new_n477), .C1(new_n483), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n477), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n482), .B2(G107), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n489), .B1(new_n490), .B2(new_n474), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n492), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G952), .ZN(new_n498));
  AOI211_X1 g312(.A(G953), .B(new_n498), .C1(G234), .C2(G237), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n292), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(G898), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n457), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n305), .A2(new_n389), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n253), .A2(G131), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n247), .A2(new_n252), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(G131), .C1(new_n508), .C2(new_n247), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n212), .A2(new_n512), .A3(new_n220), .ZN(new_n513));
  INV_X1    g327(.A(new_n347), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n266), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT30), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n347), .A2(new_n255), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n511), .B1(new_n219), .B2(new_n210), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n516), .A2(new_n332), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n332), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n515), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n272), .A2(G210), .A3(new_n391), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT27), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT26), .B(G101), .Z(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT31), .B1(new_n521), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n332), .B1(new_n518), .B2(new_n519), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT28), .A4(new_n522), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n527), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n516), .A2(new_n332), .A3(new_n520), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n528), .A4(new_n523), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NOR2_X1   g355(.A1(G472), .A2(G902), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G472), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n528), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n537), .A2(new_n527), .A3(new_n523), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n513), .A2(new_n515), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n332), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n527), .A2(new_n550), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n532), .A2(new_n552), .A3(new_n534), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n292), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n549), .A2(new_n550), .B1(KEYINPUT71), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n555), .A2(KEYINPUT71), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n546), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT72), .B1(new_n545), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n540), .A2(new_n542), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT32), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n549), .A2(new_n550), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n555), .A2(KEYINPUT71), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n557), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G472), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT72), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n476), .B1(G234), .B2(new_n292), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT22), .B(G137), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g387(.A1(G221), .A2(G234), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n272), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n270), .A2(new_n271), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT76), .B1(new_n578), .B2(new_n574), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n576), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n582), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n571), .A3(new_n580), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT73), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT67), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G128), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n590), .A3(G119), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n307), .A2(G128), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n587), .A3(new_n592), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT24), .B(G110), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT23), .B1(new_n208), .B2(G119), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n307), .B2(G128), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G110), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n411), .B2(new_n412), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n591), .A2(new_n587), .A3(new_n592), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n596), .B1(new_n606), .B2(new_n593), .ZN(new_n607));
  INV_X1    g421(.A(G110), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n599), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n412), .A2(new_n610), .A3(new_n422), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n586), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT78), .ZN(new_n613));
  INV_X1    g427(.A(new_n604), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT75), .B1(new_n423), .B2(new_n408), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n406), .A2(new_n402), .A3(KEYINPUT16), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(G146), .B1(new_n617), .B2(new_n401), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n189), .B(new_n400), .C1(new_n615), .C2(new_n616), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n412), .A2(new_n610), .A3(new_n422), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT78), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n586), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n583), .A2(new_n585), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT79), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n620), .A2(KEYINPUT79), .A3(new_n621), .A4(new_n625), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n613), .A2(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT25), .B1(new_n630), .B2(new_n292), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n613), .A2(new_n624), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n628), .A2(new_n629), .ZN(new_n633));
  AND4_X1   g447(.A1(KEYINPUT25), .A2(new_n632), .A3(new_n633), .A4(new_n292), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n570), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n570), .A2(G902), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT80), .ZN(new_n637));
  INV_X1    g451(.A(new_n630), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n559), .A2(new_n569), .A3(new_n640), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n506), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G101), .ZN(G3));
  NAND2_X1  g457(.A1(new_n540), .A2(new_n292), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G472), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n560), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n305), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n386), .B1(new_n377), .B2(new_n381), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n503), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n491), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n488), .A2(new_n491), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n488), .B(new_n491), .C1(new_n652), .C2(new_n651), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(G478), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n492), .A2(new_n493), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n493), .A2(new_n292), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n650), .A2(new_n457), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n648), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND3_X1  g479(.A1(new_n454), .A2(new_n435), .A3(new_n449), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n451), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n434), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n650), .A2(new_n497), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n648), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n221), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  INV_X1    g488(.A(new_n570), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n632), .A2(new_n633), .A3(new_n292), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT25), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n630), .A2(KEYINPUT25), .A3(new_n292), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n586), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n622), .ZN(new_n682));
  INV_X1    g496(.A(new_n637), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT100), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n635), .A2(new_n687), .A3(new_n684), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n646), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n305), .A2(new_n389), .A3(new_n505), .A4(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  NAND2_X1  g506(.A1(new_n686), .A2(new_n688), .ZN(new_n693));
  INV_X1    g507(.A(new_n499), .ZN(new_n694));
  INV_X1    g508(.A(new_n500), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n694), .B1(new_n695), .B2(G900), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n667), .A2(new_n496), .A3(new_n668), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n377), .A2(new_n381), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n385), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n305), .A3(new_n559), .A4(new_n569), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT101), .B(G128), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G30));
  XNOR2_X1  g518(.A(new_n696), .B(KEYINPUT39), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n305), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n384), .B(KEYINPUT38), .Z(new_n709));
  AOI21_X1  g523(.A(new_n527), .B1(new_n537), .B2(new_n523), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n552), .A2(new_n527), .A3(new_n523), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT102), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n292), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT102), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n563), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n457), .A2(new_n497), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n385), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n717), .A2(new_n693), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n708), .A2(new_n709), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n706), .A2(new_n707), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n197), .ZN(G45));
  AND2_X1   g538(.A1(new_n559), .A2(new_n569), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n457), .A2(new_n661), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n696), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n699), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n725), .A2(new_n305), .A3(new_n693), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AOI21_X1  g544(.A(G902), .B1(new_n288), .B2(new_n290), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n294), .B(new_n300), .C1(new_n282), .C2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n559), .A2(new_n569), .A3(new_n640), .A4(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n662), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT41), .B(G113), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  INV_X1    g552(.A(new_n670), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n309), .ZN(G18));
  NOR3_X1   g555(.A1(new_n504), .A2(new_n732), .A3(new_n699), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n559), .A3(new_n569), .A4(new_n693), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  AND3_X1   g558(.A1(new_n532), .A2(new_n552), .A3(new_n534), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n530), .B(new_n539), .C1(new_n528), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n542), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n645), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n639), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n699), .A2(new_n457), .A3(new_n497), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n503), .A4(new_n733), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  NAND2_X1  g566(.A1(new_n733), .A2(new_n649), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n727), .ZN(new_n754));
  AOI211_X1 g568(.A(KEYINPUT103), .B(new_n748), .C1(new_n686), .C2(new_n688), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT103), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n645), .A2(new_n747), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n756), .B1(new_n693), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  OAI21_X1  g574(.A(G469), .B1(new_n286), .B2(G902), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n299), .B1(new_n294), .B2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n384), .A2(new_n385), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n727), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n639), .B1(new_n563), .B2(new_n567), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(KEYINPUT42), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n559), .A2(new_n763), .A3(new_n569), .A4(new_n640), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n727), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n768), .B1(new_n770), .B2(KEYINPUT42), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT104), .B(G131), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G33));
  INV_X1    g587(.A(new_n769), .ZN(new_n774));
  INV_X1    g588(.A(new_n697), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n693), .A2(new_n646), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n661), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n457), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT43), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n778), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n276), .A2(new_n280), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n282), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n286), .A2(KEYINPUT45), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(G469), .A2(G902), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT46), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n294), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n791), .A2(new_n792), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n300), .B(new_n705), .C1(new_n795), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT105), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n798), .A2(new_n794), .A3(new_n793), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT105), .A3(new_n300), .A4(new_n705), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n779), .B(KEYINPUT106), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(KEYINPUT44), .A3(new_n784), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n384), .A2(new_n385), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n786), .A2(new_n804), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n795), .A2(new_n798), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n812), .B2(new_n299), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n802), .A2(KEYINPUT47), .A3(new_n300), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n640), .A2(new_n807), .A3(new_n727), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n559), .A2(new_n569), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT107), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT107), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n815), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(G140), .Z(G42));
  NAND3_X1  g637(.A1(new_n640), .A2(new_n385), .A3(new_n300), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT108), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n294), .B1(new_n282), .B2(new_n731), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n783), .A3(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT109), .Z(new_n829));
  OR2_X1    g643(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT110), .Z(new_n831));
  OR4_X1    g645(.A1(new_n709), .A2(new_n829), .A3(new_n716), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n295), .A2(KEYINPUT85), .A3(new_n300), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT85), .B1(new_n295), .B2(new_n300), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n693), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n817), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n669), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n808), .A2(new_n497), .A3(new_n839), .A4(new_n696), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n838), .A2(new_n841), .B1(new_n774), .B2(new_n775), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n680), .A2(KEYINPUT100), .A3(new_n685), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n687), .B1(new_n635), .B2(new_n684), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n757), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT103), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n693), .A2(new_n756), .A3(new_n757), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT111), .B1(new_n848), .B2(new_n766), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n850), .B(new_n765), .C1(new_n846), .C2(new_n847), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n842), .B(new_n771), .C1(new_n849), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n457), .A2(new_n497), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n853), .B(new_n503), .C1(new_n457), .C2(new_n782), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n305), .A2(new_n389), .A3(new_n647), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n690), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n734), .B1(new_n735), .B2(new_n739), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n743), .A2(new_n751), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n858), .A2(new_n860), .A3(new_n642), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n680), .A2(new_n685), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n762), .A2(new_n696), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n750), .A2(new_n716), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n729), .A2(new_n759), .A3(new_n702), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n871), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(KEYINPUT112), .A3(new_n871), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n833), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n863), .A2(new_n869), .A3(new_n871), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n751), .B(new_n743), .C1(new_n506), .C2(new_n641), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n857), .A3(new_n859), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n755), .A2(new_n758), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n850), .B1(new_n881), .B2(new_n765), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n848), .A2(KEYINPUT111), .A3(new_n766), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n880), .A2(new_n771), .A3(new_n884), .A4(new_n842), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n764), .A2(new_n649), .A3(new_n733), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n846), .B2(new_n847), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n700), .B1(new_n843), .B2(new_n844), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n817), .A2(new_n836), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(new_n868), .A3(new_n729), .A4(new_n866), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n867), .A2(KEYINPUT52), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT53), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT54), .B1(new_n878), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n784), .A2(new_n499), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n808), .A2(new_n733), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n767), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT48), .ZN(new_n900));
  NOR4_X1   g714(.A1(new_n897), .A2(new_n639), .A3(new_n694), .A4(new_n716), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n498), .B(G953), .C1(new_n901), .C2(new_n726), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n896), .A2(new_n639), .A3(new_n748), .ZN(new_n903));
  INV_X1    g717(.A(new_n753), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT115), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n903), .A2(KEYINPUT115), .A3(new_n904), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n900), .B(new_n902), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n749), .A2(new_n733), .ZN(new_n908));
  NOR4_X1   g722(.A1(new_n896), .A2(new_n709), .A3(new_n385), .A4(new_n908), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT50), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n898), .A2(new_n848), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n901), .A2(new_n457), .A3(new_n661), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT51), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n903), .A2(new_n808), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n813), .B(new_n814), .C1(new_n300), .C2(new_n826), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n907), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n916), .A2(KEYINPUT114), .A3(new_n917), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT114), .B1(new_n916), .B2(new_n917), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n913), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n877), .A2(new_n895), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(G952), .A2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n832), .B1(new_n925), .B2(new_n926), .ZN(G75));
  AND2_X1   g741(.A1(G210), .A2(G902), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n878), .A2(new_n894), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n346), .A2(new_n361), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n380), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n929), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n272), .A2(G952), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT117), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT116), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n929), .A2(new_n930), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n933), .ZN(new_n941));
  AOI211_X1 g755(.A(KEYINPUT116), .B(new_n934), .C1(new_n929), .C2(new_n930), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT118), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n938), .B(KEYINPUT118), .C1(new_n941), .C2(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(G51));
  XOR2_X1   g761(.A(new_n792), .B(KEYINPUT57), .Z(new_n948));
  AND3_X1   g762(.A1(new_n878), .A2(new_n894), .A3(KEYINPUT54), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n895), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n291), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n878), .A2(new_n894), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(G902), .A3(new_n790), .A4(new_n789), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n936), .B1(new_n951), .B2(new_n953), .ZN(G54));
  NAND4_X1  g768(.A1(new_n952), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n448), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n448), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n936), .ZN(G60));
  NAND2_X1  g772(.A1(new_n655), .A2(new_n656), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n659), .B(KEYINPUT59), .Z(new_n960));
  OAI211_X1 g774(.A(new_n959), .B(new_n960), .C1(new_n949), .C2(new_n895), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n937), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n877), .B2(new_n895), .ZN(new_n963));
  INV_X1    g777(.A(new_n959), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  NAND3_X1  g781(.A1(new_n878), .A2(new_n894), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n638), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n878), .A2(new_n894), .A3(new_n682), .A4(new_n967), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT119), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n937), .B(new_n969), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G66));
  NAND2_X1  g790(.A1(new_n862), .A2(new_n272), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT120), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n501), .B2(new_n355), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n342), .B(new_n345), .C1(G898), .C2(new_n272), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G69));
  AOI21_X1  g796(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n516), .A2(new_n520), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(new_n439), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n801), .A2(new_n803), .A3(new_n808), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n781), .A2(new_n785), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(KEYINPUT44), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n822), .B1(new_n989), .B2(new_n786), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n767), .A2(new_n750), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n801), .A2(new_n803), .A3(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n801), .A2(new_n803), .A3(new_n991), .A4(KEYINPUT124), .ZN(new_n995));
  AND4_X1   g809(.A1(new_n771), .A2(new_n994), .A3(new_n776), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n729), .A2(new_n759), .A3(new_n702), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT121), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n990), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n272), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n272), .A2(G900), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT125), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1000), .A2(KEYINPUT125), .A3(new_n1001), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n986), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n822), .ZN(new_n1007));
  INV_X1    g821(.A(new_n641), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n853), .B1(new_n457), .B2(new_n782), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT123), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n706), .A2(new_n1008), .A3(new_n808), .A4(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1007), .A2(new_n809), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT121), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n997), .B(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1014), .A2(new_n723), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT62), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT122), .ZN(new_n1018));
  INV_X1    g832(.A(new_n723), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n998), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1018), .B1(new_n1020), .B2(KEYINPUT62), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1015), .A2(KEYINPUT122), .A3(new_n1016), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1017), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n986), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1023), .A2(new_n578), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n984), .B1(new_n1006), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1005), .ZN(new_n1027));
  AOI21_X1  g841(.A(KEYINPUT125), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1024), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1017), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1024), .A2(new_n578), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1029), .A2(new_n1034), .A3(new_n983), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1026), .A2(new_n1035), .ZN(G72));
  NAND2_X1  g850(.A1(new_n874), .A2(new_n873), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n1037), .B(new_n876), .C1(new_n871), .C2(new_n870), .ZN(new_n1038));
  INV_X1    g852(.A(new_n548), .ZN(new_n1039));
  XNOR2_X1  g853(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n546), .A2(new_n292), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1040), .B(new_n1041), .Z(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1039), .A2(new_n710), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1042), .B1(new_n999), .B2(new_n862), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n936), .B1(new_n1046), .B2(new_n1039), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(KEYINPUT127), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1043), .B1(new_n1023), .B2(new_n880), .ZN(new_n1050));
  INV_X1    g864(.A(new_n710), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1042), .B1(new_n1032), .B2(new_n862), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1053), .A2(KEYINPUT127), .A3(new_n710), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1048), .B1(new_n1052), .B2(new_n1054), .ZN(G57));
endmodule


