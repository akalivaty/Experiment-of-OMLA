//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1042, new_n1043;
  AND2_X1   g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT27), .B(G183gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT28), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT26), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n213), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n218), .B1(new_n221), .B2(KEYINPUT24), .ZN(new_n227));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n227), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n226), .A2(KEYINPUT25), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n223), .A3(new_n225), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(KEYINPUT23), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n230), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n221), .A2(KEYINPUT24), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n218), .B(new_n238), .C1(new_n239), .C2(new_n228), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n234), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n233), .A2(KEYINPUT65), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT65), .B1(new_n233), .B2(new_n241), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n222), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G134gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G127gat), .ZN(new_n246));
  INV_X1    g045(.A(G127gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G134gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(KEYINPUT1), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(G120gat), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G113gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n259), .B1(new_n258), .B2(new_n261), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n251), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n265), .B(new_n222), .C1(new_n242), .C2(new_n243), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n202), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n269), .B(KEYINPUT34), .Z(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n202), .A3(new_n268), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n271), .A2(KEYINPUT32), .ZN(new_n272));
  XOR2_X1   g071(.A(G15gat), .B(G43gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT69), .ZN(new_n274));
  XNOR2_X1  g073(.A(G71gat), .B(G99gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT33), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n276), .B1(new_n271), .B2(KEYINPUT32), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT33), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n271), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n272), .A2(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n270), .B1(new_n283), .B2(KEYINPUT71), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n282), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n271), .A2(new_n279), .A3(KEYINPUT32), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT71), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT72), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n286), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n292), .A2(new_n293), .A3(new_n287), .A4(new_n270), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n290), .A2(new_n270), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT77), .ZN(new_n296));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT22), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n302), .B(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306));
  AND2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308));
  INV_X1    g107(.A(G155gat), .ZN(new_n309));
  INV_X1    g108(.A(G162gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  AOI211_X1 g111(.A(new_n306), .B(new_n307), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT76), .B1(new_n307), .B2(new_n306), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  INV_X1    g114(.A(G148gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n318));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n312), .A2(KEYINPUT2), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n314), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n324), .B(new_n325), .C1(G155gat), .C2(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n313), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n305), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n302), .A2(new_n304), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n303), .B1(new_n301), .B2(new_n297), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n328), .B1(new_n335), .B2(new_n329), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n296), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(G228gat), .A3(G233gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n296), .B(new_n339), .C1(new_n332), .C2(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G22gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT31), .B(G50gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT78), .B(G22gat), .Z(new_n347));
  NAND3_X1  g146(.A1(new_n338), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n348), .ZN(new_n350));
  INV_X1    g149(.A(new_n347), .ZN(new_n351));
  INV_X1    g150(.A(new_n340), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT3), .B1(new_n305), .B2(new_n331), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n328), .B2(new_n329), .ZN(new_n354));
  OAI22_X1  g153(.A1(new_n328), .A2(new_n353), .B1(new_n354), .B2(new_n305), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n339), .B1(new_n355), .B2(new_n296), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n351), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n359), .A3(new_n351), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n350), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n349), .B1(new_n361), .B2(new_n346), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n289), .A2(new_n294), .A3(new_n295), .A4(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n305), .ZN(new_n364));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n365), .B(KEYINPUT73), .Z(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(new_n244), .B2(new_n331), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n210), .B2(new_n212), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n369), .B1(new_n241), .B2(new_n233), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(new_n365), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n364), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n365), .B1(new_n370), .B2(KEYINPUT29), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT65), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT25), .B1(new_n226), .B2(new_n232), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n237), .A2(new_n240), .A3(new_n234), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n233), .A2(new_n241), .A3(KEYINPUT65), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n369), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n366), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n373), .B(new_n305), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n372), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(G8gat), .B(G36gat), .Z(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT74), .ZN(new_n384));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OR3_X1    g186(.A1(new_n382), .A2(KEYINPUT30), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n380), .B1(new_n379), .B2(KEYINPUT29), .ZN(new_n389));
  INV_X1    g188(.A(new_n371), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n305), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n381), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n372), .A2(new_n381), .A3(new_n386), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT30), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n322), .A2(new_n327), .ZN(new_n399));
  INV_X1    g198(.A(new_n313), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n265), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n264), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n262), .A3(new_n255), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n328), .B1(new_n404), .B2(new_n251), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n398), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT5), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n307), .A2(new_n306), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n408), .A2(new_n318), .B1(KEYINPUT2), .B2(new_n312), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n326), .B1(new_n409), .B2(new_n314), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(new_n410), .B2(new_n313), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(new_n330), .A3(new_n265), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n265), .B2(new_n401), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n404), .A2(new_n328), .A3(KEYINPUT4), .A4(new_n251), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n412), .A2(new_n414), .A3(new_n397), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT5), .A3(new_n397), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT0), .ZN(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n425), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n418), .A2(new_n397), .B1(KEYINPUT5), .B2(new_n406), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n416), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n419), .A3(new_n425), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n396), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT35), .B1(new_n363), .B2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT82), .B(KEYINPUT35), .Z(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n388), .B2(new_n395), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n290), .A2(new_n270), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n362), .A2(new_n439), .A3(new_n295), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n425), .B(KEYINPUT80), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n417), .A2(new_n419), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n431), .A2(new_n432), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n431), .A2(KEYINPUT81), .A3(new_n432), .A4(new_n444), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n426), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n441), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n295), .A2(new_n440), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT36), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n289), .A2(new_n294), .A3(new_n295), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(KEYINPUT36), .ZN(new_n456));
  INV_X1    g255(.A(new_n349), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n358), .A2(new_n360), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n348), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n459), .B2(new_n345), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n436), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n375), .A2(new_n376), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n331), .B1(new_n463), .B2(new_n369), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n244), .A2(new_n366), .B1(new_n464), .B2(new_n365), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n462), .B1(new_n465), .B2(new_n364), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n305), .B1(new_n367), .B2(new_n371), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT38), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n386), .B1(new_n372), .B2(new_n381), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n386), .A2(new_n462), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n470), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n393), .A2(new_n472), .B1(new_n382), .B2(KEYINPUT37), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT38), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n394), .B(new_n471), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n449), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n398), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n478), .A2(KEYINPUT39), .ZN(new_n479));
  OR3_X1    g278(.A1(new_n402), .A2(new_n405), .A3(new_n398), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(KEYINPUT39), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n442), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n482), .A2(new_n483), .B1(new_n421), .B2(new_n443), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n479), .A2(KEYINPUT40), .A3(new_n442), .A4(new_n481), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n484), .A2(new_n388), .A3(new_n395), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n362), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n461), .B1(new_n476), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n437), .A2(new_n452), .B1(new_n456), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491));
  INV_X1    g290(.A(G50gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G43gat), .ZN(new_n493));
  INV_X1    g292(.A(G43gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G50gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT83), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n493), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(KEYINPUT15), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G29gat), .ZN(new_n501));
  INV_X1    g300(.A(G36gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT14), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(G29gat), .B2(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n492), .A2(KEYINPUT86), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G50gat), .ZN(new_n511));
  AOI21_X1  g310(.A(G43gat), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n493), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n500), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT84), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT84), .ZN(new_n518));
  NAND2_X1  g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n499), .A2(KEYINPUT15), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n498), .B1(new_n493), .B2(new_n495), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n520), .B2(new_n523), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n515), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT16), .ZN(new_n529));
  INV_X1    g328(.A(G22gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G15gat), .ZN(new_n531));
  INV_X1    g330(.A(G15gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n531), .B2(new_n533), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n531), .A2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n528), .A3(new_n535), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT88), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n538), .B(new_n541), .C1(new_n542), .C2(G8gat), .ZN(new_n543));
  AOI21_X1  g342(.A(G8gat), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n543), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n500), .A2(new_n507), .A3(new_n514), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n518), .A2(new_n519), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT84), .B1(new_n503), .B2(new_n505), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT85), .B1(new_n552), .B2(new_n500), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n548), .B1(new_n555), .B2(KEYINPUT17), .ZN(new_n556));
  OAI211_X1 g355(.A(KEYINPUT17), .B(new_n515), .C1(new_n525), .C2(new_n526), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n491), .B(new_n547), .C1(new_n556), .C2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT89), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n555), .A2(new_n548), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n527), .A2(new_n563), .B1(new_n543), .B2(new_n546), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n564), .B2(new_n557), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT18), .A4(new_n491), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n555), .A2(new_n548), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n547), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n491), .B(KEYINPUT13), .Z(new_n571));
  AOI22_X1  g370(.A1(new_n559), .A2(new_n560), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G197gat), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT11), .B(G169gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT12), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n568), .A2(new_n580), .A3(new_n572), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n490), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  XOR2_X1   g384(.A(G99gat), .B(G106gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT8), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(G99gat), .B2(G106gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT99), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT8), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n587), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  AOI211_X1 g405(.A(new_n586), .B(new_n604), .C1(new_n591), .C2(new_n598), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT100), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(G64gat), .ZN(new_n612));
  OR3_X1    g411(.A1(new_n612), .A2(KEYINPUT90), .A3(G57gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(G57gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT90), .B1(new_n612), .B2(G57gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(G71gat), .A2(G78gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(G71gat), .A2(G78gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT91), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT91), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n621), .A3(new_n618), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n611), .A2(new_n616), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G57gat), .B(G64gat), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n618), .B(new_n617), .C1(new_n624), .C2(new_n609), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n594), .B1(new_n593), .B2(new_n597), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n605), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n586), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n599), .A2(new_n587), .A3(new_n605), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n608), .A2(new_n626), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n631), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n635), .A2(KEYINPUT100), .A3(new_n625), .A4(new_n623), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT10), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n623), .A2(KEYINPUT94), .A3(new_n625), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT94), .B1(new_n623), .B2(new_n625), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NOR4_X1   g440(.A1(new_n639), .A2(new_n635), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n585), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n585), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n634), .A2(new_n644), .A3(new_n636), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n643), .A2(new_n645), .A3(new_n649), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(KEYINPUT101), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n654), .A3(new_n650), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n640), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT21), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n548), .ZN(new_n659));
  XNOR2_X1  g458(.A(G127gat), .B(G155gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(G231gat), .A2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n659), .B(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT21), .B1(new_n623), .B2(new_n625), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT93), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(G183gat), .B(G211gat), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n668), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n664), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n671), .A3(new_n663), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G134gat), .B(G162gat), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n685));
  AND3_X1   g484(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n686));
  INV_X1    g485(.A(new_n635), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n527), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n635), .B1(new_n555), .B2(KEYINPUT17), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(new_n558), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G190gat), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n688), .B(new_n207), .C1(new_n689), .C2(new_n558), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n685), .B1(new_n693), .B2(new_n300), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n691), .A2(G218gat), .A3(new_n692), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n684), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n692), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n527), .A2(new_n563), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n557), .A3(new_n635), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n207), .B1(new_n699), .B2(new_n688), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n300), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  AND4_X1   g500(.A1(KEYINPUT97), .A2(new_n701), .A3(new_n695), .A4(new_n684), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n682), .B1(new_n696), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(KEYINPUT97), .A3(new_n695), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n683), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n694), .A2(new_n695), .A3(new_n684), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n706), .A3(new_n681), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n656), .B(new_n678), .C1(new_n703), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n584), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n435), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n528), .ZN(G1324gat));
  NOR2_X1   g510(.A1(new_n709), .A2(new_n396), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT16), .B(G8gat), .Z(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G8gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  MUX2_X1   g515(.A(new_n714), .B(new_n716), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g516(.A(G15gat), .B1(new_n709), .B2(new_n456), .ZN(new_n718));
  INV_X1    g517(.A(new_n453), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n532), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n709), .B2(new_n720), .ZN(G1326gat));
  NOR2_X1   g520(.A1(new_n709), .A2(new_n362), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT43), .B(G22gat), .Z(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  NAND2_X1  g523(.A1(new_n703), .A2(new_n707), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(new_n677), .A3(new_n656), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n584), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(G29gat), .A3(new_n435), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT45), .Z(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n490), .B2(new_n725), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n437), .A2(new_n452), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n456), .A2(new_n489), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n696), .A2(new_n702), .A3(new_n682), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n681), .B1(new_n705), .B2(new_n706), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(KEYINPUT44), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n568), .A2(new_n580), .A3(new_n572), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n580), .B1(new_n568), .B2(new_n572), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n579), .A2(KEYINPUT102), .A3(new_n581), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n656), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n678), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT103), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n739), .A2(KEYINPUT104), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n435), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n731), .A2(new_n738), .ZN(new_n753));
  INV_X1    g552(.A(new_n749), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n750), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n729), .B1(new_n501), .B2(new_n756), .ZN(G1328gat));
  NOR3_X1   g556(.A1(new_n727), .A2(G36gat), .A3(new_n396), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT46), .ZN(new_n759));
  INV_X1    g558(.A(new_n396), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n750), .A2(new_n760), .A3(new_n755), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n761), .B2(new_n502), .ZN(G1329gat));
  NOR3_X1   g561(.A1(new_n727), .A2(G43gat), .A3(new_n453), .ZN(new_n763));
  INV_X1    g562(.A(new_n456), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n750), .A2(new_n764), .A3(new_n755), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n763), .B1(new_n765), .B2(G43gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n753), .A2(new_n754), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n494), .B1(new_n767), .B2(new_n764), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n766), .A2(KEYINPUT47), .B1(new_n768), .B2(new_n770), .ZN(G1330gat));
  NAND2_X1  g570(.A1(new_n509), .A2(new_n511), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n362), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n727), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT105), .B1(new_n584), .B2(new_n726), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n750), .A2(new_n460), .A3(new_n755), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n772), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT48), .B1(new_n775), .B2(new_n776), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n767), .A2(new_n460), .B1(new_n509), .B2(new_n511), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n779), .A2(KEYINPUT48), .B1(new_n780), .B2(new_n781), .ZN(G1331gat));
  NAND2_X1  g581(.A1(new_n725), .A2(new_n677), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n490), .A2(new_n783), .A3(new_n747), .A4(new_n746), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n751), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n760), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT49), .B(G64gat), .Z(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(G1333gat));
  NAND2_X1  g589(.A1(new_n784), .A2(new_n764), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n453), .A2(G71gat), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n791), .A2(G71gat), .B1(new_n784), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n784), .A2(new_n460), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT107), .B(G78gat), .Z(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1335gat));
  NAND2_X1  g597(.A1(new_n751), .A2(new_n595), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT36), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n290), .A2(new_n270), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n292), .A2(new_n287), .A3(new_n270), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(KEYINPUT72), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n802), .B1(new_n805), .B2(new_n294), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n806), .A2(new_n488), .A3(new_n454), .ZN(new_n807));
  INV_X1    g606(.A(new_n436), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n805), .A2(new_n808), .A3(new_n294), .A4(new_n362), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n451), .B1(new_n809), .B2(KEYINPUT35), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n801), .B(new_n737), .C1(new_n807), .C2(new_n810), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n746), .A2(KEYINPUT108), .A3(new_n677), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT108), .B1(new_n746), .B2(new_n677), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n801), .B1(new_n734), .B2(new_n737), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n800), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT110), .B1(new_n490), .B2(new_n725), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(KEYINPUT51), .A3(new_n814), .A4(new_n811), .ZN(new_n819));
  AOI211_X1 g618(.A(new_n747), .B(new_n799), .C1(new_n817), .C2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n747), .B1(new_n812), .B2(new_n813), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n731), .A2(new_n738), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(KEYINPUT109), .A3(new_n751), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n731), .A2(new_n738), .A3(new_n751), .A4(new_n822), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT109), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n595), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n821), .A2(KEYINPUT111), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n824), .A2(new_n827), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n820), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1336gat));
  AOI21_X1  g632(.A(new_n596), .B1(new_n823), .B2(new_n760), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n747), .B1(new_n817), .B2(new_n819), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n396), .A2(G92gat), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n836), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n747), .B(new_n840), .C1(new_n817), .C2(new_n819), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT52), .B1(new_n841), .B2(new_n834), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(G1337gat));
  AOI21_X1  g642(.A(G99gat), .B1(new_n835), .B2(new_n719), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n764), .A2(G99gat), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n823), .B2(new_n845), .ZN(G1338gat));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  AOI21_X1  g646(.A(G106gat), .B1(new_n835), .B2(new_n460), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n823), .A2(G106gat), .A3(new_n460), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g650(.A(new_n362), .B(new_n747), .C1(new_n817), .C2(new_n819), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n849), .B(KEYINPUT53), .C1(new_n852), .C2(G106gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1339gat));
  NOR2_X1   g653(.A1(new_n565), .A2(new_n491), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n570), .A2(new_n571), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n577), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n581), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n656), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n581), .A2(new_n653), .A3(new_n655), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT112), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n634), .A2(new_n636), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n641), .ZN(new_n866));
  INV_X1    g665(.A(new_n642), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n644), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n868), .A2(KEYINPUT54), .A3(new_n643), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n585), .C1(new_n637), .C2(new_n642), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n650), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n864), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n872), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n868), .A2(KEYINPUT54), .A3(new_n643), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(KEYINPUT55), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n873), .A2(new_n652), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n743), .A2(new_n744), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n737), .B1(new_n863), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n652), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n581), .A2(new_n857), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(new_n703), .A3(new_n707), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n678), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n708), .A2(new_n745), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n460), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(new_n751), .A3(new_n396), .A4(new_n719), .ZN(new_n887));
  OAI21_X1  g686(.A(G113gat), .B1(new_n887), .B2(new_n583), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n878), .A2(new_n862), .A3(new_n860), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n883), .B1(new_n889), .B2(new_n725), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n885), .B1(new_n890), .B2(new_n677), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(new_n435), .A3(new_n363), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(new_n396), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT113), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n746), .A2(new_n256), .A3(new_n257), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(G1340gat));
  OAI21_X1  g696(.A(G120gat), .B1(new_n887), .B2(new_n747), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n656), .A2(new_n260), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n895), .B2(new_n899), .ZN(G1341gat));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n247), .A3(new_n677), .ZN(new_n901));
  OAI21_X1  g700(.A(G127gat), .B1(new_n887), .B2(new_n678), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(KEYINPUT114), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1342gat));
  NOR2_X1   g706(.A1(new_n725), .A2(new_n760), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n245), .A3(new_n908), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(KEYINPUT56), .ZN(new_n910));
  OAI21_X1  g709(.A(G134gat), .B1(new_n887), .B2(new_n725), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(KEYINPUT56), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G1343gat));
  NOR3_X1   g712(.A1(new_n764), .A2(new_n435), .A3(new_n760), .ZN(new_n914));
  XNOR2_X1  g713(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n891), .B2(new_n460), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n460), .A2(KEYINPUT57), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n882), .A2(new_n703), .A3(new_n707), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n876), .A2(new_n652), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n579), .B2(new_n581), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n869), .B2(new_n872), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n874), .A2(KEYINPUT116), .A3(new_n875), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n864), .A3(new_n924), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n921), .A2(new_n925), .B1(new_n656), .B2(new_n858), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n919), .B1(new_n926), .B2(new_n737), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n678), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n918), .B1(new_n928), .B2(new_n885), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n914), .B1(new_n917), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G141gat), .B1(new_n930), .B2(new_n583), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n764), .A2(new_n362), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n891), .A2(new_n751), .A3(new_n396), .A4(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n583), .A2(G141gat), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n931), .B(new_n932), .C1(new_n934), .C2(new_n936), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n746), .B(new_n914), .C1(new_n917), .C2(new_n929), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(G141gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n938), .B2(G141gat), .ZN(new_n941));
  INV_X1    g740(.A(new_n934), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(new_n935), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT118), .B1(new_n934), .B2(new_n936), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n940), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n937), .B1(new_n947), .B2(new_n932), .ZN(G1344gat));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n316), .A3(new_n656), .ZN(new_n949));
  INV_X1    g748(.A(new_n930), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT59), .B(new_n316), .C1(new_n950), .C2(new_n656), .ZN(new_n951));
  XOR2_X1   g750(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n952));
  INV_X1    g751(.A(KEYINPUT57), .ZN(new_n953));
  AOI22_X1  g752(.A1(new_n927), .A2(new_n678), .B1(new_n583), .B2(new_n708), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n362), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n362), .A2(new_n915), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n743), .A2(new_n744), .A3(new_n877), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n860), .A2(new_n862), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n725), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n677), .B1(new_n959), .B2(new_n919), .ZN(new_n960));
  INV_X1    g759(.A(new_n885), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n955), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n656), .A3(new_n914), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n952), .B1(new_n964), .B2(G148gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n949), .B1(new_n951), .B2(new_n965), .ZN(G1345gat));
  NOR3_X1   g765(.A1(new_n930), .A2(new_n309), .A3(new_n678), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT120), .B1(new_n934), .B2(new_n678), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n934), .A2(KEYINPUT120), .A3(new_n678), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n969), .A2(G155gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n967), .B1(new_n968), .B2(new_n970), .ZN(G1346gat));
  OAI21_X1  g770(.A(G162gat), .B1(new_n930), .B2(new_n725), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n891), .A2(new_n751), .A3(new_n933), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n908), .A2(new_n310), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G1347gat));
  NOR2_X1   g774(.A1(new_n751), .A2(new_n396), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n977), .A2(new_n453), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT122), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n886), .A2(new_n979), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n980), .A2(new_n214), .A3(new_n583), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n892), .A2(new_n751), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n363), .A2(new_n396), .ZN(new_n983));
  XOR2_X1   g782(.A(new_n983), .B(KEYINPUT121), .Z(new_n984));
  AND2_X1   g783(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(new_n746), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n981), .B1(new_n986), .B2(new_n214), .ZN(G1348gat));
  NAND3_X1  g786(.A1(new_n985), .A2(new_n215), .A3(new_n656), .ZN(new_n988));
  OAI21_X1  g787(.A(G176gat), .B1(new_n980), .B2(new_n747), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1349gat));
  AND2_X1   g789(.A1(new_n677), .A2(new_n211), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT123), .ZN(new_n992));
  AOI22_X1  g791(.A1(new_n985), .A2(new_n991), .B1(new_n992), .B2(KEYINPUT60), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n992), .A2(KEYINPUT60), .ZN(new_n994));
  OAI21_X1  g793(.A(G183gat), .B1(new_n980), .B2(new_n678), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n994), .B1(new_n993), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n996), .A2(new_n997), .ZN(G1350gat));
  NAND3_X1  g797(.A1(new_n985), .A2(new_n207), .A3(new_n737), .ZN(new_n999));
  OAI21_X1  g798(.A(G190gat), .B1(new_n980), .B2(new_n725), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(KEYINPUT124), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n1003), .B(G190gat), .C1(new_n980), .C2(new_n725), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1002), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n999), .B1(new_n1005), .B2(new_n1006), .ZN(G1351gat));
  NOR3_X1   g806(.A1(new_n764), .A2(new_n396), .A3(new_n362), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n982), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(G197gat), .B1(new_n1010), .B2(new_n746), .ZN(new_n1011));
  AND3_X1   g810(.A1(new_n456), .A2(KEYINPUT125), .A3(new_n976), .ZN(new_n1012));
  AOI21_X1  g811(.A(KEYINPUT125), .B1(new_n456), .B2(new_n976), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1014), .B1(new_n955), .B2(new_n962), .ZN(new_n1015));
  AND2_X1   g814(.A1(new_n582), .A2(G197gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(G1352gat));
  NOR3_X1   g816(.A1(new_n1009), .A2(G204gat), .A3(new_n747), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT62), .ZN(new_n1019));
  INV_X1    g818(.A(new_n1015), .ZN(new_n1020));
  OAI21_X1  g819(.A(G204gat), .B1(new_n1020), .B2(new_n747), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1019), .A2(new_n1021), .ZN(G1353gat));
  NAND3_X1  g821(.A1(new_n1010), .A2(new_n299), .A3(new_n677), .ZN(new_n1023));
  INV_X1    g822(.A(new_n1014), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n708), .A2(new_n583), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n928), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g825(.A(KEYINPUT57), .B1(new_n1026), .B2(new_n460), .ZN(new_n1027));
  INV_X1    g826(.A(new_n956), .ZN(new_n1028));
  AOI21_X1  g827(.A(new_n1028), .B1(new_n884), .B2(new_n885), .ZN(new_n1029));
  OAI211_X1 g828(.A(new_n1024), .B(new_n677), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1015), .A2(KEYINPUT126), .A3(new_n677), .ZN(new_n1033));
  OR2_X1    g832(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n1034));
  NAND4_X1  g833(.A1(new_n1032), .A2(G211gat), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g834(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g836(.A(new_n678), .B(new_n1014), .C1(new_n955), .C2(new_n962), .ZN(new_n1038));
  AOI21_X1  g837(.A(new_n299), .B1(new_n1038), .B2(KEYINPUT126), .ZN(new_n1039));
  AOI21_X1  g838(.A(new_n1034), .B1(new_n1039), .B2(new_n1032), .ZN(new_n1040));
  OAI21_X1  g839(.A(new_n1023), .B1(new_n1037), .B2(new_n1040), .ZN(G1354gat));
  NAND3_X1  g840(.A1(new_n1010), .A2(new_n300), .A3(new_n737), .ZN(new_n1042));
  OAI21_X1  g841(.A(G218gat), .B1(new_n1020), .B2(new_n725), .ZN(new_n1043));
  NAND2_X1  g842(.A1(new_n1042), .A2(new_n1043), .ZN(G1355gat));
endmodule


