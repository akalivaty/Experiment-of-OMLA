//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G137), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n190), .B(KEYINPUT11), .C1(new_n188), .C2(G137), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G134), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT11), .B1(new_n194), .B2(new_n190), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n189), .B1(new_n192), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n190), .B1(new_n188), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n191), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n193), .B2(G134), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT65), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  AOI211_X1 g020(.A(new_n206), .B(new_n203), .C1(new_n200), .C2(new_n191), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n197), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT0), .A3(G128), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT0), .B(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n202), .B1(new_n194), .B2(new_n189), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT66), .A2(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT66), .A2(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(G143), .B2(new_n216), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n209), .A2(new_n224), .A3(G128), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n215), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n205), .B2(new_n207), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n214), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G119), .ZN(new_n233));
  INV_X1    g047(.A(G119), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT68), .A3(G116), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT2), .B(G113), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n230), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n214), .A2(new_n241), .A3(new_n229), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n245));
  OR3_X1    g059(.A1(new_n244), .A2(KEYINPUT75), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n244), .A2(new_n245), .ZN(new_n247));
  INV_X1    g061(.A(new_n242), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(KEYINPUT28), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT75), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n246), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT69), .B(G237), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT27), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n258), .A3(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n257), .B2(new_n259), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(G902), .B1(new_n252), .B2(new_n266), .ZN(new_n267));
  AOI22_X1  g081(.A1(KEYINPUT67), .A2(new_n229), .B1(new_n208), .B2(new_n213), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n269), .B(new_n228), .C1(new_n205), .C2(new_n207), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n241), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n248), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n214), .A2(new_n274), .A3(new_n270), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n275), .B2(new_n239), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n249), .B1(new_n278), .B2(KEYINPUT28), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n263), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n214), .A2(KEYINPUT30), .A3(new_n229), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n239), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n242), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n264), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n280), .A2(new_n265), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n187), .B1(new_n267), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n245), .B1(new_n273), .B2(new_n277), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n292), .B(new_n264), .C1(new_n293), .C2(new_n249), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT31), .ZN(new_n295));
  INV_X1    g109(.A(new_n284), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n242), .A2(new_n263), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT70), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n242), .A2(new_n263), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n295), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n284), .A2(KEYINPUT31), .A3(new_n300), .A4(new_n298), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n294), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n275), .A2(new_n272), .A3(new_n239), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n242), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT28), .B1(new_n307), .B2(new_n276), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n263), .B1(new_n308), .B2(new_n250), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(new_n292), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n291), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT72), .B1(new_n279), .B2(new_n263), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n312), .A2(KEYINPUT73), .A3(new_n304), .A4(new_n294), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(G472), .A2(G902), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT74), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n290), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  AOI211_X1 g132(.A(KEYINPUT32), .B(new_n316), .C1(new_n311), .C2(new_n313), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n289), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G214), .B1(G237), .B2(G902), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT87), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G210), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n226), .A2(new_n227), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT77), .B(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n327), .B2(new_n212), .ZN(new_n329));
  INV_X1    g143(.A(G224), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT7), .B1(new_n330), .B2(G953), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G104), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT82), .B1(new_n333), .B2(G107), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n335));
  INV_X1    g149(.A(G107), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(G104), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(G107), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G101), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(KEYINPUT83), .A3(G101), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n237), .A2(new_n238), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT5), .A4(new_n236), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n232), .A2(KEYINPUT5), .A3(G119), .ZN(new_n347));
  INV_X1    g161(.A(G113), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n345), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT3), .B1(new_n333), .B2(G107), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n336), .A3(G104), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n351), .A2(new_n353), .A3(new_n354), .A4(new_n338), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G122), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n353), .A3(new_n338), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT80), .A4(new_n338), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(G101), .A3(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n362), .A2(new_n366), .A3(G101), .A4(new_n363), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n239), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n358), .B(new_n359), .C1(new_n365), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n355), .A2(new_n356), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n355), .A2(new_n356), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n370), .A2(new_n371), .B1(new_n342), .B2(new_n343), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(new_n350), .ZN(new_n373));
  INV_X1    g187(.A(new_n358), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n359), .B(KEYINPUT8), .Z(new_n376));
  OAI211_X1 g190(.A(new_n332), .B(new_n369), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n366), .B1(new_n371), .B2(new_n370), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n368), .B1(new_n364), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n382), .B2(new_n374), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n384));
  OAI211_X1 g198(.A(KEYINPUT88), .B(new_n358), .C1(new_n365), .C2(new_n368), .ZN(new_n385));
  INV_X1    g199(.A(new_n359), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT89), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n358), .B1(new_n365), .B2(new_n368), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n359), .B1(new_n389), .B2(new_n380), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n384), .A4(new_n385), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n385), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n369), .A2(KEYINPUT6), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n388), .A2(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n330), .A2(G953), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n329), .B(new_n396), .Z(new_n397));
  AOI211_X1 g211(.A(new_n325), .B(new_n379), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n388), .A2(new_n392), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n394), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n379), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n324), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n323), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT90), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n407));
  INV_X1    g221(.A(G469), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n213), .A3(new_n367), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n372), .A2(KEYINPUT10), .A3(new_n326), .ZN(new_n411));
  INV_X1    g225(.A(G128), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n220), .B1(new_n225), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n227), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n344), .A2(new_n357), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT10), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n201), .A2(new_n204), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n206), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n201), .A2(KEYINPUT65), .A3(new_n204), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n419), .A2(new_n420), .B1(G131), .B2(new_n196), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n410), .A2(new_n411), .A3(new_n417), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n254), .A2(G227), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n422), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n429));
  NAND2_X1  g243(.A1(new_n344), .A2(new_n357), .ZN(new_n430));
  INV_X1    g244(.A(new_n326), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n415), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n429), .B1(new_n433), .B2(new_n208), .ZN(new_n434));
  NOR2_X1   g248(.A1(KEYINPUT84), .A2(KEYINPUT12), .ZN(new_n435));
  AOI211_X1 g249(.A(new_n435), .B(new_n421), .C1(new_n432), .C2(new_n415), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n423), .B1(new_n422), .B2(new_n427), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n428), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n410), .A2(new_n411), .A3(new_n417), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n208), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n427), .B1(new_n441), .B2(new_n422), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n408), .B(new_n378), .C1(new_n439), .C2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n408), .A2(new_n378), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n422), .B1(new_n434), .B2(new_n436), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n422), .A2(new_n427), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n445), .A2(new_n426), .B1(new_n446), .B2(new_n441), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n447), .B2(G469), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT9), .B(G234), .ZN(new_n450));
  OAI21_X1  g264(.A(G221), .B1(new_n450), .B2(G902), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n407), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n451), .ZN(new_n453));
  AOI211_X1 g267(.A(KEYINPUT86), .B(new_n453), .C1(new_n443), .C2(new_n448), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT90), .B(new_n323), .C1(new_n398), .C2(new_n403), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n232), .A2(G122), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n336), .B1(new_n457), .B2(KEYINPUT14), .ZN(new_n458));
  XOR2_X1   g272(.A(G116), .B(G122), .Z(new_n459));
  XOR2_X1   g273(.A(new_n458), .B(new_n459), .Z(new_n460));
  NAND2_X1  g274(.A1(new_n218), .A2(G128), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT66), .B(G128), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n218), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(G134), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n461), .B(KEYINPUT13), .Z(new_n466));
  NOR2_X1   g280(.A1(new_n462), .A2(new_n218), .ZN(new_n467));
  OAI21_X1  g281(.A(G134), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n459), .B(G107), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(new_n469), .C1(G134), .C2(new_n463), .ZN(new_n470));
  INV_X1    g284(.A(G217), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n450), .A2(new_n471), .A3(G953), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n465), .B2(new_n470), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OR3_X1    g290(.A1(new_n476), .A2(KEYINPUT93), .A3(G902), .ZN(new_n477));
  INV_X1    g291(.A(G478), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT15), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n477), .B(new_n479), .Z(new_n480));
  NAND3_X1  g294(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n253), .A2(G214), .A3(new_n254), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n218), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT17), .A3(G131), .ZN(new_n485));
  INV_X1    g299(.A(G125), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(G140), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n327), .B2(G140), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT16), .ZN(new_n489));
  OR3_X1    g303(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n490));
  AOI21_X1  g304(.A(G146), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(G146), .A3(new_n490), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n485), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT91), .B1(new_n484), .B2(G131), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n484), .A2(G131), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n481), .A2(new_n498), .A3(new_n202), .A4(new_n483), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(G113), .B(G122), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(new_n333), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT18), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n202), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n484), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n484), .A2(new_n505), .ZN(new_n507));
  INV_X1    g321(.A(new_n487), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n486), .A2(G140), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n216), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n488), .B2(new_n216), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n501), .A2(new_n503), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n503), .B1(new_n501), .B2(new_n512), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n378), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT92), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n517), .B(new_n378), .C1(new_n513), .C2(new_n514), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(G475), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n521));
  INV_X1    g335(.A(new_n493), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n508), .A2(new_n509), .ZN(new_n523));
  MUX2_X1   g337(.A(new_n523), .B(new_n488), .S(KEYINPUT19), .Z(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n216), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n503), .B1(new_n526), .B2(new_n512), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n520), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT20), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT20), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n530), .B(new_n520), .C1(new_n513), .C2(new_n527), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n480), .A2(new_n519), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n254), .A2(G952), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(G234), .B2(G237), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT21), .B(G898), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT94), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI211_X1 g352(.A(new_n378), .B(new_n254), .C1(G234), .C2(G237), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  AND4_X1   g355(.A1(new_n406), .A2(new_n455), .A3(new_n456), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n471), .B1(G234), .B2(new_n378), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT22), .B(G137), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n462), .A2(new_n234), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n412), .A2(G119), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT76), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n223), .A2(G119), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT76), .ZN(new_n552));
  INV_X1    g366(.A(new_n549), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT24), .B(G110), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n234), .B2(G128), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n553), .B(new_n559), .C1(new_n551), .C2(new_n558), .ZN(new_n560));
  OAI22_X1  g374(.A1(new_n555), .A2(new_n557), .B1(G110), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n493), .A3(new_n510), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n557), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(G110), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n563), .B(new_n564), .C1(new_n522), .C2(new_n491), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT78), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT78), .B1(new_n562), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n547), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n546), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT25), .B1(new_n571), .B2(new_n378), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT25), .ZN(new_n573));
  AOI211_X1 g387(.A(new_n573), .B(G902), .C1(new_n568), .C2(new_n570), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n543), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n543), .A2(G902), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT79), .ZN(new_n577));
  INV_X1    g391(.A(new_n571), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n320), .A2(new_n542), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  NOR3_X1   g396(.A1(new_n305), .A2(new_n310), .A3(new_n291), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n309), .A2(new_n292), .B1(new_n302), .B2(new_n303), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT73), .B1(new_n584), .B2(new_n312), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n317), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n452), .A2(new_n454), .A3(new_n579), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n378), .B1(new_n583), .B2(new_n585), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n589));
  OAI21_X1  g403(.A(G472), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n311), .B2(new_n313), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT95), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n586), .B(new_n587), .C1(new_n590), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n519), .A2(new_n532), .ZN(new_n594));
  NAND2_X1  g408(.A1(G478), .A2(G902), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n378), .B1(new_n474), .B2(new_n475), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(G478), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n476), .B(KEYINPUT33), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(G478), .ZN(new_n599));
  INV_X1    g413(.A(new_n540), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n594), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n593), .A2(new_n404), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT96), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT34), .B(G104), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G6));
  NOR2_X1   g420(.A1(new_n594), .A2(new_n480), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n600), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n593), .A2(new_n404), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT35), .B(G107), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  AOI21_X1  g425(.A(new_n316), .B1(new_n311), .B2(new_n313), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n187), .B1(new_n591), .B2(KEYINPUT95), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n588), .A2(new_n589), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n455), .A2(new_n406), .A3(new_n456), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n566), .A2(new_n567), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT97), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n617), .B(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n577), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n575), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n541), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT37), .B(G110), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT98), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G12));
  OAI211_X1 g443(.A(new_n623), .B(new_n323), .C1(new_n403), .C2(new_n398), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n535), .B(KEYINPUT99), .Z(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n539), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n594), .A2(new_n480), .A3(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n631), .A2(new_n455), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n320), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  INV_X1    g453(.A(new_n480), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n594), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n623), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n323), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT102), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n635), .B(KEYINPUT39), .ZN(new_n646));
  OR3_X1    g460(.A1(new_n452), .A2(new_n454), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(KEYINPUT40), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(KEYINPUT40), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n398), .A2(new_n403), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT38), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n645), .A2(new_n648), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  OAI22_X1  g466(.A1(new_n296), .A2(new_n301), .B1(new_n263), .B2(new_n244), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n187), .B1(new_n653), .B2(new_n378), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n318), .B2(new_n319), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT100), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n586), .A2(KEYINPUT32), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n612), .A2(new_n290), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n661), .A3(new_n655), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n657), .A2(new_n662), .A3(KEYINPUT101), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n661), .B1(new_n660), .B2(new_n655), .ZN(new_n665));
  AOI211_X1 g479(.A(KEYINPUT100), .B(new_n654), .C1(new_n658), .C2(new_n659), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n652), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT103), .B(G143), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G45));
  INV_X1    g484(.A(new_n635), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n594), .A2(new_n599), .A3(new_n671), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n630), .A2(new_n452), .A3(new_n672), .A4(new_n454), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n320), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT104), .B(G146), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G48));
  NOR2_X1   g490(.A1(new_n439), .A2(new_n442), .ZN(new_n677));
  OAI21_X1  g491(.A(G469), .B1(new_n677), .B2(G902), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n451), .A3(new_n443), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n602), .A2(new_n404), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n320), .A2(new_n580), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT105), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G15));
  NOR3_X1   g498(.A1(new_n608), .A2(new_n404), .A3(new_n679), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n320), .A2(new_n580), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  NOR3_X1   g501(.A1(new_n624), .A2(new_n404), .A3(new_n679), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n320), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  NOR4_X1   g504(.A1(new_n404), .A2(new_n641), .A3(new_n679), .A4(new_n540), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n263), .B1(new_n252), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n692), .B2(new_n252), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n304), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n317), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n588), .A2(G472), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n691), .A2(new_n580), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  NOR3_X1   g513(.A1(new_n672), .A2(new_n404), .A3(new_n679), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n697), .A2(new_n700), .A3(new_n623), .A4(new_n696), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  NOR3_X1   g516(.A1(new_n398), .A2(new_n403), .A3(new_n322), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n453), .B1(new_n443), .B2(new_n448), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n672), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n320), .A2(new_n580), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G131), .ZN(G33));
  INV_X1    g526(.A(new_n607), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n705), .A2(new_n713), .A3(new_n635), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n320), .A2(new_n580), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n320), .A2(KEYINPUT108), .A3(new_n714), .A4(new_n580), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  INV_X1    g534(.A(new_n594), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n599), .ZN(new_n722));
  NAND2_X1  g536(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n599), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n615), .A2(new_n643), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n703), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n729), .B1(new_n728), .B2(KEYINPUT44), .ZN(new_n732));
  OR3_X1    g546(.A1(new_n731), .A2(KEYINPUT112), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT112), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n728), .A2(KEYINPUT44), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n421), .B1(new_n432), .B2(new_n415), .ZN(new_n737));
  INV_X1    g551(.A(new_n435), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n737), .B2(new_n429), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n427), .B1(new_n740), .B2(new_n422), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n446), .A2(new_n441), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n736), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n447), .A2(KEYINPUT45), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(G469), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n743), .A2(new_n744), .A3(new_n747), .A4(G469), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n444), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n443), .B1(new_n749), .B2(KEYINPUT46), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n751), .B(new_n444), .C1(new_n746), .C2(new_n748), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n451), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(new_n646), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n735), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n733), .A2(new_n734), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  INV_X1    g571(.A(new_n703), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n320), .A2(new_n580), .A3(new_n672), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(KEYINPUT47), .B(new_n451), .C1(new_n750), .C2(new_n752), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  INV_X1    g579(.A(KEYINPUT120), .ZN(new_n766));
  NOR2_X1   g580(.A1(G952), .A2(G953), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n579), .B1(new_n660), .B2(new_n289), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n768), .A2(new_n542), .B1(new_n615), .B2(new_n625), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n288), .B1(new_n658), .B2(new_n659), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n631), .A2(new_n455), .A3(new_n636), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n701), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT52), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n406), .A2(new_n456), .A3(new_n601), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT114), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n406), .A2(new_n456), .A3(new_n600), .A4(new_n607), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n406), .A2(new_n777), .A3(new_n601), .A4(new_n456), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n615), .A3(new_n587), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n769), .A2(new_n773), .A3(KEYINPUT53), .A4(new_n780), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n623), .A2(new_n706), .A3(new_n697), .A4(new_n696), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n643), .A2(new_n533), .A3(new_n635), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n455), .A3(new_n703), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n783), .B1(new_n770), .B2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n784), .A2(new_n455), .A3(new_n703), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n320), .A2(new_n787), .A3(KEYINPUT115), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n782), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n719), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n781), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n594), .A2(new_n599), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n631), .A2(new_n455), .A3(new_n793), .A4(new_n671), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n770), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n772), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n641), .A2(new_n404), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n643), .A2(new_n704), .A3(new_n671), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n665), .B2(new_n666), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n801), .A2(KEYINPUT52), .B1(new_n709), .B2(new_n710), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n796), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n681), .A2(new_n689), .A3(new_n698), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(KEYINPUT116), .A3(new_n686), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n681), .A2(new_n686), .A3(new_n689), .A4(new_n698), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n791), .A2(new_n802), .A3(new_n804), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  INV_X1    g626(.A(new_n799), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n657), .B2(new_n662), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n638), .A2(new_n674), .A3(new_n701), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n804), .A2(new_n816), .A3(new_n711), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n626), .B(new_n581), .C1(new_n818), .C2(new_n593), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n681), .A2(new_n686), .A3(new_n689), .A4(new_n698), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n719), .A3(new_n821), .A4(new_n789), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n812), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n824));
  AND3_X1   g638(.A1(new_n811), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n805), .A2(new_n769), .A3(new_n686), .A4(new_n780), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n790), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n773), .A2(new_n812), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n802), .A3(new_n804), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n826), .B1(new_n830), .B2(new_n823), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n632), .B1(new_n724), .B2(new_n726), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n758), .A2(new_n679), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n697), .A2(new_n623), .A3(new_n696), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n323), .B(new_n679), .C1(KEYINPUT119), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(new_n651), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n697), .A2(new_n580), .A3(new_n696), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n842), .A3(new_n833), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n838), .A2(KEYINPUT119), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n678), .A2(new_n453), .A3(new_n443), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n761), .A2(new_n762), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n844), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n847), .A2(new_n703), .B1(new_n848), .B2(new_n840), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n842), .A2(new_n833), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n837), .B(new_n845), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n834), .A2(new_n580), .A3(new_n535), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n594), .A2(new_n599), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n852), .B(new_n854), .C1(new_n667), .C2(new_n663), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT118), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT51), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  OAI211_X1 g672(.A(KEYINPUT118), .B(new_n858), .C1(new_n851), .C2(new_n855), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n850), .A2(new_n404), .A3(new_n679), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n534), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n835), .A2(new_n770), .A3(new_n579), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT48), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n852), .B1(new_n667), .B2(new_n663), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n866), .B1(new_n793), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n857), .A2(new_n859), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n767), .B1(new_n832), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n667), .A2(new_n663), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n678), .A2(new_n443), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(KEYINPUT49), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT113), .Z(new_n874));
  NAND3_X1  g688(.A1(new_n580), .A2(new_n323), .A3(new_n451), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n722), .B(new_n875), .C1(KEYINPUT49), .C2(new_n872), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n871), .A2(new_n651), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n766), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n857), .A2(new_n859), .A3(new_n868), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n825), .A3(new_n831), .ZN(new_n881));
  OAI211_X1 g695(.A(KEYINPUT120), .B(new_n877), .C1(new_n881), .C2(new_n767), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(G75));
  AOI21_X1  g697(.A(new_n378), .B1(new_n811), .B2(new_n823), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(KEYINPUT121), .A3(G210), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n395), .B(new_n397), .Z(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT121), .B1(new_n884), .B2(G210), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n254), .A2(G952), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n884), .B2(G210), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n888), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n891), .A2(new_n895), .ZN(G51));
  NAND2_X1  g710(.A1(new_n811), .A2(new_n823), .ZN(new_n897));
  INV_X1    g711(.A(new_n824), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n811), .A2(new_n823), .A3(new_n824), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(KEYINPUT122), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n902), .A3(new_n898), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n444), .B(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n677), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n884), .A2(new_n748), .A3(new_n746), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n892), .B1(new_n907), .B2(new_n908), .ZN(G54));
  NOR2_X1   g723(.A1(new_n513), .A2(new_n527), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(KEYINPUT58), .A2(G475), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n884), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n884), .B2(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n892), .ZN(G60));
  XOR2_X1   g729(.A(new_n595), .B(KEYINPUT59), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n830), .A2(new_n823), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT54), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n918), .B2(new_n900), .ZN(new_n919));
  INV_X1    g733(.A(new_n598), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n893), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n901), .A2(new_n903), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n598), .A2(new_n916), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G63));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT125), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n926), .B(new_n927), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n897), .A2(new_n620), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n928), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n811), .B2(new_n823), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n571), .B(KEYINPUT126), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n929), .B(new_n893), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT61), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT61), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(G66));
  OAI21_X1  g752(.A(G953), .B1(new_n538), .B2(new_n330), .ZN(new_n939));
  INV_X1    g753(.A(new_n827), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(G953), .ZN(new_n941));
  INV_X1    g755(.A(new_n395), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(G898), .B2(new_n254), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  NAND2_X1  g758(.A1(new_n282), .A2(new_n283), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(new_n524), .Z(new_n946));
  NAND2_X1  g760(.A1(G900), .A2(G953), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n754), .A2(new_n797), .ZN(new_n948));
  AOI22_X1  g762(.A1(new_n948), .A2(new_n768), .B1(new_n763), .B2(new_n759), .ZN(new_n949));
  AND4_X1   g763(.A1(new_n711), .A2(new_n949), .A3(new_n719), .A4(new_n796), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n756), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n946), .B(new_n947), .C1(new_n951), .C2(G953), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n668), .A2(new_n796), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n758), .B(new_n647), .C1(new_n792), .C2(new_n713), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n768), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n764), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n953), .B2(KEYINPUT62), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n756), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n254), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n946), .B(KEYINPUT127), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n952), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n254), .B1(G227), .B2(G900), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n963), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(new_n952), .C1(new_n960), .C2(new_n961), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(G72));
  INV_X1    g781(.A(new_n285), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n756), .A2(new_n940), .A3(new_n954), .A4(new_n958), .ZN(new_n969));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  AOI211_X1 g785(.A(new_n264), .B(new_n968), .C1(new_n969), .C2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n756), .A2(new_n950), .A3(new_n940), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n263), .B(new_n285), .C1(new_n973), .C2(new_n971), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n286), .B1(new_n296), .B2(new_n301), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n917), .A2(new_n971), .A3(new_n975), .ZN(new_n976));
  NOR4_X1   g790(.A1(new_n972), .A2(new_n974), .A3(new_n892), .A4(new_n976), .ZN(G57));
endmodule


