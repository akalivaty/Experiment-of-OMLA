//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n207), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n207), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT0), .ZN(new_n219));
  AND2_X1   g0019(.A1(KEYINPUT64), .A2(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(KEYINPUT64), .A2(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(new_n203), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(new_n218), .A2(KEYINPUT0), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n215), .A2(new_n219), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n214), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n223), .B1(new_n207), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n222), .A2(G33), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n204), .A2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  INV_X1    g0054(.A(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n248), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n249), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n255), .A3(G1), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n249), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n260), .B1(new_n201), .B2(new_n269), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n258), .A2(new_n259), .B1(G50), .B2(new_n265), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT70), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  OAI211_X1 g0074(.A(G1), .B(G13), .C1(new_n248), .C2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G41), .A2(G45), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G1), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n277), .A3(G274), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT66), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n278), .B(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n276), .B2(G1), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G226), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n248), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G222), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G223), .A2(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n294), .B(new_n281), .C1(G77), .C2(new_n290), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n280), .A2(new_n286), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G169), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n272), .A2(new_n273), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n273), .B1(new_n272), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n296), .A2(G179), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT71), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n296), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n296), .ZN(new_n307));
  INV_X1    g0107(.A(new_n272), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n272), .A2(KEYINPUT74), .A3(KEYINPUT9), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT74), .B1(new_n272), .B2(KEYINPUT9), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n310), .B(new_n315), .C1(new_n312), .C2(new_n311), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n304), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n269), .A2(new_n203), .ZN(new_n318));
  INV_X1    g0118(.A(new_n265), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT12), .B1(new_n319), .B2(new_n203), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT12), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n265), .A2(new_n321), .A3(G68), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n318), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G20), .A2(G33), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n325));
  INV_X1    g0125(.A(G77), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n250), .B2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n327), .A2(KEYINPUT76), .A3(new_n249), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT76), .B1(new_n327), .B2(new_n249), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT11), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT11), .B1(new_n328), .B2(new_n329), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n323), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n285), .A2(G238), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n234), .A2(G1698), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(G226), .B2(G1698), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n336), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n281), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n280), .A2(new_n335), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n280), .A2(new_n335), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n344), .B1(KEYINPUT75), .B2(new_n345), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT75), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n347), .A2(new_n353), .A3(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(G179), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n350), .B1(new_n349), .B2(G169), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n334), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G200), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n346), .B2(new_n348), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n334), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n352), .A2(G190), .A3(new_n354), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT77), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT77), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n358), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n265), .A2(G77), .ZN(new_n368));
  INV_X1    g0168(.A(new_n269), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(G77), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n222), .A2(new_n326), .B1(new_n251), .B2(new_n256), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT72), .ZN(new_n372));
  XOR2_X1   g0172(.A(KEYINPUT15), .B(G87), .Z(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n250), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n371), .A2(KEYINPUT72), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n249), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n285), .A2(G244), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G238), .A2(G1698), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n290), .B(new_n381), .C1(new_n234), .C2(G1698), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n382), .B(new_n281), .C1(G107), .C2(new_n290), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n280), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G200), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT73), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n370), .A2(new_n385), .A3(KEYINPUT73), .A4(new_n377), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n306), .B2(new_n384), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n384), .A2(G179), .ZN(new_n390));
  INV_X1    g0190(.A(G169), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n378), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n317), .A2(new_n365), .A3(new_n367), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n319), .A2(new_n251), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n269), .B2(new_n251), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(G223), .A2(G1698), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G226), .B2(new_n291), .ZN(new_n401));
  INV_X1    g0201(.A(G87), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n401), .A2(new_n341), .B1(new_n248), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n285), .A2(G232), .B1(new_n403), .B2(new_n281), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n280), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n359), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n306), .A3(new_n280), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT78), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G58), .A2(G68), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n255), .B1(new_n225), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G159), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n256), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n410), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G58), .A2(G68), .ZN(new_n416));
  OAI21_X1  g0216(.A(G20), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n324), .A2(G159), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(KEYINPUT78), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n288), .A2(new_n255), .A3(new_n289), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n203), .B1(new_n421), .B2(KEYINPUT7), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n222), .A2(new_n341), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n420), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n249), .ZN(new_n427));
  OR2_X1    g0227(.A1(KEYINPUT64), .A2(G20), .ZN(new_n428));
  NAND2_X1  g0228(.A1(KEYINPUT64), .A2(G20), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT7), .B1(new_n430), .B2(new_n290), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n341), .A2(new_n423), .A3(new_n255), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(G68), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n411), .A2(new_n413), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT16), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n427), .A2(KEYINPUT79), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT79), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n414), .A2(new_n419), .B1(new_n422), .B2(new_n424), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n266), .B1(new_n438), .B2(KEYINPUT16), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n433), .A2(new_n434), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT16), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n437), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n399), .B(new_n408), .C1(new_n436), .C2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT80), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT79), .B1(new_n427), .B2(new_n435), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n439), .A2(new_n437), .A3(new_n442), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n398), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT80), .B1(new_n449), .B2(new_n408), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT17), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n399), .B1(new_n436), .B2(new_n443), .ZN(new_n453));
  INV_X1    g0253(.A(G179), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n405), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n391), .B1(new_n404), .B2(new_n280), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n452), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n449), .A2(KEYINPUT18), .A3(new_n457), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n444), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n451), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n396), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n250), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n402), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n336), .A2(new_n467), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n430), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n428), .B(new_n429), .C1(new_n339), .C2(new_n340), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n469), .B(new_n473), .C1(new_n203), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n249), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n319), .A2(new_n374), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n267), .A2(G33), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n479), .B(KEYINPUT83), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n265), .A2(new_n266), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(G87), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G45), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n483), .A2(G1), .A3(G274), .ZN(new_n484));
  AOI21_X1  g0284(.A(G250), .B1(new_n267), .B2(G45), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n281), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G244), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G1698), .ZN(new_n488));
  OAI221_X1 g0288(.A(new_n488), .B1(G238), .B2(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n486), .B1(new_n491), .B2(new_n281), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n359), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(G190), .B2(new_n492), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n482), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n265), .A2(new_n266), .A3(new_n480), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n476), .B(new_n477), .C1(new_n374), .C2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n492), .A2(G169), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n454), .B2(new_n492), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n319), .A2(new_n468), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n496), .B2(new_n468), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n431), .A2(G107), .A3(new_n432), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n324), .A2(G77), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT81), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT6), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n509), .A2(new_n468), .A3(G107), .ZN(new_n510));
  XNOR2_X1  g0310(.A(G97), .B(G107), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n508), .B1(new_n222), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n249), .B1(new_n505), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n249), .C1(new_n505), .C2(new_n513), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n503), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT5), .ZN(new_n520));
  AOI211_X1 g0320(.A(G1), .B(new_n483), .C1(new_n520), .C2(G41), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT85), .B1(new_n520), .B2(G41), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT85), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n274), .A3(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n281), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G257), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n521), .A2(G274), .A3(new_n275), .A4(new_n525), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G250), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT84), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n291), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  OAI211_X1 g0333(.A(G244), .B(new_n291), .C1(new_n339), .C2(new_n340), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n529), .B1(new_n537), .B2(new_n281), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n454), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n530), .B(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(new_n532), .A3(new_n533), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n281), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n527), .A3(new_n528), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n391), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n519), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(G200), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT86), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n538), .B2(G190), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n544), .A2(KEYINPUT86), .A3(new_n306), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n518), .B(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT25), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n265), .B2(G107), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n470), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n554), .A2(new_n555), .B1(new_n481), .B2(G107), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT87), .B1(new_n474), .B2(new_n402), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT87), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n290), .A2(new_n222), .A3(new_n558), .A4(G87), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(KEYINPUT22), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT88), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT22), .A4(new_n559), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n474), .A2(new_n402), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n222), .A2(KEYINPUT23), .A3(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n255), .A2(G33), .A3(G116), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT23), .B1(new_n255), .B2(G107), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT24), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT24), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n567), .A2(new_n575), .A3(new_n572), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT89), .B1(new_n577), .B2(new_n249), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n560), .A2(KEYINPUT88), .B1(new_n565), .B2(new_n564), .ZN(new_n579));
  AOI211_X1 g0379(.A(KEYINPUT24), .B(new_n571), .C1(new_n579), .C2(new_n563), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n575), .B1(new_n567), .B2(new_n572), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT89), .B(new_n249), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n556), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n290), .A2(G250), .A3(new_n291), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n290), .A2(G257), .A3(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G294), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n281), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n526), .A2(G264), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n590), .A3(new_n528), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(G179), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n391), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n584), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n359), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G190), .B2(new_n591), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n556), .B(new_n596), .C1(new_n578), .C2(new_n583), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n533), .B1(new_n468), .B2(G33), .ZN(new_n600));
  OAI221_X1 g0400(.A(new_n249), .B1(new_n255), .B2(G116), .C1(new_n430), .C2(new_n600), .ZN(new_n601));
  XOR2_X1   g0401(.A(new_n601), .B(KEYINPUT20), .Z(new_n602));
  NAND2_X1  g0402(.A1(new_n481), .A2(G116), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n602), .B(new_n603), .C1(G116), .C2(new_n265), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n526), .A2(G270), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n291), .A2(G257), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G264), .A2(G1698), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n290), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(G303), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n341), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n281), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n606), .A2(new_n528), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G169), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n599), .B1(new_n605), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n604), .A2(KEYINPUT21), .A3(G169), .A4(new_n613), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n528), .ZN(new_n617));
  INV_X1    g0417(.A(G270), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n618), .B(new_n281), .C1(new_n521), .C2(new_n525), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n604), .A2(G179), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n615), .A2(new_n616), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(G190), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n359), .B2(new_n620), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n604), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n598), .A2(new_n626), .ZN(new_n627));
  NOR4_X1   g0427(.A1(new_n466), .A2(new_n501), .A3(new_n552), .A4(new_n627), .ZN(G372));
  NAND3_X1  g0428(.A1(new_n453), .A2(new_n452), .A3(new_n458), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT18), .B1(new_n449), .B2(new_n457), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n363), .A2(new_n394), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n358), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n444), .A2(new_n445), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n449), .A2(KEYINPUT80), .A3(new_n408), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n462), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n463), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n631), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n314), .ZN(new_n640));
  INV_X1    g0440(.A(new_n316), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n303), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n500), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n482), .B2(new_n494), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n518), .B1(new_n391), .B2(new_n544), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT26), .A4(new_n539), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n501), .B2(new_n546), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n622), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT90), .B1(new_n584), .B2(new_n593), .ZN(new_n654));
  INV_X1    g0454(.A(new_n556), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n249), .B1(new_n580), .B2(new_n581), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n658), .B2(new_n582), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  INV_X1    g0460(.A(new_n593), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n653), .B1(new_n654), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n546), .A2(new_n551), .A3(new_n495), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n597), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n652), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n644), .B1(new_n466), .B2(new_n667), .ZN(G369));
  NAND3_X1  g0468(.A1(new_n222), .A2(new_n267), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n626), .B1(new_n605), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT91), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n622), .A2(new_n604), .A3(new_n674), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n677), .B1(new_n676), .B2(new_n678), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n584), .A2(new_n593), .A3(new_n674), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n594), .A2(new_n597), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n659), .A2(new_n675), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n584), .A2(KEYINPUT90), .A3(new_n593), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n675), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n653), .A2(new_n674), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n598), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n688), .A2(new_n691), .A3(new_n693), .ZN(G399));
  NAND2_X1  g0494(.A1(new_n216), .A2(new_n274), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n267), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n471), .A2(G116), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n227), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  AOI21_X1  g0500(.A(new_n622), .B1(new_n584), .B2(new_n593), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n651), .B1(new_n701), .B2(new_n665), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n663), .A2(new_n666), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n674), .B1(new_n704), .B2(new_n651), .ZN(new_n705));
  XNOR2_X1  g0505(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n703), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n552), .A2(new_n501), .A3(new_n674), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n594), .A2(new_n709), .A3(new_n597), .A4(new_n626), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n589), .A2(new_n492), .A3(new_n590), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n606), .A2(G179), .A3(new_n528), .A4(new_n612), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT30), .B1(new_n713), .B2(new_n538), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n492), .A2(G179), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n591), .A2(new_n715), .A3(new_n613), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n538), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT92), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n588), .A2(new_n281), .B1(new_n526), .B2(G264), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n620), .A2(G179), .A3(new_n720), .A4(new_n492), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n721), .B2(new_n544), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT92), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n544), .A2(new_n591), .A3(new_n613), .A4(new_n715), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n713), .A2(new_n538), .A3(KEYINPUT30), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n718), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n674), .A2(KEYINPUT31), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n727), .A2(KEYINPUT93), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT93), .B1(new_n727), .B2(new_n728), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n722), .A2(new_n726), .A3(new_n724), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n731), .B2(new_n674), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n710), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n708), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n700), .B1(new_n736), .B2(G1), .ZN(G364));
  OAI21_X1  g0537(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n738));
  INV_X1    g0538(.A(new_n682), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(G330), .A3(new_n679), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n430), .A2(new_n261), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G45), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n697), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n738), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n676), .A2(new_n678), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n744), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n290), .A2(new_n216), .ZN(new_n751));
  INV_X1    g0551(.A(G355), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(new_n752), .B1(G116), .B2(new_n216), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n243), .A2(G45), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n341), .A2(new_n216), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n483), .B2(new_n227), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n223), .B1(G20), .B2(new_n391), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n748), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT96), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n750), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT97), .Z(new_n762));
  NOR2_X1   g0562(.A1(G179), .A2(G200), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n430), .A2(new_n306), .A3(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G159), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT32), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n222), .A2(new_n454), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G190), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(G68), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n359), .A2(G179), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n430), .A2(new_n306), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n470), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n772), .A2(G20), .A3(G190), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT98), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT98), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n402), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n222), .A2(new_n454), .A3(G190), .A4(G200), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n774), .B(new_n779), .C1(G77), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n763), .A2(G190), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n430), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n306), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n768), .A2(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n290), .B1(new_n783), .B2(new_n468), .C1(new_n785), .C2(new_n202), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n769), .A2(new_n306), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(G50), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n771), .A2(new_n781), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G294), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n341), .B1(new_n783), .B2(new_n790), .C1(new_n778), .C2(new_n610), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G326), .B2(new_n787), .ZN(new_n792));
  INV_X1    g0592(.A(new_n773), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G311), .A2(new_n780), .B1(new_n793), .B2(G283), .ZN(new_n794));
  INV_X1    g0594(.A(new_n785), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G322), .B1(G329), .B2(new_n765), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n770), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n792), .A2(new_n794), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(KEYINPUT99), .B1(new_n789), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n758), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n789), .A2(new_n799), .A3(KEYINPUT99), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n762), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n749), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n745), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  OAI22_X1  g0607(.A1(new_n386), .A2(new_n388), .B1(new_n379), .B2(new_n675), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n393), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n394), .A2(new_n675), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n395), .A2(new_n675), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n705), .A2(new_n812), .B1(new_n667), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n750), .B1(new_n814), .B2(new_n735), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n735), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n758), .A2(new_n746), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT100), .Z(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n744), .B1(new_n326), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n793), .A2(G87), .ZN(new_n821));
  INV_X1    g0621(.A(new_n783), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n290), .B1(new_n822), .B2(G97), .ZN(new_n823));
  INV_X1    g0623(.A(new_n770), .ZN(new_n824));
  INV_X1    g0624(.A(G283), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n821), .B(new_n823), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G303), .B2(new_n787), .ZN(new_n827));
  INV_X1    g0627(.A(new_n778), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(G107), .B1(G116), .B2(new_n780), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n795), .A2(G294), .B1(G311), .B2(new_n765), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n795), .A2(G143), .B1(G159), .B2(new_n780), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n787), .A2(G137), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n254), .C2(new_n824), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT34), .Z(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n290), .B1(new_n764), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT101), .Z(new_n838));
  NAND2_X1  g0638(.A1(new_n828), .A2(G50), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n822), .A2(G58), .B1(new_n793), .B2(G68), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n831), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n758), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n820), .B1(new_n843), .B2(new_n845), .C1(new_n812), .C2(new_n747), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n816), .A2(new_n846), .ZN(G384));
  INV_X1    g0647(.A(new_n512), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(G116), .A3(new_n224), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT36), .Z(new_n852));
  NAND3_X1  g0652(.A1(new_n227), .A2(G77), .A3(new_n410), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n201), .A2(G68), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n267), .B(G13), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT104), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n622), .B1(new_n689), .B2(new_n690), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n651), .B1(new_n858), .B2(new_n665), .ZN(new_n859));
  INV_X1    g0659(.A(new_n813), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n859), .A2(new_n860), .B1(new_n394), .B2(new_n675), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n334), .A2(new_n862), .A3(new_n674), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n334), .B2(new_n674), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n364), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n358), .A2(new_n865), .A3(new_n363), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n857), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n810), .B1(new_n667), .B2(new_n813), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(KEYINPUT104), .A3(new_n869), .ZN(new_n873));
  INV_X1    g0673(.A(new_n672), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n453), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n634), .A2(new_n875), .A3(new_n635), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT106), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n453), .A2(new_n879), .A3(new_n458), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT106), .B1(new_n449), .B2(new_n457), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n439), .B1(KEYINPUT16), .B2(new_n438), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n399), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n458), .B2(new_n874), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n634), .A2(new_n885), .A3(new_n635), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n878), .A2(new_n882), .B1(KEYINPUT37), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n874), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n464), .A2(KEYINPUT105), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT105), .B1(new_n464), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT38), .B(new_n888), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n871), .A2(new_n873), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n631), .A2(new_n672), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n358), .A2(new_n674), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n895), .B2(new_n896), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT107), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n880), .A2(new_n881), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n905), .B2(new_n877), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n446), .A2(new_n450), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n449), .A2(new_n672), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n907), .A2(KEYINPUT107), .A3(new_n882), .A4(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n444), .B1(new_n457), .B2(new_n449), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT37), .B1(new_n911), .B2(new_n908), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n906), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n464), .A2(new_n908), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n894), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n896), .A2(new_n916), .A3(new_n902), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n901), .B1(new_n903), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n898), .A2(new_n899), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT108), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n465), .B(new_n703), .C1(new_n705), .C2(new_n707), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n644), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n921), .B(new_n923), .Z(new_n924));
  AOI21_X1  g0724(.A(new_n732), .B1(new_n728), .B2(new_n731), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n710), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n811), .B1(new_n867), .B2(new_n868), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(KEYINPUT40), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n896), .B2(new_n916), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n927), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT105), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n636), .A2(new_n631), .A3(new_n637), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n932), .B1(new_n933), .B2(new_n889), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n464), .A2(KEYINPUT105), .A3(new_n890), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n936), .B2(new_n888), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n894), .B(new_n887), .C1(new_n934), .C2(new_n935), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n931), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n929), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT110), .Z(new_n943));
  NAND2_X1  g0743(.A1(new_n465), .A2(new_n926), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n681), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n924), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n267), .B2(new_n741), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n924), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n856), .B1(new_n949), .B2(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n482), .A2(new_n675), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT111), .Z(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(new_n645), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(KEYINPUT112), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(KEYINPUT112), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n953), .A2(new_n501), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT43), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n546), .B(new_n551), .C1(new_n518), .C2(new_n675), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n647), .A2(new_n539), .A3(new_n674), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n598), .A2(new_n692), .A3(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT42), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n546), .B1(new_n594), .B2(new_n962), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n965), .A2(KEYINPUT42), .B1(new_n675), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n960), .A2(new_n961), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n968), .A3(new_n958), .A4(new_n959), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n964), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n688), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT113), .B(KEYINPUT41), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n695), .B(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n683), .A2(KEYINPUT114), .A3(new_n687), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n693), .A2(new_n691), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(new_n973), .ZN(new_n982));
  AOI211_X1 g0782(.A(KEYINPUT44), .B(new_n964), .C1(new_n693), .C2(new_n691), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n981), .B2(new_n973), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n691), .A4(new_n964), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n979), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n684), .B1(new_n653), .B2(new_n674), .C1(new_n685), .C2(new_n686), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n693), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n683), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n740), .A2(new_n693), .A3(new_n991), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n735), .A3(new_n708), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n984), .A2(new_n979), .A3(new_n988), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n990), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n978), .B1(new_n999), .B2(new_n736), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n743), .A2(G1), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n975), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n958), .A2(new_n748), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n238), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n759), .B1(new_n216), .B2(new_n374), .C1(new_n1004), .C2(new_n755), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n750), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n828), .A2(G116), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT46), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n773), .A2(new_n468), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G317), .B2(new_n765), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n780), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1008), .B(new_n1010), .C1(new_n825), .C2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n341), .B1(new_n783), .B2(new_n470), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G303), .B2(new_n795), .ZN(new_n1014));
  INV_X1    g0814(.A(G311), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n787), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1014), .B1(new_n824), .B2(new_n790), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(KEYINPUT115), .B(G137), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G77), .A2(new_n793), .B1(new_n765), .B2(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n202), .B2(new_n778), .C1(new_n254), .C2(new_n785), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n290), .B1(new_n783), .B2(new_n203), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G50), .B2(new_n780), .ZN(new_n1022));
  INV_X1    g0822(.A(G143), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1022), .B1(new_n824), .B2(new_n412), .C1(new_n1023), .C2(new_n1016), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1012), .A2(new_n1017), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT47), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1006), .B1(new_n1026), .B2(new_n758), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1003), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1002), .A2(new_n1028), .ZN(G387));
  NAND2_X1  g0829(.A1(new_n708), .A2(new_n735), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(new_n994), .A3(new_n993), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1031), .A2(new_n274), .A3(new_n216), .A4(new_n996), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n684), .B(new_n748), .C1(new_n685), .C2(new_n686), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n751), .A2(new_n698), .B1(G107), .B2(new_n216), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n235), .A2(G45), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n698), .ZN(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n1036), .C1(G68), .C2(G77), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n251), .A2(G50), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n755), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n750), .B1(new_n1041), .B2(new_n760), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1016), .A2(new_n412), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n783), .A2(new_n374), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1043), .A2(new_n341), .A3(new_n1009), .A4(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n778), .A2(new_n326), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1011), .A2(new_n203), .B1(new_n201), .B2(new_n785), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(G150), .C2(new_n765), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1045), .B(new_n1048), .C1(new_n251), .C2(new_n824), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n290), .B1(new_n765), .B2(G326), .ZN(new_n1050));
  INV_X1    g0850(.A(G116), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n778), .A2(new_n790), .B1(new_n825), .B2(new_n783), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n795), .A2(G317), .B1(G303), .B2(new_n780), .ZN(new_n1053));
  INV_X1    g0853(.A(G322), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1053), .B1(new_n824), .B2(new_n1015), .C1(new_n1054), .C2(new_n1016), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT49), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1050), .B1(new_n1051), .B2(new_n773), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1049), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1042), .B1(new_n1062), .B2(new_n758), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n995), .A2(new_n1001), .B1(new_n1033), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1032), .A2(new_n1064), .ZN(G393));
  NAND3_X1  g0865(.A1(new_n984), .A2(new_n688), .A3(new_n988), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1001), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n688), .B1(new_n984), .B2(new_n988), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n973), .A2(new_n748), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n759), .B1(new_n468), .B2(new_n216), .C1(new_n246), .C2(new_n755), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n750), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n787), .A2(G317), .B1(new_n795), .B2(G311), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  OAI22_X1  g0875(.A1(new_n778), .A2(new_n825), .B1(new_n1054), .B2(new_n764), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G294), .B2(new_n780), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n341), .B1(new_n783), .B2(new_n1051), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n774), .B(new_n1078), .C1(G303), .C2(new_n770), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1075), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n787), .A2(G150), .B1(new_n795), .B2(G159), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n778), .A2(new_n203), .B1(new_n1023), .B2(new_n764), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n251), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n780), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n821), .B(new_n290), .C1(new_n326), .C2(new_n783), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G50), .B2(new_n770), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1080), .B1(new_n1083), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1073), .B1(new_n1091), .B2(new_n758), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1070), .B1(new_n1071), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n996), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n999), .A3(new_n696), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(G390));
  NAND3_X1  g0896(.A1(new_n734), .A2(G330), .A3(new_n812), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n870), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n702), .A2(new_n675), .A3(new_n809), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n870), .B1(new_n1100), .B2(new_n810), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n896), .A2(new_n916), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n900), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(KEYINPUT39), .B1(new_n937), .B2(new_n938), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n917), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n901), .B1(new_n872), .B2(new_n869), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1099), .B(new_n1104), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n896), .A2(new_n916), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1109), .A2(new_n1101), .A3(new_n901), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n903), .A2(new_n918), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n900), .B1(new_n861), .B2(new_n870), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n681), .B1(new_n710), .B2(new_n925), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n927), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1108), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT117), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1097), .A2(new_n870), .B1(new_n927), .B2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n861), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n681), .B(new_n811), .C1(new_n710), .C2(new_n733), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1115), .B1(new_n1120), .B2(new_n869), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(KEYINPUT117), .A3(new_n872), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1100), .A2(new_n810), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n869), .B1(new_n1114), .B2(new_n812), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1098), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n465), .A2(new_n1114), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n922), .A2(new_n644), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1116), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1115), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1134), .A2(new_n1137), .A3(new_n1108), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(new_n696), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1001), .A3(new_n1108), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n750), .B1(new_n1085), .B2(new_n818), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n290), .B(new_n779), .C1(G77), .C2(new_n822), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n470), .B2(new_n824), .C1(new_n825), .C2(new_n1016), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G97), .A2(new_n780), .B1(new_n793), .B2(G68), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n1051), .B2(new_n785), .C1(new_n790), .C2(new_n764), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n770), .A2(new_n1018), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n787), .A2(G128), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n795), .A2(G132), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n341), .B1(new_n822), .B2(G159), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n778), .A2(new_n254), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT53), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G50), .A2(new_n793), .B1(new_n765), .B2(G125), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n1153), .C1(new_n1011), .C2(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1143), .A2(new_n1145), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1141), .B1(new_n1156), .B2(new_n758), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1106), .B2(new_n747), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1140), .A2(KEYINPUT118), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT118), .B1(new_n1140), .B2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1139), .B1(new_n1159), .B2(new_n1160), .ZN(G378));
  OAI21_X1  g0961(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n341), .B2(new_n274), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1046), .A2(G41), .A3(new_n290), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n793), .A2(G58), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n825), .C2(new_n764), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT119), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n795), .A2(G107), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G68), .A2(new_n822), .B1(new_n780), .B2(new_n373), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G97), .A2(new_n770), .B1(new_n787), .B2(G116), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1163), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1172), .B2(new_n1171), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(G41), .C1(new_n765), .C2(G124), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1154), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n828), .A2(new_n1176), .B1(G137), .B2(new_n780), .ZN(new_n1177));
  INV_X1    g0977(.A(G128), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n785), .C1(new_n836), .C2(new_n824), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n787), .A2(G125), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n254), .B2(new_n783), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1181), .A2(KEYINPUT120), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT120), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT59), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1175), .B1(new_n412), .B2(new_n773), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1185), .B2(new_n1184), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n758), .B1(new_n1174), .B2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n750), .C1(G50), .C2(new_n818), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n308), .A2(new_n874), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT55), .Z(new_n1191));
  XNOR2_X1  g0991(.A(new_n317), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1192), .B(new_n1193), .Z(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1189), .B1(new_n1195), .B2(new_n746), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1131), .B1(new_n1116), .B2(new_n1132), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n928), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1103), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n930), .B1(new_n895), .B2(new_n896), .ZN(new_n1200));
  OAI211_X1 g1000(.A(G330), .B(new_n1199), .C1(new_n1200), .C2(new_n940), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1201), .A2(new_n1195), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1194), .B1(new_n942), .B2(G330), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n920), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1195), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1106), .A2(new_n901), .B1(new_n631), .B2(new_n672), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n939), .A2(new_n941), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1207), .A2(G330), .A3(new_n1194), .A4(new_n1199), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .A4(new_n898), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1204), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1197), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT57), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n695), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1196), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT123), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1205), .A2(new_n1215), .A3(new_n1208), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT122), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n920), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1205), .A2(new_n1215), .A3(new_n1208), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n1217), .A3(new_n920), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1209), .A2(KEYINPUT123), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n696), .A2(new_n1212), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1138), .B2(new_n1131), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1001), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1214), .A2(new_n1226), .ZN(G375));
  AOI21_X1  g1027(.A(new_n1126), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT124), .B1(new_n1228), .B2(new_n1068), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n818), .A2(G68), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n290), .B(new_n1044), .C1(G77), .C2(new_n793), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n1051), .B2(new_n824), .C1(new_n790), .C2(new_n1016), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G107), .A2(new_n780), .B1(new_n765), .B2(G303), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n468), .B2(new_n778), .C1(new_n825), .C2(new_n785), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n290), .B1(new_n783), .B2(new_n201), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G58), .B2(new_n793), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n824), .B2(new_n1154), .C1(new_n836), .C2(new_n1016), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n795), .A2(new_n1018), .B1(G150), .B2(new_n780), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n1178), .B2(new_n764), .C1(new_n412), .C2(new_n778), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1232), .A2(new_n1234), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n744), .B(new_n1230), .C1(new_n1240), .C2(new_n758), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n869), .B2(new_n747), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1229), .A2(new_n1242), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1228), .A2(KEYINPUT124), .A3(new_n1068), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1228), .A2(new_n1130), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1132), .A2(new_n977), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(G381));
  NAND4_X1  g1048(.A1(new_n1002), .A2(new_n1028), .A3(new_n1095), .A4(new_n1093), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1032), .A2(new_n806), .A3(new_n1064), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(new_n1249), .A2(G384), .A3(G381), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(G378), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1226), .A4(new_n1214), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n673), .A2(G213), .ZN(new_n1254));
  OR3_X1    g1054(.A1(G375), .A2(G378), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(new_n1255), .A3(G213), .ZN(G409));
  INV_X1    g1056(.A(new_n974), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n972), .B(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n984), .A2(new_n979), .A3(new_n988), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(new_n989), .A3(new_n996), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n977), .B1(new_n1260), .B2(new_n1030), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1258), .B1(new_n1261), .B2(new_n1068), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1028), .ZN(new_n1263));
  OAI21_X1  g1063(.A(G390), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G393), .A2(G396), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1250), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1264), .A2(new_n1249), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1264), .B2(new_n1249), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1246), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1134), .A2(new_n695), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1123), .A2(new_n1130), .A3(KEYINPUT60), .A4(new_n1127), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT125), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(KEYINPUT125), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1272), .B(new_n1273), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(G384), .A3(new_n1245), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1277), .B2(new_n1245), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1214), .A2(new_n1226), .A3(G378), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n978), .B1(new_n1138), .B2(new_n1131), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1223), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1196), .B1(new_n1210), .B2(new_n1001), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1254), .B(new_n1281), .C1(new_n1282), .C2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT126), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1252), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1214), .A2(new_n1226), .A3(G378), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1254), .A4(new_n1281), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1288), .A2(new_n1289), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1254), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n673), .A2(G213), .A3(G2897), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1277), .A2(new_n1245), .ZN(new_n1301));
  INV_X1    g1101(.A(G384), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n1278), .A3(new_n1298), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1297), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1270), .B1(new_n1296), .B2(new_n1309), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1291), .A2(new_n1292), .B1(G213), .B2(new_n673), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1269), .B(new_n1308), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1287), .A2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT63), .B1(new_n1288), .B2(new_n1295), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1316), .B1(new_n1317), .B2(KEYINPUT127), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n1319), .B(KEYINPUT63), .C1(new_n1288), .C2(new_n1295), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1310), .B1(new_n1318), .B2(new_n1320), .ZN(G405));
  XNOR2_X1  g1121(.A(G375), .B(G378), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1270), .A2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1270), .A2(new_n1322), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1281), .ZN(new_n1325));
  OR3_X1    g1125(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1325), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


