//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT92), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n205), .A2(new_n206), .A3(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT92), .B1(new_n208), .B2(KEYINPUT16), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n203), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(KEYINPUT93), .A3(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n211), .B(G8gat), .C1(KEYINPUT93), .C2(new_n210), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n210), .A2(KEYINPUT94), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(KEYINPUT94), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n204), .A4(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT89), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT14), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n218), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n218), .A2(new_n220), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(KEYINPUT15), .B2(new_n217), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n226), .B(KEYINPUT90), .Z(new_n230));
  OAI21_X1  g029(.A(new_n227), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT17), .B1(new_n231), .B2(new_n232), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n212), .B(new_n216), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n212), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n231), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n202), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n241), .A4(new_n239), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n238), .B(new_n231), .Z(new_n245));
  XOR2_X1   g044(.A(new_n241), .B(KEYINPUT13), .Z(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G169gat), .B(G197gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT12), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n255), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n243), .A2(new_n244), .A3(new_n248), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT87), .ZN(new_n261));
  AND2_X1   g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262));
  INV_X1    g061(.A(G169gat), .ZN(new_n263));
  INV_X1    g062(.A(G176gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(G190gat), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT23), .ZN(new_n271));
  INV_X1    g070(.A(G190gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n267), .A2(new_n270), .A3(new_n271), .A4(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n266), .B1(G169gat), .B2(G176gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT64), .ZN(new_n276));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n271), .A2(new_n275), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT25), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n269), .A2(G190gat), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n272), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(new_n268), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n271), .A2(new_n275), .A3(new_n277), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n283), .A2(new_n284), .B1(new_n278), .B2(KEYINPUT25), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n265), .B(KEYINPUT65), .C1(new_n262), .C2(KEYINPUT26), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n265), .B2(KEYINPUT26), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT26), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(KEYINPUT66), .A3(new_n293), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n286), .A2(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G183gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT27), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G183gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n299), .A3(new_n272), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT28), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT27), .B(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n272), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI22_X1  g105(.A1(new_n280), .A2(new_n285), .B1(new_n295), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G120gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G113gat), .ZN(new_n309));
  INV_X1    g108(.A(G113gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G120gat), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT1), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G127gat), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT67), .B1(new_n315), .B2(G134gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(G134gat), .ZN(new_n317));
  INV_X1    g116(.A(G134gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G127gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(new_n320), .B2(KEYINPUT67), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n314), .B1(new_n321), .B2(new_n312), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G227gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n286), .A2(new_n290), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n292), .A2(new_n294), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n274), .A2(new_n279), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT64), .A4(KEYINPUT25), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n334), .A3(new_n322), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n324), .A2(new_n326), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(G15gat), .B(G43gat), .Z(new_n339));
  XNOR2_X1  g138(.A(G71gat), .B(G99gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT34), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n325), .B2(KEYINPUT68), .ZN(new_n344));
  AOI211_X1 g143(.A(new_n326), .B(new_n344), .C1(new_n324), .C2(new_n335), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n324), .A2(new_n335), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n325), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n344), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n342), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n344), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n347), .B2(new_n325), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n338), .B(new_n341), .C1(new_n352), .C2(new_n345), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n350), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n350), .B2(new_n353), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT35), .ZN(new_n359));
  XNOR2_X1  g158(.A(G197gat), .B(G204gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT22), .ZN(new_n361));
  INV_X1    g160(.A(G211gat), .ZN(new_n362));
  INV_X1    g161(.A(G218gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n360), .A3(new_n364), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(KEYINPUT70), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n365), .A2(new_n371), .A3(new_n367), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT71), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(KEYINPUT71), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  INV_X1    g177(.A(G141gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G148gat), .ZN(new_n380));
  INV_X1    g179(.A(G148gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G141gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n380), .A2(new_n382), .B1(KEYINPUT2), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n385));
  INV_X1    g184(.A(new_n383), .ZN(new_n386));
  NOR2_X1   g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G155gat), .ZN(new_n389));
  INV_X1    g188(.A(G162gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT76), .A3(new_n383), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n384), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n383), .ZN(new_n394));
  XNOR2_X1  g193(.A(G141gat), .B(G148gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT2), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(G155gat), .B2(G162gat), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n394), .B(new_n385), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT77), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT77), .ZN(new_n402));
  AOI211_X1 g201(.A(new_n402), .B(KEYINPUT3), .C1(new_n393), .C2(new_n398), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n378), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n400), .B1(new_n373), .B2(KEYINPUT29), .ZN(new_n407));
  INV_X1    g206(.A(new_n399), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n406), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n368), .A2(new_n412), .A3(new_n369), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(new_n378), .C1(new_n412), .C2(new_n369), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n400), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n377), .A2(new_n404), .B1(new_n415), .B2(new_n408), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n410), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G22gat), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n410), .B(new_n420), .C1(new_n416), .C2(new_n411), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G50gat), .ZN(new_n423));
  XOR2_X1   g222(.A(G78gat), .B(G106gat), .Z(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND4_X1  g224(.A1(new_n418), .A2(new_n419), .A3(new_n421), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n418), .A2(new_n421), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n421), .A2(KEYINPUT85), .ZN(new_n428));
  INV_X1    g227(.A(new_n425), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n358), .A2(new_n359), .A3(new_n426), .A4(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n377), .ZN(new_n433));
  INV_X1    g232(.A(G226gat), .ZN(new_n434));
  INV_X1    g233(.A(G233gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n330), .A2(new_n327), .B1(new_n332), .B2(new_n333), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(KEYINPUT29), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n331), .B2(new_n334), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n439), .B1(KEYINPUT72), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n442), .B(new_n437), .C1(new_n438), .C2(KEYINPUT29), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n433), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(KEYINPUT73), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT73), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n438), .B2(new_n437), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n433), .A2(new_n445), .A3(new_n439), .A4(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT74), .ZN(new_n451));
  XNOR2_X1  g250(.A(G8gat), .B(G36gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(G64gat), .B(G92gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  NAND4_X1  g253(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT30), .A4(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n436), .B1(new_n307), .B2(new_n378), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT72), .B1(new_n307), .B2(new_n436), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n443), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n377), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n459), .A2(KEYINPUT30), .A3(new_n448), .A4(new_n454), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n454), .B1(new_n459), .B2(new_n448), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(KEYINPUT74), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n448), .A3(new_n454), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n463), .A2(KEYINPUT75), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT75), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n455), .B(new_n462), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n393), .A2(KEYINPUT3), .A3(new_n398), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n468), .A2(new_n322), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n401), .B2(new_n403), .ZN(new_n470));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n313), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n309), .A2(new_n311), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n473), .A2(new_n316), .B1(KEYINPUT1), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n399), .A2(new_n475), .A3(new_n314), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n323), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n470), .A2(new_n471), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n481));
  NAND3_X1  g280(.A1(new_n322), .A2(new_n398), .A3(new_n393), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n471), .B1(new_n482), .B2(new_n476), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(KEYINPUT78), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n485));
  AOI211_X1 g284(.A(new_n485), .B(new_n471), .C1(new_n482), .C2(new_n476), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n480), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(G1gat), .B(G29gat), .Z(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G85gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n478), .A2(new_n479), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(new_n471), .A3(new_n470), .A4(new_n481), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n487), .A2(KEYINPUT6), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n487), .A2(new_n494), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n498), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n492), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n494), .ZN(new_n503));
  INV_X1    g302(.A(new_n492), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n497), .A2(new_n499), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n467), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n261), .B1(new_n432), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n462), .A2(new_n455), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n501), .A3(new_n500), .ZN(new_n510));
  INV_X1    g309(.A(new_n497), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n463), .A2(new_n464), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n463), .A2(KEYINPUT75), .A3(new_n464), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n509), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n519), .A2(new_n431), .A3(KEYINPUT87), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n350), .A2(new_n353), .A3(new_n355), .ZN(new_n521));
  INV_X1    g320(.A(new_n357), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n430), .A2(new_n521), .A3(new_n522), .A4(new_n426), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT82), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n467), .B2(new_n506), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n509), .A2(new_n513), .A3(new_n518), .A4(KEYINPUT82), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI22_X1  g326(.A1(new_n508), .A2(new_n520), .B1(new_n527), .B2(new_n359), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n358), .B2(KEYINPUT69), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n522), .A2(new_n521), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT69), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT36), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n430), .A2(new_n426), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n525), .B2(new_n526), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT37), .B1(new_n444), .B2(new_n449), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n454), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n537), .B(new_n539), .C1(new_n461), .C2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n454), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n444), .B2(new_n449), .ZN(new_n544));
  INV_X1    g343(.A(new_n541), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n445), .A2(new_n439), .A3(new_n447), .A4(new_n377), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n540), .B1(new_n458), .B2(new_n433), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n542), .B1(new_n548), .B2(new_n539), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n506), .A3(new_n463), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT40), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n493), .A2(new_n470), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT39), .ZN(new_n553));
  INV_X1    g352(.A(new_n471), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n504), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n482), .A2(new_n476), .A3(new_n471), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT39), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n552), .B2(new_n554), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n551), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n500), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n556), .A2(new_n551), .A3(new_n559), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n467), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n534), .B1(new_n550), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n530), .B(new_n533), .C1(new_n536), .C2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n260), .B1(new_n528), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n570));
  AOI211_X1 g369(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(KEYINPUT7), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n570), .B2(KEYINPUT7), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT98), .B(G85gat), .Z(new_n573));
  NAND2_X1  g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n573), .A2(new_n569), .B1(KEYINPUT8), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n576));
  OAI211_X1 g375(.A(KEYINPUT97), .B(new_n576), .C1(new_n568), .C2(new_n569), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G99gat), .B(G106gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n235), .B2(new_n236), .ZN(new_n581));
  INV_X1    g380(.A(new_n579), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n578), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n231), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G190gat), .B(G218gat), .Z(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G134gat), .B(G162gat), .Z(new_n589));
  AOI21_X1  g388(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n591), .A2(KEYINPUT99), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(new_n587), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(KEYINPUT99), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT100), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G57gat), .B(G64gat), .Z(new_n605));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(KEYINPUT9), .B2(new_n602), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT20), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n614), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G183gat), .B(G211gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n238), .B1(KEYINPUT21), .B2(new_n611), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n601), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G230gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n435), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n580), .A2(new_n609), .A3(new_n610), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n583), .A2(new_n611), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n583), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n628), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n635), .B1(new_n629), .B2(new_n630), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G120gat), .B(G148gat), .Z(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n567), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT101), .Z(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n513), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n208), .ZN(G1324gat));
  INV_X1    g447(.A(new_n467), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n214), .B2(new_n650), .ZN(new_n653));
  MUX2_X1   g452(.A(new_n652), .B(new_n653), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g453(.A1(new_n530), .A2(new_n533), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT102), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n530), .A2(new_n533), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(G15gat), .B1(new_n646), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n531), .A2(G15gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n646), .B2(new_n662), .ZN(G1326gat));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n535), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  INV_X1    g465(.A(new_n625), .ZN(new_n667));
  INV_X1    g466(.A(new_n643), .ZN(new_n668));
  AND4_X1   g467(.A1(new_n567), .A2(new_n667), .A3(new_n600), .A4(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n221), .A3(new_n506), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n656), .B(new_n658), .C1(new_n536), .C2(new_n565), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n528), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n528), .A2(new_n673), .A3(new_n672), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n601), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n528), .A2(new_n566), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n600), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT105), .B1(new_n681), .B2(KEYINPUT44), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n601), .B1(new_n528), .B2(new_n566), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n679), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n643), .B(KEYINPUT103), .Z(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n667), .A3(new_n259), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT104), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n692), .A2(new_n506), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n671), .B1(new_n694), .B2(new_n221), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n669), .A2(new_n222), .A3(new_n467), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT46), .Z(new_n697));
  AND3_X1   g496(.A1(new_n692), .A2(new_n467), .A3(new_n693), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n698), .B2(new_n222), .ZN(G1329gat));
  OAI21_X1  g498(.A(G43gat), .B1(new_n691), .B2(new_n660), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n531), .A2(G43gat), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n669), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n692), .A2(new_n659), .A3(new_n693), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n702), .B1(new_n706), .B2(G43gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n707), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g507(.A(G50gat), .B1(new_n691), .B2(new_n535), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n535), .A2(G50gat), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n669), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n692), .A2(new_n534), .A3(new_n693), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n711), .B1(new_n715), .B2(G50gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n716), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g516(.A1(new_n675), .A2(new_n676), .ZN(new_n718));
  NOR4_X1   g517(.A1(new_n718), .A2(new_n259), .A3(new_n626), .A4(new_n688), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n506), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  INV_X1    g520(.A(new_n719), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n649), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  AND2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n723), .B2(new_n724), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n722), .B2(new_n660), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n531), .A2(G71gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n722), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g530(.A1(new_n719), .A2(new_n534), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n681), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n528), .A2(new_n673), .A3(new_n672), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n674), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n735), .A2(new_n736), .B1(new_n738), .B2(new_n678), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n625), .A2(new_n259), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n643), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n734), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n741), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n687), .A2(KEYINPUT109), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n742), .A2(new_n506), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n528), .A2(new_n673), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n601), .A2(new_n259), .A3(new_n625), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n746), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT51), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n643), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n506), .A2(new_n573), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n745), .A2(new_n573), .B1(new_n751), .B2(new_n752), .ZN(G1336gat));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n742), .A2(new_n467), .A3(new_n744), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G92gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n688), .A2(G92gat), .A3(new_n649), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n748), .B2(new_n749), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n754), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n687), .A2(new_n467), .A3(new_n743), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n754), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AOI211_X1 g564(.A(KEYINPUT110), .B(new_n763), .C1(new_n761), .C2(G92gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT111), .B1(new_n759), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n736), .A2(new_n735), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n741), .B1(new_n769), .B2(new_n679), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n569), .B1(new_n770), .B2(new_n467), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT110), .B1(new_n771), .B2(new_n763), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n762), .A2(new_n760), .A3(new_n764), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n755), .A2(G92gat), .B1(new_n750), .B2(new_n757), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n774), .B(new_n775), .C1(new_n776), .C2(new_n754), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n768), .A2(new_n777), .ZN(G1337gat));
  NAND3_X1  g577(.A1(new_n742), .A2(new_n659), .A3(new_n744), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G99gat), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n531), .A2(G99gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n751), .B2(new_n781), .ZN(G1338gat));
  INV_X1    g581(.A(G106gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n770), .B2(new_n534), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n688), .A2(G106gat), .A3(new_n535), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n750), .A2(new_n785), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n784), .A2(KEYINPUT53), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n742), .A2(new_n534), .A3(new_n744), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n788), .A2(new_n789), .A3(G106gat), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n788), .B2(G106gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n790), .A2(new_n791), .A3(new_n786), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(G1339gat));
  NAND2_X1  g593(.A1(new_n632), .A2(new_n633), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n635), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n632), .A2(new_n633), .A3(new_n628), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n640), .B1(new_n634), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n798), .A2(new_n800), .A3(new_n801), .A4(KEYINPUT55), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n642), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n798), .A2(new_n800), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT113), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n259), .A2(new_n803), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n245), .A2(new_n247), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT115), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n240), .A2(KEYINPUT114), .A3(new_n242), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT114), .B1(new_n240), .B2(new_n242), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n254), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n258), .A3(new_n643), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n808), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n808), .A2(KEYINPUT116), .A3(new_n815), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n601), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n600), .A2(new_n258), .A3(new_n814), .A4(new_n807), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n625), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n644), .A2(new_n260), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n467), .A2(new_n513), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n828), .A2(new_n358), .A3(new_n535), .A4(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n310), .A3(new_n260), .ZN(new_n831));
  INV_X1    g630(.A(new_n523), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n828), .A2(new_n506), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT117), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n259), .A3(new_n649), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n831), .B1(new_n835), .B2(new_n310), .ZN(G1340gat));
  OAI21_X1  g635(.A(G120gat), .B1(new_n830), .B2(new_n688), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT118), .Z(new_n838));
  NAND2_X1  g637(.A1(new_n834), .A2(new_n649), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n643), .A2(new_n308), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(G1341gat));
  OAI21_X1  g640(.A(G127gat), .B1(new_n830), .B2(new_n667), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n625), .A2(new_n315), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n839), .B2(new_n843), .ZN(G1342gat));
  NAND4_X1  g643(.A1(new_n834), .A2(new_n318), .A3(new_n649), .A4(new_n600), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n846));
  OAI21_X1  g645(.A(G134gat), .B1(new_n830), .B2(new_n601), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n660), .A2(new_n829), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n534), .B1(new_n825), .B2(new_n827), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n815), .A2(KEYINPUT120), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n804), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n798), .A2(KEYINPUT121), .A3(new_n800), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n259), .A2(new_n860), .A3(new_n806), .A4(new_n803), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n815), .A2(KEYINPUT120), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n855), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n823), .B1(new_n863), .B2(new_n601), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n826), .B1(new_n864), .B2(new_n625), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(KEYINPUT57), .A3(new_n534), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n854), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT119), .B1(new_n852), .B2(new_n853), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n259), .B(new_n851), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT123), .B1(new_n869), .B2(G141gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n660), .A2(new_n534), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n828), .A2(new_n506), .A3(new_n872), .ZN(new_n873));
  NOR4_X1   g672(.A1(new_n873), .A2(G141gat), .A3(new_n260), .A4(new_n467), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n869), .B2(G141gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n870), .A2(new_n875), .A3(KEYINPUT58), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  AOI221_X4 g676(.A(new_n874), .B1(KEYINPUT123), .B2(new_n877), .C1(new_n869), .C2(G141gat), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n828), .A2(KEYINPUT57), .A3(new_n534), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n534), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n853), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n882), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n643), .B(new_n851), .C1(new_n883), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n880), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n880), .A2(G148gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n867), .A2(new_n868), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n850), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n643), .ZN(new_n892));
  INV_X1    g691(.A(new_n873), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n649), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n643), .A2(new_n381), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n888), .A2(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1345gat));
  NOR3_X1   g695(.A1(new_n894), .A2(KEYINPUT125), .A3(new_n667), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(G155gat), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT125), .B1(new_n894), .B2(new_n667), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n667), .A2(new_n389), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n898), .A2(new_n899), .B1(new_n891), .B2(new_n900), .ZN(G1346gat));
  OAI211_X1 g700(.A(new_n600), .B(new_n851), .C1(new_n867), .C2(new_n868), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n390), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n903), .B2(new_n902), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n600), .A2(new_n390), .A3(new_n649), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n873), .B2(new_n906), .ZN(G1347gat));
  NOR3_X1   g706(.A1(new_n649), .A2(new_n506), .A3(new_n531), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n828), .A2(new_n535), .A3(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n263), .A3(new_n260), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n828), .A2(new_n513), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n467), .A3(new_n832), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n259), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n914), .B2(new_n263), .ZN(G1348gat));
  OAI21_X1  g714(.A(G176gat), .B1(new_n909), .B2(new_n688), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n643), .A2(new_n264), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n912), .B2(new_n917), .ZN(G1349gat));
  OAI21_X1  g717(.A(G183gat), .B1(new_n909), .B2(new_n667), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n625), .A2(new_n302), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n913), .A2(new_n272), .A3(new_n600), .ZN(new_n923));
  OAI21_X1  g722(.A(G190gat), .B1(new_n909), .B2(new_n601), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1351gat));
  NOR2_X1   g726(.A1(new_n871), .A2(new_n649), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT127), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(G197gat), .B1(new_n931), .B2(new_n259), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n883), .A2(new_n886), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n659), .A2(new_n506), .A3(new_n649), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n259), .A2(G197gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G1352gat));
  OAI21_X1  g737(.A(G204gat), .B1(new_n935), .B2(new_n688), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n930), .A2(G204gat), .A3(new_n668), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1353gat));
  NAND3_X1  g741(.A1(new_n931), .A2(new_n362), .A3(new_n625), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n625), .B(new_n934), .C1(new_n883), .C2(new_n886), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1354gat));
  OAI21_X1  g746(.A(G218gat), .B1(new_n935), .B2(new_n601), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n363), .A3(new_n600), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1355gat));
endmodule


