//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087;
  XOR2_X1   g000(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G107), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n195), .A2(KEYINPUT76), .A3(new_n196), .A4(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(new_n192), .A3(new_n196), .A4(new_n194), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n191), .A2(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n194), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n198), .A2(new_n201), .B1(G101), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G116), .B(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT5), .ZN(new_n206));
  INV_X1    g020(.A(G116), .ZN(new_n207));
  NOR3_X1   g021(.A1(new_n207), .A2(KEYINPUT5), .A3(G119), .ZN(new_n208));
  INV_X1    g022(.A(G113), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT2), .B(G113), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n206), .A2(new_n210), .B1(new_n212), .B2(new_n205), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n204), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n204), .A2(new_n213), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n189), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT72), .B(G125), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT0), .B(G128), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G143), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n230), .A3(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT66), .B1(new_n225), .B2(G146), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n223), .A3(G143), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n233), .A2(new_n235), .A3(new_n228), .A4(new_n226), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n218), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n225), .A2(G146), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g054(.A(G128), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n227), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(KEYINPUT1), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n233), .A2(new_n235), .A3(new_n226), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n237), .A2(new_n238), .B1(new_n247), .B2(new_n218), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n233), .A2(new_n235), .A3(new_n226), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n222), .A2(new_n231), .B1(new_n249), .B2(new_n228), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT82), .B1(new_n250), .B2(new_n218), .ZN(new_n251));
  INV_X1    g065(.A(G224), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT7), .B1(new_n252), .B2(G953), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n248), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n205), .B(new_n211), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n197), .A2(new_n192), .A3(new_n194), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(G101), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT78), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n257), .A2(new_n258), .A3(new_n261), .A4(G101), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(G101), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n199), .A2(new_n200), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n199), .A2(new_n200), .ZN(new_n266));
  OAI211_X1 g080(.A(KEYINPUT4), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n188), .A3(new_n214), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n217), .A2(new_n255), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n220), .A2(new_n221), .A3(new_n219), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT65), .B1(new_n227), .B2(new_n230), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n236), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G125), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT72), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G125), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n238), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n247), .A2(new_n218), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n251), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n253), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT85), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT85), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n285), .A3(new_n253), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n271), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n188), .B1(new_n268), .B2(new_n214), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(KEYINPUT81), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n290), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n263), .A2(new_n267), .B1(new_n204), .B2(new_n213), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n188), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n294), .B2(new_n288), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n252), .A2(G953), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT83), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n248), .B2(new_n251), .ZN(new_n298));
  AND4_X1   g112(.A1(new_n251), .A2(new_n280), .A3(new_n281), .A4(new_n297), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n287), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT87), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n303), .B(KEYINPUT86), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n284), .A2(new_n286), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n302), .B1(new_n307), .B2(new_n270), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n298), .A2(new_n299), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n269), .A2(new_n290), .ZN(new_n310));
  INV_X1    g124(.A(new_n288), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n309), .B1(new_n312), .B2(new_n291), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n306), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n284), .A2(new_n286), .ZN(new_n315));
  AOI21_X1  g129(.A(G902), .B1(new_n315), .B2(new_n271), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n301), .A4(new_n303), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n305), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT80), .B(G469), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n203), .A2(G101), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n265), .B2(new_n266), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n247), .ZN(new_n324));
  AND4_X1   g138(.A1(new_n233), .A2(new_n235), .A3(new_n226), .A4(new_n244), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n233), .A2(new_n235), .A3(new_n226), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT79), .B1(new_n328), .B2(new_n241), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n329), .B2(new_n325), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n204), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G137), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT11), .ZN(new_n334));
  INV_X1    g148(.A(G134), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT67), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G134), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(KEYINPUT11), .A3(G134), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT11), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G137), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G131), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n340), .A2(new_n342), .ZN(new_n345));
  INV_X1    g159(.A(G131), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT12), .B1(new_n332), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT12), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n339), .A2(G131), .A3(new_n343), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n346), .B1(new_n345), .B2(new_n347), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n351), .B(new_n354), .C1(new_n324), .C2(new_n331), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n331), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n260), .A2(new_n262), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n267), .A2(new_n250), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n247), .A2(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n204), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(new_n354), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G110), .B(G140), .ZN(new_n364));
  INV_X1    g178(.A(G227), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G953), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n364), .B(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n360), .A3(new_n362), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n349), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(new_n372), .B2(new_n363), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n302), .B(new_n321), .C1(new_n370), .C2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n363), .B1(new_n350), .B2(new_n355), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n367), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n363), .A2(new_n368), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n372), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G469), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n374), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT9), .B(G234), .ZN(new_n382));
  OAI21_X1  g196(.A(G221), .B1(new_n382), .B2(G902), .ZN(new_n383));
  OAI21_X1  g197(.A(G214), .B1(G237), .B2(G902), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT95), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n218), .A2(KEYINPUT16), .A3(G140), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT73), .ZN(new_n389));
  INV_X1    g203(.A(G140), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n276), .B2(new_n278), .ZN(new_n391));
  NOR2_X1   g205(.A1(G125), .A2(G140), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n389), .B(KEYINPUT16), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n392), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n218), .B2(new_n390), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n389), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n388), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n223), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n392), .B1(new_n279), .B2(G140), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT16), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT73), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n387), .B1(new_n402), .B2(new_n393), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G146), .ZN(new_n404));
  INV_X1    g218(.A(G237), .ZN(new_n405));
  INV_X1    g219(.A(G953), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(G214), .ZN(new_n407));
  AND2_X1   g221(.A1(KEYINPUT88), .A2(G143), .ZN(new_n408));
  NOR2_X1   g222(.A1(KEYINPUT88), .A2(G143), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(G237), .A2(G953), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n411), .B(G214), .C1(KEYINPUT88), .C2(G143), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G131), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT17), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n346), .A3(new_n412), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n346), .B1(new_n410), .B2(new_n412), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT17), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n399), .A2(new_n404), .A3(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(G113), .B(G122), .Z(new_n422));
  XOR2_X1   g236(.A(KEYINPUT92), .B(G104), .Z(new_n423));
  XOR2_X1   g237(.A(new_n422), .B(new_n423), .Z(new_n424));
  AND2_X1   g238(.A1(new_n424), .A2(KEYINPUT94), .ZN(new_n425));
  AND2_X1   g239(.A1(KEYINPUT89), .A2(KEYINPUT18), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n410), .A2(new_n346), .A3(new_n412), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n418), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n413), .A2(new_n426), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(G146), .B(new_n395), .C1(new_n218), .C2(new_n390), .ZN(new_n432));
  XNOR2_X1  g246(.A(G125), .B(G140), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n223), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n432), .A2(KEYINPUT90), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT90), .B1(new_n432), .B2(new_n434), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n431), .A2(new_n437), .A3(KEYINPUT91), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n414), .A2(new_n416), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n429), .B1(new_n440), .B2(new_n426), .ZN(new_n441));
  INV_X1    g255(.A(new_n436), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(KEYINPUT90), .A3(new_n434), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n421), .B(new_n425), .C1(new_n438), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n302), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT91), .B1(new_n431), .B2(new_n437), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n441), .A2(new_n444), .A3(new_n439), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n425), .B1(new_n450), .B2(new_n421), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n386), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n421), .B1(new_n438), .B2(new_n445), .ZN(new_n453));
  INV_X1    g267(.A(new_n425), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(KEYINPUT95), .A3(new_n302), .A4(new_n446), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(G475), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n424), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT19), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n433), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n396), .B2(new_n459), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G146), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n414), .B2(new_n416), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n458), .B1(new_n463), .B2(new_n404), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n453), .A2(new_n458), .B1(new_n450), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n466));
  NOR2_X1   g280(.A1(G475), .A2(G902), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n465), .A2(KEYINPUT93), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n450), .A2(new_n464), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n403), .A2(G146), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n223), .B(new_n387), .C1(new_n402), .C2(new_n393), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n474), .A2(new_n420), .B1(new_n448), .B2(new_n449), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n470), .B(new_n471), .C1(new_n475), .C2(new_n424), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n476), .A2(new_n466), .B1(new_n465), .B2(new_n467), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n457), .B1(new_n469), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n207), .A2(KEYINPUT14), .A3(G122), .ZN(new_n479));
  XNOR2_X1  g293(.A(G116), .B(G122), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(G107), .B(new_n479), .C1(new_n481), .C2(KEYINPUT14), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n191), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT67), .B(G134), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n225), .A2(G128), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n243), .A2(G143), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n482), .B(new_n483), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n480), .B(new_n191), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n486), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n485), .A2(new_n492), .ZN(new_n495));
  OAI21_X1  g309(.A(G134), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n496), .A3(new_n487), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G217), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n382), .A2(new_n499), .A3(G953), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n498), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n302), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G478), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n505), .A3(G478), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(G234), .A2(G237), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(G952), .A3(new_n406), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(G902), .A3(G953), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NOR4_X1   g331(.A1(new_n320), .A2(new_n385), .A3(new_n478), .A4(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n406), .A2(G221), .A3(G234), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n519), .B(new_n520), .Z(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n243), .A2(G119), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT23), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G128), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G110), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n523), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT24), .B(G110), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(KEYINPUT74), .A3(new_n534), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n434), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(new_n473), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n529), .A2(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n399), .B2(new_n404), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n522), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n541), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n472), .B2(new_n473), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n404), .A2(new_n538), .A3(new_n434), .A4(new_n537), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n521), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n547), .A3(new_n302), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n543), .A2(new_n547), .A3(new_n302), .A4(new_n550), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n499), .B1(G234), .B2(new_n302), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(G902), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n543), .A2(new_n547), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G131), .B1(new_n335), .B2(new_n333), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n484), .B2(new_n333), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n343), .B1(new_n334), .B2(new_n484), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(new_n346), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n349), .A2(new_n250), .B1(new_n563), .B2(new_n246), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n256), .ZN(new_n565));
  INV_X1    g379(.A(new_n561), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n246), .A2(new_n348), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n354), .B2(new_n274), .ZN(new_n568));
  INV_X1    g382(.A(new_n256), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT71), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT28), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n232), .B(new_n236), .C1(new_n352), .C2(new_n353), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n256), .B1(new_n574), .B2(new_n567), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n575), .B2(KEYINPUT71), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n572), .A2(new_n576), .B1(new_n573), .B2(new_n565), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n411), .A2(G210), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT27), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT26), .B(G101), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT70), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT29), .B1(new_n577), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n574), .A2(new_n256), .A3(new_n567), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT64), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT30), .B1(new_n568), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT30), .ZN(new_n590));
  AOI211_X1 g404(.A(KEYINPUT64), .B(new_n590), .C1(new_n574), .C2(new_n567), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n569), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT68), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n590), .B1(new_n564), .B2(KEYINPUT64), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n568), .A2(new_n588), .A3(KEYINPUT30), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT68), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n569), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n587), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n582), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n586), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n565), .A2(new_n570), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT28), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n565), .A2(new_n573), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT29), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n582), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n587), .A2(new_n582), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n597), .B1(new_n596), .B2(new_n569), .ZN(new_n613));
  AOI211_X1 g427(.A(KEYINPUT68), .B(new_n256), .C1(new_n594), .C2(new_n595), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n577), .A2(new_n585), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT31), .ZN(new_n617));
  INV_X1    g431(.A(new_n611), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n593), .B2(new_n598), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(G472), .A2(G902), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT32), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n610), .A2(G472), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n621), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n623), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n559), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n518), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT96), .B(G101), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G3));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n620), .A2(new_n302), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n626), .ZN(new_n635));
  INV_X1    g449(.A(new_n559), .ZN(new_n636));
  INV_X1    g450(.A(new_n383), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n375), .A2(new_n367), .B1(new_n377), .B2(new_n372), .ZN(new_n638));
  OAI21_X1  g452(.A(G469), .B1(new_n638), .B2(G902), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n637), .B1(new_n639), .B2(new_n374), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n632), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n381), .A2(new_n383), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n559), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n644), .A2(KEYINPUT97), .A3(new_n626), .A4(new_n634), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n502), .B(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G478), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(G902), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT98), .B(G478), .Z(new_n652));
  OAI22_X1  g466(.A1(new_n648), .A2(new_n651), .B1(new_n504), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n478), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n384), .ZN(new_n655));
  INV_X1    g469(.A(new_n303), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n308), .B2(new_n313), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n655), .B1(new_n657), .B2(new_n304), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n654), .A2(new_n659), .A3(new_n516), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n646), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NAND2_X1  g477(.A1(new_n465), .A2(new_n467), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n466), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n467), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n457), .A2(new_n509), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n516), .B(KEYINPUT99), .Z(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n659), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  INV_X1    g487(.A(new_n555), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n552), .B2(new_n553), .ZN(new_n675));
  OAI22_X1  g489(.A1(new_n542), .A2(new_n540), .B1(KEYINPUT36), .B2(new_n522), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n545), .A2(new_n546), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n557), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n676), .A2(KEYINPUT100), .A3(new_n557), .A4(new_n678), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n635), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n518), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  NAND2_X1  g502(.A1(new_n620), .A2(new_n624), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n587), .A2(new_n575), .A3(KEYINPUT71), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT28), .B1(new_n570), .B2(new_n571), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n604), .B(new_n585), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n607), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n565), .B1(new_n613), .B2(new_n614), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n693), .B1(new_n694), .B2(new_n582), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n606), .A2(new_n608), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n302), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n577), .A2(new_n585), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n699), .B1(new_n700), .B2(KEYINPUT31), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n622), .B1(new_n701), .B2(new_n615), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n689), .B(new_n698), .C1(new_n702), .C2(KEYINPUT32), .ZN(new_n703));
  INV_X1    g517(.A(new_n684), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n514), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n511), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n667), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n657), .A2(new_n304), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n381), .A2(new_n710), .A3(new_n383), .A4(new_n384), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n703), .A2(new_n704), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n684), .B1(new_n625), .B2(new_n627), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(KEYINPUT101), .A3(new_n709), .A4(new_n711), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n602), .A2(new_n584), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n302), .B1(new_n722), .B2(new_n619), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G472), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n689), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT32), .B1(new_n620), .B2(new_n621), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n719), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n627), .A2(KEYINPUT103), .A3(new_n689), .A4(new_n724), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n509), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n476), .A2(new_n466), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n664), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n468), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n731), .B1(new_n734), .B2(new_n457), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n384), .A3(new_n684), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n707), .B(KEYINPUT39), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n643), .A2(KEYINPUT40), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT40), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n640), .B2(new_n737), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n736), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n319), .A2(KEYINPUT38), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n319), .A2(KEYINPUT38), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n730), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G143), .ZN(G45));
  AND3_X1   g561(.A1(new_n478), .A2(new_n653), .A3(new_n707), .ZN(new_n748));
  AND4_X1   g562(.A1(new_n703), .A2(new_n748), .A3(new_n704), .A4(new_n711), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n223), .ZN(G48));
  INV_X1    g564(.A(new_n363), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n331), .A2(new_n357), .B1(new_n361), .B2(new_n204), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n354), .B1(new_n752), .B2(new_n360), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n367), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n363), .B(new_n368), .C1(new_n350), .C2(new_n355), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n380), .B1(new_n756), .B2(new_n302), .ZN(new_n757));
  INV_X1    g571(.A(new_n321), .ZN(new_n758));
  AOI211_X1 g572(.A(G902), .B(new_n758), .C1(new_n754), .C2(new_n755), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n383), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n628), .A2(new_n660), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT41), .B(G113), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G15));
  NAND3_X1  g579(.A1(new_n628), .A2(new_n670), .A3(new_n762), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G116), .ZN(G18));
  NAND3_X1  g581(.A1(new_n658), .A2(new_n760), .A3(new_n383), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n478), .A3(new_n517), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n715), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G119), .ZN(G21));
  NAND2_X1  g585(.A1(new_n605), .A2(new_n584), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n619), .B2(new_n617), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT104), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n773), .A2(new_n774), .B1(new_n619), .B2(new_n612), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT104), .B(new_n772), .C1(new_n619), .C2(new_n617), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n622), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(G472), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n620), .B2(new_n302), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n777), .A2(new_n559), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n478), .A2(new_n658), .A3(new_n509), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n761), .A3(new_n669), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G122), .ZN(G24));
  NOR4_X1   g598(.A1(new_n777), .A2(new_n768), .A3(new_n779), .A4(new_n684), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n478), .A2(new_n653), .A3(new_n707), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT105), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT105), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n478), .A2(new_n788), .A3(new_n653), .A4(new_n707), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G125), .ZN(G27));
  NOR2_X1   g606(.A1(new_n385), .A2(new_n319), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n793), .A3(new_n789), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n698), .A2(new_n689), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT106), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n797), .B1(new_n798), .B2(new_n627), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n726), .A2(KEYINPUT106), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n559), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n628), .A2(new_n787), .A3(new_n789), .A4(new_n793), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n796), .A2(new_n801), .B1(new_n802), .B2(new_n795), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT107), .B(G131), .Z(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G33));
  NAND3_X1  g619(.A1(new_n628), .A2(new_n709), .A3(new_n793), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G134), .ZN(G36));
  NOR2_X1   g621(.A1(new_n380), .A2(new_n302), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n376), .A2(KEYINPUT45), .A3(new_n378), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT108), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n638), .A2(new_n811), .A3(KEYINPUT45), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n638), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n380), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n808), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n374), .B1(new_n817), .B2(KEYINPUT46), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n819), .B(new_n808), .C1(new_n813), .C2(new_n816), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n383), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n821), .A2(KEYINPUT109), .A3(new_n738), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT109), .B1(new_n821), .B2(new_n738), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n457), .B(new_n653), .C1(new_n469), .C2(new_n477), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT43), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT43), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n734), .A2(new_n826), .A3(new_n457), .A4(new_n653), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n635), .A2(new_n704), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT44), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n305), .A2(new_n314), .A3(new_n318), .A4(new_n384), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n828), .B2(KEYINPUT44), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n822), .A2(new_n823), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G137), .ZN(G39));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n821), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(KEYINPUT47), .B(new_n383), .C1(new_n818), .C2(new_n820), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n830), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n703), .A2(new_n636), .A3(new_n786), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G140), .ZN(G42));
  NOR3_X1   g655(.A1(new_n675), .A2(new_n683), .A3(new_n708), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n735), .A2(new_n842), .A3(new_n640), .A4(new_n658), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n727), .B2(new_n728), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n749), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n717), .A3(new_n791), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT113), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n717), .A2(new_n791), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n714), .A2(new_n716), .B1(new_n785), .B2(new_n790), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT112), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n844), .A2(new_n749), .A3(new_n847), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT52), .B1(new_n853), .B2(new_n845), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n849), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n783), .A2(new_n763), .A3(new_n766), .A4(new_n770), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n803), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n509), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n507), .A2(KEYINPUT111), .A3(new_n508), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n654), .B1(new_n866), .B2(new_n478), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n320), .A2(new_n655), .A3(new_n669), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n642), .A2(new_n645), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n518), .B1(new_n685), .B2(new_n628), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n707), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n457), .A2(new_n665), .A3(new_n666), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n684), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n703), .A3(new_n640), .A4(new_n838), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n777), .A2(new_n779), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n704), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n806), .B(new_n875), .C1(new_n877), .C2(new_n794), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n862), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n860), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n846), .A2(new_n847), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n862), .B(new_n879), .C1(new_n883), .C2(new_n857), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT53), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(KEYINPUT54), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n796), .A2(new_n801), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n802), .A2(new_n795), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n861), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT114), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n871), .A2(new_n878), .A3(new_n880), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT114), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n803), .B2(new_n861), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n860), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n884), .A2(new_n880), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n825), .A2(new_n512), .A3(new_n827), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT115), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n825), .A2(new_n827), .A3(new_n902), .A4(new_n512), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n762), .A2(new_n838), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT118), .B1(new_n761), .B2(new_n830), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n904), .A2(new_n704), .A3(new_n876), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n559), .A2(new_n511), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n478), .A2(new_n653), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n729), .A2(new_n908), .A3(new_n910), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(KEYINPUT50), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n775), .A2(new_n776), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n621), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n636), .A3(new_n634), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n901), .B2(new_n903), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n761), .A2(new_n384), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n743), .A2(new_n922), .A3(new_n744), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n917), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n914), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n904), .A2(KEYINPUT116), .A3(new_n923), .A4(new_n780), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n916), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT50), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n921), .A2(new_n838), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n760), .A2(new_n637), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n835), .A2(new_n836), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n925), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT51), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n835), .A2(KEYINPUT119), .A3(new_n836), .A4(new_n931), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n939), .A3(new_n930), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n940), .A2(KEYINPUT51), .A3(new_n929), .A4(new_n925), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n921), .A2(new_n658), .A3(new_n762), .ZN(new_n942));
  INV_X1    g756(.A(new_n654), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n729), .A2(new_n908), .A3(new_n943), .A4(new_n910), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n942), .A2(G952), .A3(new_n944), .A4(new_n406), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n801), .A2(new_n904), .A3(new_n908), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT48), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(KEYINPUT48), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n936), .A2(new_n941), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n886), .A2(new_n899), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(G952), .A2(G953), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n730), .A2(new_n745), .ZN(new_n954));
  NOR4_X1   g768(.A1(new_n824), .A2(new_n559), .A3(new_n637), .A4(new_n655), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(KEYINPUT110), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(KEYINPUT110), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n760), .B(KEYINPUT49), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n954), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n953), .A2(KEYINPUT120), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G75));
  INV_X1    g779(.A(KEYINPUT122), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n406), .A2(G952), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT121), .Z(new_n968));
  AOI22_X1  g782(.A1(new_n860), .A2(new_n895), .B1(new_n884), .B2(new_n880), .ZN(new_n969));
  INV_X1    g783(.A(new_n306), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n302), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n295), .A2(new_n300), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n313), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT55), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT56), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n968), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n896), .A2(new_n898), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(G210), .A3(G902), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n979), .B2(new_n975), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n966), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n968), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n978), .A2(G902), .A3(new_n306), .ZN(new_n983));
  INV_X1    g797(.A(new_n976), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n969), .A2(new_n302), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT56), .B1(new_n986), .B2(G210), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n985), .B(KEYINPUT122), .C1(new_n987), .C2(new_n974), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n981), .A2(new_n988), .ZN(G51));
  NAND3_X1  g803(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n990));
  AOI211_X1 g804(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n853), .C2(new_n845), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n858), .B1(new_n846), .B2(new_n847), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n990), .B1(new_n993), .B2(new_n856), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n846), .B(new_n847), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n862), .A2(new_n879), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT53), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT54), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(KEYINPUT123), .A3(new_n899), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT123), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n978), .A2(new_n1000), .A3(KEYINPUT54), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n808), .B(KEYINPUT57), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n756), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n986), .A2(new_n813), .A3(new_n816), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n967), .B1(new_n1004), .B2(new_n1005), .ZN(G54));
  NAND3_X1  g820(.A1(new_n986), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1007));
  INV_X1    g821(.A(new_n465), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1009), .A2(new_n1010), .A3(new_n967), .ZN(G60));
  NAND2_X1  g825(.A1(G478), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT59), .Z(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n886), .B2(new_n899), .ZN(new_n1014));
  INV_X1    g828(.A(new_n648), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n968), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n648), .A2(new_n1013), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n999), .A2(new_n1001), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT124), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT124), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n999), .A2(new_n1020), .A3(new_n1001), .A4(new_n1017), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1016), .B1(new_n1019), .B2(new_n1021), .ZN(G63));
  NAND2_X1  g836(.A1(G217), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT60), .Z(new_n1024));
  NAND2_X1  g838(.A1(new_n978), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n543), .A2(new_n547), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n978), .A2(new_n678), .A3(new_n676), .A4(new_n1024), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1027), .A2(new_n968), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT61), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1027), .A2(KEYINPUT61), .A3(new_n968), .A4(new_n1028), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(G66));
  OAI21_X1  g847(.A(G953), .B1(new_n515), .B2(new_n252), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n871), .A2(new_n861), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(G953), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n312), .B(new_n291), .C1(G898), .C2(new_n406), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(G69));
  OAI21_X1  g852(.A(G953), .B1(new_n365), .B2(new_n705), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1039), .B(KEYINPUT127), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  AND2_X1   g855(.A1(new_n628), .A2(new_n793), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n803), .B1(new_n709), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n822), .A2(new_n823), .ZN(new_n1044));
  INV_X1    g858(.A(new_n781), .ZN(new_n1045));
  AOI22_X1  g859(.A1(new_n829), .A2(new_n831), .B1(new_n1045), .B2(new_n801), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1043), .B(new_n840), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g861(.A(new_n749), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n852), .A2(new_n1048), .A3(new_n854), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n406), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n705), .A2(G953), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT126), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g868(.A(KEYINPUT126), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1055));
  XNOR2_X1  g869(.A(new_n596), .B(new_n461), .ZN(new_n1056));
  NOR3_X1   g870(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1056), .A2(new_n406), .ZN(new_n1058));
  NAND4_X1  g872(.A1(new_n852), .A2(new_n746), .A3(new_n854), .A4(new_n1048), .ZN(new_n1059));
  INV_X1    g873(.A(KEYINPUT62), .ZN(new_n1060));
  XNOR2_X1  g874(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1042), .A2(new_n737), .A3(new_n867), .ZN(new_n1062));
  AND3_X1   g876(.A1(new_n832), .A2(new_n840), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g878(.A(KEYINPUT125), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n1061), .A2(KEYINPUT125), .A3(new_n1063), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1058), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n1041), .B1(new_n1057), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g883(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1070));
  OAI21_X1  g884(.A(new_n1070), .B1(new_n1053), .B2(new_n1052), .ZN(new_n1071));
  AND3_X1   g885(.A1(new_n1061), .A2(KEYINPUT125), .A3(new_n1063), .ZN(new_n1072));
  AOI21_X1  g886(.A(KEYINPUT125), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1073));
  OAI211_X1 g887(.A(new_n406), .B(new_n1056), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g888(.A1(new_n1071), .A2(new_n1074), .A3(new_n1040), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1069), .A2(new_n1075), .ZN(G72));
  NOR4_X1   g890(.A1(new_n1047), .A2(new_n861), .A3(new_n871), .A4(new_n1049), .ZN(new_n1077));
  NAND2_X1  g891(.A1(G472), .A2(G902), .ZN(new_n1078));
  XOR2_X1   g892(.A(new_n1078), .B(KEYINPUT63), .Z(new_n1079));
  INV_X1    g893(.A(new_n1079), .ZN(new_n1080));
  OAI211_X1 g894(.A(new_n582), .B(new_n599), .C1(new_n1077), .C2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g895(.A(new_n700), .B1(new_n599), .B2(new_n600), .ZN(new_n1082));
  NAND4_X1  g896(.A1(new_n882), .A2(new_n885), .A3(new_n1079), .A4(new_n1082), .ZN(new_n1083));
  OAI211_X1 g897(.A(new_n1081), .B(new_n1083), .C1(G952), .C2(new_n406), .ZN(new_n1084));
  NAND3_X1  g898(.A1(new_n1066), .A2(new_n1035), .A3(new_n1067), .ZN(new_n1085));
  NAND2_X1  g899(.A1(new_n1085), .A2(new_n1079), .ZN(new_n1086));
  NOR2_X1   g900(.A1(new_n599), .A2(new_n582), .ZN(new_n1087));
  AOI21_X1  g901(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(G57));
endmodule


