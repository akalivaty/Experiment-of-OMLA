//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT75), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  OAI21_X1  g006(.A(G214), .B1(G237), .B2(G902), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT77), .B1(new_n195), .B2(G104), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G107), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n195), .A2(KEYINPUT3), .A3(G104), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT3), .B1(new_n195), .B2(G104), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n196), .B(new_n199), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n198), .B2(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n195), .A2(KEYINPUT3), .A3(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n207), .A2(new_n208), .A3(new_n196), .A4(new_n199), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G116), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT2), .B(G113), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n202), .A2(new_n218), .A3(G101), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n215), .A2(new_n216), .ZN(new_n221));
  INV_X1    g035(.A(G113), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n212), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n212), .A3(new_n214), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n221), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n231));
  XNOR2_X1  g045(.A(G104), .B(G107), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n208), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n195), .A2(G104), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n198), .A2(G107), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT78), .A3(G101), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n230), .A2(new_n209), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n220), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n220), .A2(new_n239), .A3(new_n241), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(KEYINPUT6), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT6), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n246), .A3(new_n242), .ZN(new_n247));
  XNOR2_X1  g061(.A(G143), .B(G146), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT64), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n251), .A3(G146), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n249), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n250), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G125), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT1), .ZN(new_n264));
  INV_X1    g078(.A(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G143), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n266), .A3(new_n253), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n248), .A2(KEYINPUT68), .A3(new_n264), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n255), .B1(new_n251), .B2(G146), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n265), .A2(KEYINPUT64), .A3(G143), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n262), .B1(G125), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G224), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G953), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n245), .A2(new_n247), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n245), .A2(KEYINPUT83), .A3(new_n247), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT8), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n241), .B(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT78), .B1(new_n236), .B2(G101), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n231), .B(new_n208), .C1(new_n234), .C2(new_n235), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n209), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n292), .B2(new_n230), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT84), .ZN(new_n294));
  OAI21_X1  g108(.A(G113), .B1(new_n228), .B2(new_n212), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT5), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n209), .B(new_n238), .C1(new_n297), .C2(new_n221), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n293), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n294), .B1(new_n293), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT7), .B1(new_n280), .B2(G953), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n279), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n302), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n262), .B(new_n304), .C1(G125), .C2(new_n278), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n244), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n190), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT85), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(KEYINPUT85), .B(new_n190), .C1(new_n301), .C2(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n287), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G210), .B1(G237), .B2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n287), .A2(new_n311), .A3(new_n313), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n194), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n275), .A2(G128), .B1(new_n266), .B2(new_n253), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n269), .B2(new_n270), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT79), .B1(new_n292), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n266), .A2(new_n253), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n276), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT68), .B1(new_n248), .B2(new_n264), .ZN(new_n323));
  AND4_X1   g137(.A1(KEYINPUT68), .A2(new_n264), .A3(new_n266), .A4(new_n253), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n209), .A4(new_n238), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n278), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n292), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT11), .ZN(new_n332));
  INV_X1    g146(.A(G134), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(G137), .ZN(new_n334));
  INV_X1    g148(.A(G137), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT11), .A3(G134), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(G137), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G131), .ZN(new_n339));
  INV_X1    g153(.A(G131), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n334), .A2(new_n336), .A3(new_n340), .A4(new_n337), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT12), .B1(new_n342), .B2(KEYINPUT80), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n331), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n320), .A2(new_n327), .B1(new_n329), .B2(new_n292), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n339), .A2(new_n341), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n328), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n274), .A2(new_n259), .B1(new_n248), .B2(new_n249), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n210), .A2(new_n352), .A3(new_n219), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n278), .A2(KEYINPUT10), .A3(new_n209), .A4(new_n238), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n355), .A3(new_n347), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G953), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G227), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT76), .ZN(new_n360));
  XNOR2_X1  g174(.A(G110), .B(G140), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT10), .B1(new_n320), .B2(new_n327), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n353), .A2(new_n354), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n364), .A2(new_n365), .A3(new_n342), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(new_n363), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n342), .B1(new_n364), .B2(new_n365), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n357), .A2(new_n363), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G469), .B1(new_n369), .B2(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n356), .A2(new_n368), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n367), .A2(new_n349), .B1(new_n371), .B2(new_n363), .ZN(new_n372));
  NOR4_X1   g186(.A1(new_n372), .A2(KEYINPUT81), .A3(G469), .A4(G902), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n344), .B1(new_n331), .B2(new_n342), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n346), .A2(new_n347), .A3(new_n343), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n356), .B(new_n362), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n347), .B1(new_n351), .B2(new_n355), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n363), .B1(new_n378), .B2(new_n366), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G469), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n370), .B1(new_n373), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G475), .ZN(new_n384));
  XNOR2_X1  g198(.A(G113), .B(G122), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n198), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n358), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n251), .A2(KEYINPUT86), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G143), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(G237), .A2(G953), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n393), .A2(G214), .B1(new_n390), .B2(G143), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT18), .B(G131), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT87), .B1(new_n396), .B2(new_n265), .ZN(new_n397));
  INV_X1    g211(.A(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G125), .ZN(new_n399));
  INV_X1    g213(.A(G125), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G146), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n388), .A2(new_n391), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT86), .B(G143), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n405), .B(new_n406), .C1(new_n388), .C2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(KEYINPUT87), .A3(G146), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n395), .A2(new_n404), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n392), .B2(new_n394), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT17), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n405), .B(new_n340), .C1(new_n388), .C2(new_n407), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT17), .B(G131), .C1(new_n392), .C2(new_n394), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT16), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n398), .A3(G125), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n402), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n265), .ZN(new_n419));
  OAI211_X1 g233(.A(G146), .B(new_n417), .C1(new_n402), .C2(new_n416), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n386), .B(new_n410), .C1(new_n414), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT88), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n424), .A2(new_n419), .A3(new_n420), .A4(new_n415), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n386), .A4(new_n410), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n425), .A2(new_n410), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n386), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n384), .B1(new_n430), .B2(new_n190), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(G475), .A2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n411), .A2(new_n413), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n402), .B(KEYINPUT19), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(G146), .B2(new_n436), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n420), .A2(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n420), .A2(KEYINPUT72), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n410), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n386), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n434), .B1(new_n428), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n428), .A2(new_n443), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT89), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n445), .A2(new_n449), .A3(new_n447), .A4(new_n433), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n432), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G116), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n195), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n251), .A2(G128), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT13), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n263), .A2(G143), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n455), .A2(new_n456), .ZN(new_n460));
  OAI21_X1  g274(.A(G134), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n458), .A3(new_n333), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n454), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n189), .A2(G217), .A3(new_n358), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n213), .A2(G122), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(KEYINPUT14), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n213), .A2(G122), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n468), .B2(KEYINPUT14), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n469), .B2(KEYINPUT90), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(KEYINPUT90), .B2(new_n469), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n471), .A2(G107), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n453), .A2(new_n195), .ZN(new_n473));
  INV_X1    g287(.A(new_n462), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n333), .B1(new_n455), .B2(new_n458), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n463), .B(new_n465), .C1(new_n472), .C2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n471), .B2(G107), .ZN(new_n478));
  INV_X1    g292(.A(new_n463), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n464), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n481), .A2(new_n190), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n481), .B2(new_n190), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G952), .ZN(new_n488));
  AOI211_X1 g302(.A(G953), .B(new_n488), .C1(G234), .C2(G237), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n190), .B(new_n358), .C1(G234), .C2(G237), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT21), .B(G898), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n452), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  AND4_X1   g307(.A1(new_n192), .A2(new_n317), .A3(new_n383), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n263), .A2(G119), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n211), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT24), .B(G110), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n419), .A2(new_n420), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT23), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n211), .B2(G128), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n263), .A2(KEYINPUT23), .A3(G119), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n503), .A2(new_n504), .A3(new_n496), .ZN(new_n505));
  INV_X1    g319(.A(G110), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n497), .A2(new_n498), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n509), .A2(new_n510), .B1(new_n265), .B2(new_n396), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n439), .A3(new_n438), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT22), .B(G137), .Z(new_n515));
  AND3_X1   g329(.A1(new_n358), .A2(G221), .A3(G234), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n513), .B1(new_n508), .B2(new_n512), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n513), .B(new_n518), .C1(new_n508), .C2(new_n512), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(KEYINPUT74), .B(KEYINPUT25), .C1(new_n523), .C2(G902), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n508), .A2(new_n512), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n514), .A3(new_n518), .ZN(new_n528));
  INV_X1    g342(.A(new_n522), .ZN(new_n529));
  AOI21_X1  g343(.A(G902), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G217), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(G234), .B2(new_n190), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n524), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(G902), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n521), .B2(new_n522), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n341), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n335), .A2(G134), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n340), .B1(new_n540), .B2(new_n337), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n541), .A2(KEYINPUT66), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT66), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n543), .B(new_n340), .C1(new_n540), .C2(new_n337), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n539), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n546), .A2(new_n278), .B1(new_n352), .B2(new_n342), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT30), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n541), .A2(KEYINPUT66), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n341), .B1(new_n549), .B2(new_n544), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n550), .A2(KEYINPUT67), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n550), .A2(KEYINPUT67), .B1(new_n271), .B2(new_n277), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT65), .B1(new_n347), .B2(new_n261), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT65), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n352), .A2(new_n554), .A3(new_n342), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n217), .B(new_n548), .C1(new_n556), .C2(KEYINPUT30), .ZN(new_n557));
  INV_X1    g371(.A(new_n217), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n393), .A2(G210), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT27), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(G101), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n557), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT31), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n559), .A2(KEYINPUT28), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT28), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n547), .B2(new_n558), .ZN(new_n568));
  OAI22_X1  g382(.A1(new_n566), .A2(new_n568), .B1(new_n558), .B2(new_n556), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n563), .B(KEYINPUT70), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n572));
  NAND4_X1  g386(.A1(new_n557), .A2(new_n559), .A3(new_n563), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n565), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(G472), .A2(G902), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT32), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT32), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n547), .A2(new_n558), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n566), .B2(new_n568), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n563), .A2(KEYINPUT29), .ZN(new_n585));
  AOI21_X1  g399(.A(G902), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n557), .A2(new_n559), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n563), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n569), .B2(new_n570), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n538), .B1(new_n580), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n494), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n574), .A2(new_n596), .A3(new_n190), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n574), .B2(new_n190), .ZN(new_n598));
  INV_X1    g412(.A(G472), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n600), .A2(KEYINPUT92), .B1(new_n575), .B2(new_n574), .ZN(new_n601));
  OR3_X1    g415(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n538), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n383), .A2(new_n605), .A3(new_n192), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n601), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT93), .ZN(new_n608));
  INV_X1    g422(.A(new_n492), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n287), .A2(new_n311), .A3(new_n313), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n313), .B1(new_n287), .B2(new_n311), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n193), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n449), .B1(new_n428), .B2(new_n443), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n423), .A2(new_n427), .B1(new_n442), .B2(new_n441), .ZN(new_n614));
  OAI22_X1  g428(.A1(new_n613), .A2(KEYINPUT20), .B1(new_n614), .B2(new_n434), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n431), .B1(new_n615), .B2(new_n450), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n481), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n481), .A2(new_n617), .A3(KEYINPUT33), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n482), .A2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n481), .A2(new_n190), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n622), .A2(new_n623), .B1(new_n482), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n616), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n612), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n608), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  XNOR2_X1  g445(.A(new_n444), .B(KEYINPUT20), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n431), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n487), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n612), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n608), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n518), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n526), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n536), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n535), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n494), .A2(new_n601), .A3(new_n604), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  AND3_X1   g459(.A1(new_n574), .A2(new_n578), .A3(new_n575), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n578), .B1(new_n574), .B2(new_n575), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n592), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n642), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n317), .A2(new_n192), .A3(new_n383), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n490), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n489), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n634), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT95), .B(G128), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G30));
  NAND2_X1  g474(.A1(new_n377), .A2(new_n379), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n381), .A3(new_n190), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT81), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n380), .A2(new_n374), .A3(new_n381), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n191), .B1(new_n665), .B2(new_n370), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n655), .B(KEYINPUT39), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT40), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n582), .A2(new_n559), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n587), .A2(new_n563), .B1(new_n570), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(G902), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n642), .B1(new_n580), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n610), .A2(new_n611), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n452), .A2(new_n487), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n674), .A2(new_n676), .A3(new_n194), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n669), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  INV_X1    g494(.A(KEYINPUT96), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n626), .B2(new_n655), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n616), .A2(new_n625), .A3(KEYINPUT96), .A4(new_n656), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n642), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n580), .B2(new_n592), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n684), .A2(new_n686), .A3(new_n666), .A4(new_n317), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  OAI21_X1  g502(.A(G469), .B1(new_n380), .B2(KEYINPUT97), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT97), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n372), .A2(new_n690), .A3(G902), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT98), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n380), .A2(KEYINPUT97), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n690), .B1(new_n372), .B2(G902), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT98), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .A4(G469), .ZN(new_n696));
  AND4_X1   g510(.A1(new_n192), .A2(new_n692), .A3(new_n665), .A4(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n648), .A2(new_n605), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n628), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n635), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NAND4_X1  g519(.A1(new_n697), .A2(new_n686), .A3(new_n317), .A4(new_n493), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  NAND2_X1  g521(.A1(new_n583), .A2(KEYINPUT99), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT99), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n709), .B(new_n582), .C1(new_n566), .C2(new_n568), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n570), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n565), .A3(new_n573), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n575), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n599), .B1(new_n574), .B2(new_n190), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI211_X1 g530(.A(KEYINPUT100), .B(new_n599), .C1(new_n574), .C2(new_n190), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n538), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n193), .B1(new_n610), .B2(new_n611), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n719), .A2(new_n492), .A3(new_n677), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n697), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR3_X1   g536(.A1(new_n716), .A2(new_n685), .A3(new_n717), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n697), .A3(new_n684), .A4(new_n317), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND2_X1  g540(.A1(G469), .A2(G902), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT101), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n369), .B2(G469), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n191), .B1(new_n665), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n610), .A2(new_n611), .A3(new_n194), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n726), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n729), .B1(new_n373), .B2(new_n382), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n726), .A2(new_n731), .A3(new_n192), .A4(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n593), .B(new_n684), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n731), .A2(new_n192), .A3(new_n733), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT102), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n730), .A2(new_n726), .A3(new_n731), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n699), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT42), .B1(new_n741), .B2(new_n684), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT103), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n735), .A2(new_n736), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(KEYINPUT42), .A3(new_n684), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  OAI211_X1 g563(.A(new_n593), .B(new_n657), .C1(new_n732), .C2(new_n734), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND2_X1  g565(.A1(new_n622), .A2(new_n623), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n624), .A2(new_n482), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n616), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT43), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n685), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n576), .B1(new_n602), .B2(new_n603), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n600), .A2(KEYINPUT92), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n757), .B(KEYINPUT44), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT104), .Z(new_n761));
  NAND2_X1  g575(.A1(new_n601), .A2(new_n604), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT44), .B1(new_n762), .B2(new_n757), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n367), .A2(new_n368), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n366), .B1(new_n345), .B2(new_n348), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n765), .B2(new_n362), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n381), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  INV_X1    g583(.A(new_n728), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n665), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n192), .B(new_n667), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n731), .B(KEYINPUT105), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n763), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n761), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  OAI21_X1  g595(.A(new_n192), .B1(new_n774), .B2(new_n775), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT47), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n452), .A2(new_n754), .A3(new_n655), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n626), .A2(new_n681), .A3(new_n655), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n731), .ZN(new_n788));
  OR4_X1    g602(.A1(new_n648), .A2(new_n787), .A3(new_n788), .A4(new_n605), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n398), .ZN(G42));
  AND2_X1   g605(.A1(new_n665), .A2(new_n696), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n692), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT106), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n580), .A2(new_n672), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n538), .A2(new_n755), .A3(new_n191), .A4(new_n194), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n676), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n797), .B(new_n800), .C1(new_n795), .C2(new_n794), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n574), .A2(new_n190), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(G472), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT100), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n714), .A2(new_n715), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n642), .A3(new_n806), .A4(new_n713), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n787), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n734), .B2(new_n732), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n487), .A2(new_n656), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n666), .A2(new_n633), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n686), .A3(new_n731), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n750), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n452), .A2(new_n486), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n626), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n612), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n601), .A2(new_n604), .A3(new_n816), .A4(new_n606), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n643), .A2(new_n817), .A3(new_n594), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n697), .B(new_n593), .C1(new_n628), .C2(new_n635), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n706), .A3(new_n721), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n813), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n723), .A2(new_n684), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n792), .A2(new_n192), .A3(new_n317), .A4(new_n692), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n666), .A2(new_n648), .A3(new_n317), .A4(new_n642), .ZN(new_n824));
  INV_X1    g638(.A(new_n657), .ZN(new_n825));
  OAI22_X1  g639(.A1(new_n822), .A2(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n719), .A2(new_n677), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n673), .A2(new_n655), .A3(new_n827), .A4(new_n730), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n687), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT107), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(KEYINPUT108), .B(KEYINPUT52), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT107), .B(new_n831), .C1(new_n826), .C2(new_n829), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n748), .A2(new_n802), .A3(new_n821), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n826), .B2(new_n829), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n733), .A2(new_n192), .A3(new_n655), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n616), .A2(new_n486), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n840), .B(new_n193), .C1(new_n611), .C2(new_n610), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n651), .A2(new_n684), .B1(new_n842), .B2(new_n673), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n658), .A4(new_n724), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n821), .A2(new_n743), .A3(new_n845), .A4(new_n747), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n820), .A2(KEYINPUT109), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT109), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n819), .A2(new_n706), .A3(new_n721), .A4(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n849), .B(new_n851), .C1(new_n737), .C2(new_n742), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT110), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n813), .A2(new_n818), .A3(new_n802), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n744), .A2(new_n746), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT110), .A3(new_n851), .A4(new_n849), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n854), .A2(new_n835), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n846), .A2(new_n802), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n848), .B1(KEYINPUT54), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n698), .A2(new_n788), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n756), .A2(new_n654), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n593), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT48), .Z(new_n865));
  NAND2_X1  g679(.A1(new_n358), .A2(G952), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n718), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n823), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n605), .A2(new_n862), .A3(new_n489), .A4(new_n798), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n866), .B(new_n868), .C1(new_n626), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n616), .A3(new_n625), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT113), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n783), .B1(new_n192), .B2(new_n793), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n718), .A3(new_n777), .A4(new_n863), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n862), .A2(new_n723), .A3(new_n863), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n676), .A2(new_n194), .A3(new_n697), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT111), .B1(new_n867), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT50), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT51), .ZN(new_n882));
  OAI221_X1 g696(.A(new_n872), .B1(new_n871), .B2(new_n870), .C1(new_n878), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n881), .A2(KEYINPUT112), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n881), .A2(KEYINPUT112), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n878), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n861), .B(new_n883), .C1(new_n884), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n801), .B1(new_n888), .B2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n358), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n190), .B1(new_n858), .B2(new_n859), .ZN(new_n893));
  AOI211_X1 g707(.A(KEYINPUT116), .B(KEYINPUT56), .C1(new_n893), .C2(G210), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n245), .A2(new_n247), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT115), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n282), .B(KEYINPUT55), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n892), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n898), .B2(new_n894), .ZN(G51));
  XOR2_X1   g714(.A(new_n769), .B(KEYINPUT120), .Z(new_n901));
  AND2_X1   g715(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n728), .B(KEYINPUT57), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n858), .A2(new_n859), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n904), .B1(new_n858), .B2(new_n859), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n661), .B(KEYINPUT118), .ZN(new_n910));
  OAI211_X1 g724(.A(KEYINPUT117), .B(new_n903), .C1(new_n905), .C2(new_n906), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n902), .B1(new_n912), .B2(KEYINPUT119), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n909), .A2(new_n914), .A3(new_n910), .A4(new_n911), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n891), .B1(new_n913), .B2(new_n915), .ZN(G54));
  AND3_X1   g730(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n892), .B1(new_n917), .B2(new_n445), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n445), .B2(new_n917), .ZN(G60));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n861), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n622), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(KEYINPUT121), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n905), .A2(new_n906), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n622), .A2(new_n922), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n892), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT121), .B1(new_n923), .B2(new_n924), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT60), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n860), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n891), .B1(new_n933), .B2(new_n523), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n640), .B(KEYINPUT122), .Z(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g751(.A(G953), .B1(new_n491), .B2(new_n280), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n818), .A2(new_n820), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n896), .B1(G898), .B2(new_n358), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  INV_X1    g756(.A(new_n547), .ZN(new_n943));
  MUX2_X1   g757(.A(new_n556), .B(new_n943), .S(KEYINPUT30), .Z(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(new_n436), .Z(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n358), .B1(G227), .B2(G900), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n790), .B1(new_n761), .B2(new_n779), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n776), .A2(new_n699), .A3(new_n841), .ZN(new_n952));
  INV_X1    g766(.A(new_n687), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n826), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n748), .A2(new_n750), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n748), .A2(new_n958), .A3(new_n750), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n358), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n946), .B1(G900), .B2(G953), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n826), .A2(new_n953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n679), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  INV_X1    g780(.A(new_n815), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(KEYINPUT123), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n731), .B1(new_n967), .B2(KEYINPUT123), .ZN(new_n969));
  OR4_X1    g783(.A1(new_n699), .A2(new_n968), .A3(new_n969), .A4(new_n668), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n966), .A2(new_n951), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n945), .B1(new_n971), .B2(new_n358), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n950), .B1(new_n963), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n962), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n960), .B2(new_n358), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n976), .A2(KEYINPUT126), .A3(new_n972), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n949), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n963), .A2(new_n950), .A3(new_n973), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT126), .B1(new_n976), .B2(new_n972), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n979), .A2(new_n980), .A3(new_n947), .A4(new_n948), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(G72));
  INV_X1    g796(.A(new_n587), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n960), .A2(new_n939), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  AOI211_X1 g800(.A(new_n563), .B(new_n983), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n983), .A2(new_n563), .ZN(new_n988));
  INV_X1    g802(.A(new_n939), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n986), .B1(new_n971), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n992), .B(new_n986), .C1(new_n971), .C2(new_n989), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n988), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n587), .B(new_n563), .ZN(new_n995));
  AND4_X1   g809(.A1(new_n847), .A2(new_n836), .A3(new_n986), .A4(new_n995), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n987), .A2(new_n994), .A3(new_n891), .A4(new_n996), .ZN(G57));
endmodule


