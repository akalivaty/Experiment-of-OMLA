//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n191), .A2(new_n192), .A3(new_n195), .A4(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G137), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n204), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G137), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n197), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G131), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n205), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(KEYINPUT69), .A3(new_n205), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n193), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(new_n191), .B2(new_n192), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT0), .A3(G128), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n221), .A2(KEYINPUT65), .A3(new_n225), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n219), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n210), .B1(new_n217), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G116), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT68), .A3(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NOR3_X1   g055(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n243));
  INV_X1    g057(.A(G113), .ZN(new_n244));
  OAI22_X1  g058(.A1(new_n241), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n243), .A3(new_n244), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n240), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT2), .A2(G113), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n237), .A2(new_n249), .A3(new_n250), .A4(new_n238), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n231), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n231), .A2(KEYINPUT70), .A3(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n213), .ZN(new_n259));
  INV_X1    g073(.A(new_n219), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n221), .A2(KEYINPUT65), .A3(new_n225), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT65), .B1(new_n221), .B2(new_n225), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n259), .B1(new_n263), .B2(KEYINPUT66), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n230), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n210), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(new_n253), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT28), .B1(new_n258), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT28), .B1(new_n231), .B2(new_n253), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G237), .A2(G953), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G210), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n274), .B(KEYINPUT27), .Z(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G101), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n275), .B(new_n276), .Z(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT31), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n217), .A2(new_n230), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n209), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n282), .B(new_n252), .C1(new_n267), .C2(KEYINPUT30), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n283), .A2(new_n256), .A3(new_n257), .A4(new_n277), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n257), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT70), .B1(new_n231), .B2(new_n253), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n289), .A2(KEYINPUT71), .A3(new_n277), .A4(new_n283), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n280), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n284), .A2(new_n280), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n279), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(KEYINPUT32), .A3(new_n294), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n256), .B(new_n257), .C1(new_n253), .C2(new_n231), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n270), .B1(new_n299), .B2(KEYINPUT28), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n278), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(G902), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n289), .A2(new_n283), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n301), .B1(new_n304), .B2(new_n277), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n269), .A2(new_n271), .A3(new_n277), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G472), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n297), .A2(new_n298), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G125), .B(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT16), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G125), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n313), .A2(KEYINPUT16), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(G146), .A3(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n315), .A2(KEYINPUT74), .ZN(new_n316));
  INV_X1    g130(.A(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G146), .ZN(new_n320));
  INV_X1    g134(.A(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G119), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(KEYINPUT23), .A3(G119), .ZN(new_n325));
  INV_X1    g139(.A(G110), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n233), .A2(G128), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(new_n327), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT24), .B(G110), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n320), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n315), .A2(KEYINPUT74), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n316), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n316), .A2(new_n332), .A3(new_n333), .A4(KEYINPUT75), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n329), .A2(new_n330), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(G110), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n315), .ZN(new_n342));
  AOI21_X1  g156(.A(G146), .B1(new_n311), .B2(new_n314), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G953), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(G221), .A3(G234), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT76), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n353));
  INV_X1    g167(.A(G902), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n338), .A2(new_n344), .A3(new_n350), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT72), .B(G217), .Z(new_n357));
  INV_X1    g171(.A(G234), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(G902), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n359), .B(KEYINPUT73), .Z(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n350), .B1(new_n338), .B2(new_n344), .ZN(new_n363));
  INV_X1    g177(.A(new_n344), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n364), .B(new_n351), .C1(new_n336), .C2(new_n337), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n353), .B1(new_n366), .B2(new_n354), .ZN(new_n367));
  INV_X1    g181(.A(new_n366), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n361), .A2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI22_X1  g184(.A1(new_n362), .A2(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI221_X1 g187(.A(KEYINPUT77), .B1(new_n368), .B2(new_n370), .C1(new_n362), .C2(new_n367), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G214), .B1(G237), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT87), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n346), .A2(G224), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n228), .A2(new_n229), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n317), .B1(new_n380), .B2(new_n260), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n194), .A2(new_n317), .A3(new_n196), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT82), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n194), .A2(new_n384), .A3(new_n317), .A4(new_n196), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n379), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n385), .B(new_n383), .C1(new_n230), .C2(new_n317), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT85), .A3(new_n379), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n390), .B2(new_n379), .ZN(new_n394));
  INV_X1    g208(.A(new_n386), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n263), .A2(G125), .ZN(new_n396));
  INV_X1    g210(.A(new_n379), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n395), .A2(KEYINPUT86), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n401));
  AOI221_X4 g215(.A(new_n401), .B1(G116), .B2(new_n233), .C1(new_n234), .C2(new_n236), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n233), .A3(G116), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT79), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n405), .A2(new_n401), .A3(new_n233), .A4(G116), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(G113), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n251), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G104), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(new_n409), .B2(G107), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n411));
  INV_X1    g225(.A(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(G104), .ZN(new_n413));
  INV_X1    g227(.A(G101), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(G107), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n410), .A2(new_n413), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n409), .A2(G107), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n412), .A2(G104), .ZN(new_n418));
  OAI21_X1  g232(.A(G101), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT83), .B1(new_n408), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n237), .A2(KEYINPUT5), .A3(new_n238), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n422), .A2(G113), .A3(new_n406), .A4(new_n404), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n424));
  INV_X1    g238(.A(new_n420), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n251), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n408), .A2(new_n420), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n421), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT8), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n429), .B1(new_n428), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n377), .B1(new_n400), .B2(new_n434), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n389), .A2(new_n391), .B1(new_n394), .B2(new_n398), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n428), .A2(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT84), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(new_n440), .A3(KEYINPUT87), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n410), .A2(new_n413), .A3(new_n415), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G101), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT4), .A3(new_n416), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT4), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n445), .A3(G101), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n252), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n423), .A2(new_n251), .A3(new_n425), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n430), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n435), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G210), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n447), .A2(KEYINPUT80), .A3(new_n448), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT80), .B1(new_n447), .B2(new_n448), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(KEYINPUT6), .B(new_n455), .C1(new_n456), .C2(new_n457), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n449), .A3(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n390), .B(new_n378), .Z(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n450), .A2(new_n454), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n454), .B1(new_n450), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n376), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT99), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT95), .ZN(new_n469));
  INV_X1    g283(.A(G122), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT95), .A2(G122), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G116), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n412), .B1(new_n474), .B2(KEYINPUT14), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n470), .A2(G116), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n235), .B1(new_n471), .B2(new_n472), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n476), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n474), .B(new_n479), .C1(KEYINPUT14), .C2(new_n412), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n187), .A2(G128), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n321), .A2(G143), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT97), .ZN(new_n484));
  XNOR2_X1  g298(.A(G128), .B(G143), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT97), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n484), .A2(new_n487), .A3(new_n199), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(KEYINPUT97), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n486), .ZN(new_n490));
  AOI21_X1  g304(.A(G134), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n478), .B(new_n480), .C1(new_n488), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n485), .A2(KEYINPUT13), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n493), .B(G134), .C1(KEYINPUT13), .C2(new_n481), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT98), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT98), .B(G134), .C1(new_n489), .C2(new_n490), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT96), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n474), .A2(new_n499), .A3(new_n479), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT96), .B1(new_n477), .B2(new_n476), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n412), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n501), .A3(G107), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n492), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT9), .B(G234), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n346), .A3(new_n357), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n509), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n492), .B(new_n511), .C1(new_n498), .C2(new_n505), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI211_X1 g331(.A(G902), .B(new_n515), .C1(new_n510), .C2(new_n512), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n468), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n512), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n199), .B1(new_n484), .B2(new_n487), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT98), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n491), .A2(new_n495), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n524), .A2(new_n494), .A3(new_n504), .A4(new_n503), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n511), .B1(new_n525), .B2(new_n492), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n354), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n515), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n513), .A2(new_n516), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT99), .ZN(new_n530));
  NOR2_X1   g344(.A1(G475), .A2(G902), .ZN(new_n531));
  INV_X1    g345(.A(G237), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n346), .A3(G214), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(KEYINPUT89), .B2(new_n187), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT89), .B(G143), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G131), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n187), .A2(KEYINPUT89), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n187), .A2(KEYINPUT89), .ZN(new_n540));
  OAI211_X1 g354(.A(G214), .B(new_n273), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n203), .A3(new_n534), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n536), .A2(KEYINPUT17), .A3(G131), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT94), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n342), .A2(new_n343), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n203), .B1(new_n541), .B2(new_n534), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT17), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n543), .A2(new_n545), .A3(new_n546), .A4(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n551), .A2(KEYINPUT90), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n542), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(new_n547), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n541), .A2(new_n552), .A3(new_n534), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n319), .A2(G146), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n310), .A2(new_n190), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT91), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT91), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G113), .B(G122), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(new_n409), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT93), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n550), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n537), .A2(new_n542), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT19), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n319), .A2(KEYINPUT92), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n569), .A2(KEYINPUT92), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n569), .A2(KEYINPUT92), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n310), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n190), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n568), .A2(new_n316), .A3(new_n333), .A4(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n565), .B1(new_n563), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n531), .B1(new_n567), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT20), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n563), .A2(new_n575), .ZN(new_n579));
  INV_X1    g393(.A(new_n565), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n550), .A2(new_n563), .A3(new_n566), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n531), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n565), .B1(new_n550), .B2(new_n563), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n354), .B1(new_n567), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n578), .A2(new_n585), .B1(G475), .B2(new_n587), .ZN(new_n588));
  OR2_X1    g402(.A1(KEYINPUT100), .A2(G952), .ZN(new_n589));
  NAND2_X1  g403(.A1(KEYINPUT100), .A2(G952), .ZN(new_n590));
  AOI21_X1  g404(.A(G953), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n358), .B2(new_n532), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(G902), .B(G953), .C1(new_n358), .C2(new_n532), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT101), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT21), .B(G898), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n519), .A2(new_n530), .A3(new_n588), .A4(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G469), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n230), .A2(new_n444), .A3(new_n446), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n215), .A2(new_n216), .ZN(new_n603));
  INV_X1    g417(.A(new_n196), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n188), .A2(G128), .B1(new_n191), .B2(new_n192), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n416), .B(new_n419), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n425), .A2(new_n197), .A3(KEYINPUT10), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n602), .A2(new_n603), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(G110), .B(G140), .ZN(new_n611));
  INV_X1    g425(.A(G227), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(G953), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n611), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n420), .A2(new_n196), .A3(new_n194), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n606), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n217), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT78), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT12), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n215), .A2(new_n216), .B1(new_n617), .B2(new_n606), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT78), .B1(new_n623), .B2(KEYINPUT12), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n618), .A2(KEYINPUT12), .A3(new_n213), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n616), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n260), .B(new_n446), .C1(new_n261), .C2(new_n262), .ZN(new_n628));
  INV_X1    g442(.A(new_n444), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n608), .B(new_n609), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n217), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n615), .B1(new_n610), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n601), .B(new_n354), .C1(new_n627), .C2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n630), .A2(new_n217), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n614), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n631), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n625), .B2(new_n626), .ZN(new_n637));
  OAI211_X1 g451(.A(G469), .B(new_n636), .C1(new_n637), .C2(new_n615), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n601), .A2(new_n354), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n633), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(G221), .B1(new_n507), .B2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n600), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n467), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n309), .A2(new_n375), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT102), .B(G101), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G3));
  NAND2_X1  g462(.A1(new_n293), .A2(new_n354), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n649), .A2(G472), .B1(new_n293), .B2(new_n294), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n641), .A2(new_n642), .ZN(new_n651));
  AND4_X1   g465(.A1(new_n373), .A2(new_n651), .A3(new_n374), .A4(new_n599), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n441), .A2(new_n449), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT87), .B1(new_n436), .B2(new_n440), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n464), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n451), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n450), .A2(new_n452), .A3(new_n464), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n376), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n527), .A2(new_n514), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT103), .B1(new_n520), .B2(new_n526), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT33), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT33), .ZN(new_n664));
  OAI211_X1 g478(.A(KEYINPUT103), .B(new_n664), .C1(new_n520), .C2(new_n526), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n514), .A2(G902), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n588), .B1(new_n661), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n654), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT104), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT34), .B(G104), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  NAND2_X1  g488(.A1(new_n578), .A2(new_n585), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(KEYINPUT105), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n587), .A2(G475), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n677), .B1(new_n578), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n519), .A2(new_n530), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n660), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n654), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT35), .B(G107), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G9));
  NOR2_X1   g500(.A1(new_n351), .A2(KEYINPUT36), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n345), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n369), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n362), .B2(new_n367), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n645), .A2(new_n650), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  INV_X1    g507(.A(new_n376), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n657), .B2(new_n451), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n695), .A2(new_n659), .A3(new_n690), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n592), .B(KEYINPUT106), .Z(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n698), .B1(new_n699), .B2(new_n596), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n680), .A2(new_n681), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n643), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n298), .A2(new_n308), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT32), .B1(new_n293), .B2(new_n294), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n696), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XOR2_X1   g521(.A(new_n700), .B(KEYINPUT39), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n651), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT108), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT40), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n465), .A2(new_n466), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT38), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n690), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n588), .B1(new_n519), .B2(new_n530), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n717), .A2(new_n376), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n712), .A2(new_n713), .A3(new_n716), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n299), .A2(new_n278), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT107), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n286), .A2(new_n290), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n354), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G472), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n297), .A2(new_n725), .A3(new_n298), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n720), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n187), .ZN(G45));
  NAND3_X1  g543(.A1(new_n651), .A2(new_n668), .A3(new_n701), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n696), .B(new_n731), .C1(new_n704), .C2(new_n705), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  AOI21_X1  g547(.A(new_n620), .B1(new_n619), .B2(new_n621), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n623), .A2(KEYINPUT78), .A3(KEYINPUT12), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n626), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n632), .B1(new_n736), .B2(new_n635), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n737), .B2(G902), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n642), .A3(new_n633), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT109), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n738), .A2(new_n741), .A3(new_n642), .A4(new_n633), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n740), .A2(KEYINPUT110), .A3(new_n742), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n598), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n309), .A3(new_n375), .A4(new_n670), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT41), .B(G113), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G15));
  NAND4_X1  g564(.A1(new_n747), .A2(new_n309), .A3(new_n375), .A4(new_n683), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G116), .ZN(G18));
  NOR2_X1   g566(.A1(new_n743), .A2(new_n600), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n696), .B(new_n753), .C1(new_n704), .C2(new_n705), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  NAND4_X1  g569(.A1(new_n658), .A2(new_n376), .A3(new_n659), .A4(new_n718), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n695), .A2(KEYINPUT112), .A3(new_n659), .A4(new_n718), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n747), .ZN(new_n761));
  OAI22_X1  g575(.A1(new_n291), .A2(new_n292), .B1(new_n277), .B2(new_n300), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n649), .A2(G472), .B1(new_n294), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n764));
  INV_X1    g578(.A(new_n371), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT111), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n761), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n470), .ZN(G24));
  NOR2_X1   g584(.A1(new_n660), .A2(new_n743), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n668), .A2(new_n701), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n763), .A2(new_n771), .A3(new_n690), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  NOR3_X1   g589(.A1(new_n465), .A2(new_n466), .A3(new_n694), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n730), .A3(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n298), .B(new_n308), .C1(new_n705), .C2(KEYINPUT114), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n705), .A2(KEYINPUT114), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n779), .B(new_n765), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n465), .A2(new_n466), .A3(new_n643), .A4(new_n694), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n309), .A2(new_n375), .A3(new_n773), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n778), .B1(new_n784), .B2(new_n785), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  OAI211_X1 g604(.A(new_n783), .B(new_n375), .C1(new_n704), .C2(new_n705), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(new_n702), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND2_X1  g607(.A1(new_n667), .A2(new_n661), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n588), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT43), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n675), .A2(new_n677), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n796), .A2(new_n800), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n650), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n690), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n736), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n614), .B1(new_n810), .B2(new_n634), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(KEYINPUT45), .A3(new_n636), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT115), .Z(new_n813));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n811), .B2(new_n636), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n601), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n639), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n633), .B1(new_n816), .B2(KEYINPUT46), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT46), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n818), .B(new_n639), .C1(new_n813), .C2(new_n815), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n642), .A3(new_n708), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n809), .A2(new_n821), .A3(new_n777), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n201), .ZN(G39));
  INV_X1    g637(.A(new_n309), .ZN(new_n824));
  INV_X1    g638(.A(new_n375), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n773), .A4(new_n776), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(KEYINPUT47), .A3(new_n642), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n642), .B1(new_n817), .B2(new_n819), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT47), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n826), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(new_n312), .ZN(G42));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n765), .A2(new_n376), .A3(new_n642), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n835), .B2(new_n796), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n738), .B(new_n633), .C1(KEYINPUT118), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n834), .A2(KEYINPUT117), .A3(new_n795), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n836), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n716), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n727), .A3(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n774), .A2(new_n706), .A3(new_n732), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n643), .A2(new_n690), .A3(new_n700), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n760), .A2(new_n726), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n774), .A2(new_n706), .A3(new_n732), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n760), .A2(new_n726), .A3(new_n847), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT52), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n849), .A2(KEYINPUT120), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT120), .B1(new_n849), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n748), .A2(new_n751), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n517), .A2(new_n518), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n798), .A2(new_n858), .A3(KEYINPUT119), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n528), .A2(new_n529), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(new_n588), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n859), .A2(new_n668), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n467), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n650), .A2(new_n652), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n646), .A2(new_n691), .A3(new_n866), .A4(new_n754), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n769), .A2(new_n857), .A3(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n858), .A2(new_n680), .A3(new_n690), .A4(new_n701), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n309), .A2(new_n783), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n763), .A2(new_n690), .A3(new_n731), .A4(new_n776), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n870), .B(new_n871), .C1(new_n791), .C2(new_n702), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n868), .A2(new_n789), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n855), .A2(new_n856), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n849), .A2(new_n852), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(KEYINPUT53), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n874), .A2(new_n856), .A3(new_n876), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n856), .B1(new_n855), .B2(new_n874), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n738), .A2(new_n633), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n827), .B(new_n830), .C1(new_n642), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n697), .B1(new_n802), .B2(new_n804), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n766), .B2(new_n768), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(new_n776), .A3(new_n890), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n825), .A2(new_n777), .A3(new_n592), .A4(new_n743), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n794), .A2(new_n798), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n727), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n763), .A2(new_n690), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n743), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n888), .A2(new_n900), .A3(new_n776), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n896), .A2(new_n897), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n891), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n716), .A2(new_n376), .A3(new_n743), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n890), .A2(KEYINPUT50), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT121), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT50), .B1(new_n890), .B2(new_n904), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n906), .A2(new_n907), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n903), .A2(KEYINPUT51), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n890), .A2(new_n771), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n892), .A2(new_n727), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n591), .B1(new_n913), .B2(new_n669), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n901), .B(new_n765), .C1(new_n781), .C2(new_n780), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT48), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n917), .B(KEYINPUT48), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n891), .A2(new_n910), .A3(new_n902), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n908), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n911), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n885), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(G952), .A2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n844), .B1(new_n929), .B2(new_n930), .ZN(G75));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n846), .B1(new_n845), .B2(new_n848), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT52), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n849), .A2(new_n852), .A3(KEYINPUT120), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n768), .A2(new_n766), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n747), .A3(new_n760), .ZN(new_n939));
  INV_X1    g753(.A(new_n857), .ZN(new_n940));
  INV_X1    g754(.A(new_n867), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n873), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n782), .ZN(new_n943));
  INV_X1    g757(.A(new_n788), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n786), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT53), .B1(new_n937), .B2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(G210), .B(G902), .C1(new_n947), .C2(new_n880), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n462), .B(new_n463), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT55), .Z(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(KEYINPUT124), .B2(new_n949), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n948), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n948), .B2(new_n949), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n346), .A2(G952), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(G51));
  XNOR2_X1  g771(.A(new_n639), .B(KEYINPUT57), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n947), .A2(KEYINPUT54), .A3(new_n880), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n737), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n881), .A2(new_n882), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n964), .A2(G902), .A3(new_n813), .A4(new_n815), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n956), .B1(new_n963), .B2(new_n965), .ZN(G54));
  NAND2_X1  g780(.A1(KEYINPUT58), .A2(G475), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n964), .A2(G902), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n581), .A3(new_n582), .ZN(new_n970));
  INV_X1    g784(.A(new_n956), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n964), .A2(G902), .A3(new_n583), .A4(new_n968), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(G60));
  AND2_X1   g787(.A1(new_n663), .A2(new_n665), .ZN(new_n974));
  NAND2_X1  g788(.A1(G478), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT59), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n885), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n974), .A2(new_n976), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n959), .B2(new_n960), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n971), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n977), .A2(new_n980), .ZN(G63));
  XOR2_X1   g795(.A(KEYINPUT125), .B(KEYINPUT60), .Z(new_n982));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n947), .B2(new_n880), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n368), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n688), .B(new_n984), .C1(new_n947), .C2(new_n880), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n986), .A2(new_n971), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT61), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n986), .A2(KEYINPUT61), .A3(new_n971), .A4(new_n987), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(G66));
  INV_X1    g806(.A(new_n597), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n346), .B1(new_n993), .B2(G224), .ZN(new_n994));
  INV_X1    g808(.A(new_n868), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n346), .ZN(new_n996));
  INV_X1    g810(.A(G898), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n462), .B1(new_n997), .B2(G953), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n996), .B(new_n998), .ZN(G69));
  OAI21_X1  g813(.A(new_n845), .B1(new_n720), .B2(new_n727), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n822), .A2(new_n831), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n710), .A2(new_n776), .A3(new_n864), .ZN(new_n1004));
  OR3_X1    g818(.A1(new_n1004), .A2(new_n825), .A3(new_n824), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n282), .B1(new_n267), .B2(KEYINPUT30), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT126), .Z(new_n1008));
  OR2_X1    g822(.A1(new_n570), .A2(new_n573), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1006), .A2(new_n346), .A3(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n820), .A2(new_n642), .A3(new_n708), .A4(new_n760), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n765), .B1(new_n780), .B2(new_n781), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n792), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1015), .A2(new_n850), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1003), .A2(new_n1016), .A3(new_n346), .A4(new_n789), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G900), .A2(G953), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1011), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n346), .B1(G227), .B2(G900), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT127), .ZN(new_n1021));
  OR3_X1    g835(.A1(new_n1012), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1021), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1022), .A2(new_n1023), .ZN(G72));
  NOR2_X1   g838(.A1(new_n875), .A2(new_n878), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  NOR2_X1   g841(.A1(new_n304), .A2(new_n277), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(new_n723), .ZN(new_n1029));
  OR2_X1    g843(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1027), .B1(new_n1006), .B2(new_n995), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n304), .A2(new_n278), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1003), .A2(new_n1016), .A3(new_n789), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1027), .B1(new_n1034), .B2(new_n995), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(new_n278), .A3(new_n304), .ZN(new_n1036));
  AND4_X1   g850(.A1(new_n971), .A2(new_n1030), .A3(new_n1033), .A4(new_n1036), .ZN(G57));
endmodule


