

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  INV_X1 U322 ( .A(KEYINPUT112), .ZN(n420) );
  XNOR2_X1 U323 ( .A(n420), .B(KEYINPUT48), .ZN(n421) );
  XNOR2_X1 U324 ( .A(n422), .B(n421), .ZN(n524) );
  XOR2_X1 U325 ( .A(n562), .B(KEYINPUT36), .Z(n580) );
  NOR2_X1 U326 ( .A1(n526), .A2(n444), .ZN(n563) );
  XNOR2_X1 U327 ( .A(n408), .B(n407), .ZN(n562) );
  XNOR2_X1 U328 ( .A(KEYINPUT124), .B(G183GAT), .ZN(n445) );
  XNOR2_X1 U329 ( .A(n446), .B(n445), .ZN(G1350GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n291) );
  XNOR2_X1 U331 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n296) );
  XNOR2_X1 U333 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n292), .B(KEYINPUT70), .ZN(n380) );
  XOR2_X1 U335 ( .A(n380), .B(G155GAT), .Z(n294) );
  XOR2_X1 U336 ( .A(G15GAT), .B(G1GAT), .Z(n368) );
  XNOR2_X1 U337 ( .A(G22GAT), .B(n368), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n309) );
  XOR2_X1 U340 ( .A(G78GAT), .B(G211GAT), .Z(n298) );
  XNOR2_X1 U341 ( .A(G127GAT), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U343 ( .A(KEYINPUT80), .B(G64GAT), .Z(n300) );
  XNOR2_X1 U344 ( .A(G8GAT), .B(G71GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U346 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U347 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n304) );
  NAND2_X1 U348 ( .A1(G231GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U350 ( .A(KEYINPUT77), .B(n305), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U352 ( .A(n309), .B(n308), .Z(n575) );
  XOR2_X1 U353 ( .A(G120GAT), .B(G71GAT), .Z(n385) );
  XOR2_X1 U354 ( .A(G99GAT), .B(G15GAT), .Z(n311) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(G43GAT), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U357 ( .A(n385), .B(n312), .Z(n314) );
  NAND2_X1 U358 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U360 ( .A(G176GAT), .B(KEYINPUT20), .Z(n316) );
  XNOR2_X1 U361 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U363 ( .A(n318), .B(n317), .Z(n327) );
  XNOR2_X1 U364 ( .A(G127GAT), .B(KEYINPUT83), .ZN(n319) );
  XNOR2_X1 U365 ( .A(n319), .B(KEYINPUT0), .ZN(n320) );
  XOR2_X1 U366 ( .A(n320), .B(KEYINPUT82), .Z(n322) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(G134GAT), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n441) );
  XOR2_X1 U369 ( .A(KEYINPUT19), .B(G190GAT), .Z(n324) );
  XNOR2_X1 U370 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U372 ( .A(KEYINPUT18), .B(n325), .ZN(n356) );
  XOR2_X1 U373 ( .A(n441), .B(n356), .Z(n326) );
  XOR2_X1 U374 ( .A(n327), .B(n326), .Z(n517) );
  INV_X1 U375 ( .A(n517), .ZN(n526) );
  XOR2_X1 U376 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n329) );
  XNOR2_X1 U377 ( .A(KEYINPUT90), .B(KEYINPUT24), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n332) );
  XOR2_X1 U379 ( .A(G78GAT), .B(G148GAT), .Z(n331) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n381) );
  XOR2_X1 U382 ( .A(n332), .B(n381), .Z(n343) );
  XNOR2_X1 U383 ( .A(G211GAT), .B(KEYINPUT88), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n333), .B(KEYINPUT87), .ZN(n335) );
  INV_X1 U385 ( .A(KEYINPUT21), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n337) );
  XNOR2_X1 U387 ( .A(G197GAT), .B(G218GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n348) );
  XNOR2_X1 U389 ( .A(G50GAT), .B(G22GAT), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n338), .B(G141GAT), .ZN(n365) );
  XOR2_X1 U391 ( .A(n365), .B(KEYINPUT86), .Z(n340) );
  NAND2_X1 U392 ( .A1(G228GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n348), .B(n341), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U396 ( .A(KEYINPUT89), .B(G162GAT), .Z(n345) );
  XNOR2_X1 U397 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U399 ( .A(KEYINPUT3), .B(n346), .Z(n437) );
  XOR2_X1 U400 ( .A(n347), .B(n437), .Z(n462) );
  XOR2_X1 U401 ( .A(G176GAT), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U402 ( .A(n376), .B(n348), .ZN(n350) );
  AND2_X1 U403 ( .A1(G226GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n352) );
  INV_X1 U405 ( .A(G92GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n355) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(G36GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n353), .B(G8GAT), .ZN(n364) );
  XNOR2_X1 U409 ( .A(n364), .B(G204GAT), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n357) );
  XOR2_X1 U411 ( .A(n357), .B(n356), .Z(n492) );
  INV_X1 U412 ( .A(n492), .ZN(n515) );
  XOR2_X1 U413 ( .A(KEYINPUT7), .B(KEYINPUT67), .Z(n359) );
  XNOR2_X1 U414 ( .A(G43GAT), .B(G29GAT), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT8), .B(n360), .Z(n406) );
  XOR2_X1 U417 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n362) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U420 ( .A(n363), .B(KEYINPUT29), .Z(n367) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n369) );
  XOR2_X1 U423 ( .A(n369), .B(n368), .Z(n371) );
  XNOR2_X1 U424 ( .A(G197GAT), .B(G113GAT), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U426 ( .A(n406), .B(n372), .Z(n500) );
  INV_X1 U427 ( .A(n500), .ZN(n568) );
  XOR2_X1 U428 ( .A(G92GAT), .B(KEYINPUT72), .Z(n374) );
  XNOR2_X1 U429 ( .A(G99GAT), .B(G85GAT), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n401) );
  XNOR2_X1 U431 ( .A(n401), .B(KEYINPUT33), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n375), .B(KEYINPUT32), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n376), .B(KEYINPUT31), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n377), .B(KEYINPUT71), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n387) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n386) );
  XOR2_X1 U440 ( .A(n387), .B(n386), .Z(n572) );
  XOR2_X1 U441 ( .A(KEYINPUT41), .B(n572), .Z(n549) );
  NAND2_X1 U442 ( .A1(n568), .A2(n549), .ZN(n389) );
  INV_X1 U443 ( .A(KEYINPUT46), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n410) );
  XOR2_X1 U445 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n391) );
  XNOR2_X1 U446 ( .A(G36GAT), .B(KEYINPUT64), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U448 ( .A(KEYINPUT10), .B(G106GAT), .Z(n393) );
  XNOR2_X1 U449 ( .A(G134GAT), .B(G162GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U451 ( .A(n395), .B(n394), .Z(n400) );
  XOR2_X1 U452 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n397) );
  NAND2_X1 U453 ( .A1(G232GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U455 ( .A(KEYINPUT76), .B(n398), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n405) );
  XOR2_X1 U457 ( .A(KEYINPUT74), .B(n401), .Z(n403) );
  XNOR2_X1 U458 ( .A(G190GAT), .B(G218GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U460 ( .A(n405), .B(n404), .Z(n408) );
  XNOR2_X1 U461 ( .A(n406), .B(G50GAT), .ZN(n407) );
  OR2_X1 U462 ( .A1(n562), .A2(n575), .ZN(n409) );
  NOR2_X1 U463 ( .A1(n410), .A2(n409), .ZN(n412) );
  XNOR2_X1 U464 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n419) );
  XOR2_X1 U466 ( .A(n568), .B(KEYINPUT69), .Z(n555) );
  INV_X1 U467 ( .A(n575), .ZN(n482) );
  NOR2_X1 U468 ( .A1(n482), .A2(n580), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n413), .B(KEYINPUT45), .ZN(n414) );
  INV_X1 U470 ( .A(n572), .ZN(n447) );
  NAND2_X1 U471 ( .A1(n414), .A2(n447), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n415), .B(KEYINPUT110), .ZN(n416) );
  NOR2_X1 U473 ( .A1(n555), .A2(n416), .ZN(n417) );
  XOR2_X1 U474 ( .A(n417), .B(KEYINPUT111), .Z(n418) );
  NOR2_X1 U475 ( .A1(n419), .A2(n418), .ZN(n422) );
  NAND2_X1 U476 ( .A1(n515), .A2(n524), .ZN(n424) );
  XOR2_X1 U477 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n442) );
  XOR2_X1 U479 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n426) );
  XNOR2_X1 U480 ( .A(G1GAT), .B(G120GAT), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U482 ( .A(KEYINPUT91), .B(G57GAT), .Z(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U485 ( .A(n430), .B(n429), .Z(n439) );
  XOR2_X1 U486 ( .A(G85GAT), .B(G148GAT), .Z(n432) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(G141GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U489 ( .A(KEYINPUT92), .B(n433), .Z(n435) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U494 ( .A(n441), .B(n440), .Z(n513) );
  INV_X1 U495 ( .A(n513), .ZN(n488) );
  NAND2_X1 U496 ( .A1(n442), .A2(n488), .ZN(n566) );
  NOR2_X1 U497 ( .A1(n462), .A2(n566), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n443), .B(KEYINPUT55), .ZN(n444) );
  NAND2_X1 U499 ( .A1(n575), .A2(n563), .ZN(n446) );
  NAND2_X1 U500 ( .A1(n555), .A2(n447), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT73), .B(n448), .Z(n485) );
  NOR2_X1 U502 ( .A1(n562), .A2(n482), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n449), .B(KEYINPUT16), .ZN(n468) );
  XNOR2_X1 U504 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n450), .B(KEYINPUT25), .ZN(n454) );
  NAND2_X1 U506 ( .A1(n515), .A2(n517), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT94), .B(n451), .Z(n452) );
  NOR2_X1 U508 ( .A1(n462), .A2(n452), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(n458) );
  XOR2_X1 U510 ( .A(KEYINPUT93), .B(KEYINPUT26), .Z(n456) );
  NAND2_X1 U511 ( .A1(n462), .A2(n526), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(n567) );
  XNOR2_X1 U513 ( .A(n492), .B(KEYINPUT27), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n567), .A2(n461), .ZN(n457) );
  NOR2_X1 U515 ( .A1(n458), .A2(n457), .ZN(n459) );
  OR2_X1 U516 ( .A1(n513), .A2(n459), .ZN(n460) );
  XNOR2_X1 U517 ( .A(KEYINPUT97), .B(n460), .ZN(n466) );
  NOR2_X1 U518 ( .A1(n461), .A2(n488), .ZN(n525) );
  XOR2_X1 U519 ( .A(n462), .B(KEYINPUT66), .Z(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT28), .B(n463), .Z(n519) );
  INV_X1 U521 ( .A(n519), .ZN(n527) );
  NAND2_X1 U522 ( .A1(n525), .A2(n527), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n517), .A2(n464), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n480) );
  INV_X1 U525 ( .A(n480), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n501) );
  NOR2_X1 U527 ( .A1(n485), .A2(n501), .ZN(n476) );
  NAND2_X1 U528 ( .A1(n476), .A2(n513), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n470) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U533 ( .A1(n476), .A2(n515), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(G15GAT), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n517), .ZN(n474) );
  XNOR2_X1 U537 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NAND2_X1 U538 ( .A1(n476), .A2(n519), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n477), .B(KEYINPUT100), .ZN(n478) );
  XNOR2_X1 U540 ( .A(G22GAT), .B(n478), .ZN(G1327GAT) );
  INV_X1 U541 ( .A(KEYINPUT38), .ZN(n487) );
  XNOR2_X1 U542 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n479), .B(KEYINPUT101), .ZN(n484) );
  NOR2_X1 U544 ( .A1(n580), .A2(n480), .ZN(n481) );
  NAND2_X1 U545 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(n512) );
  NOR2_X1 U547 ( .A1(n512), .A2(n485), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n498) );
  NOR2_X1 U549 ( .A1(n498), .A2(n488), .ZN(n491) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT103), .B(n489), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  OR2_X1 U553 ( .A1(n498), .A2(n492), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n493), .ZN(n494) );
  XNOR2_X1 U555 ( .A(KEYINPUT104), .B(n494), .ZN(G1329GAT) );
  INV_X1 U556 ( .A(KEYINPUT40), .ZN(n496) );
  NOR2_X1 U557 ( .A1(n526), .A2(n498), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NOR2_X1 U560 ( .A1(n498), .A2(n527), .ZN(n499) );
  XOR2_X1 U561 ( .A(G50GAT), .B(n499), .Z(G1331GAT) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  XOR2_X1 U563 ( .A(KEYINPUT105), .B(n549), .Z(n557) );
  NAND2_X1 U564 ( .A1(n500), .A2(n557), .ZN(n511) );
  NOR2_X1 U565 ( .A1(n511), .A2(n501), .ZN(n507) );
  NAND2_X1 U566 ( .A1(n513), .A2(n507), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U568 ( .A1(n507), .A2(n515), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n517), .A2(n507), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U574 ( .A1(n507), .A2(n519), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n510), .Z(G1335GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n513), .A2(n520), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n520), .A2(n515), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n520), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n522) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n523), .Z(G1339GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n543) );
  NOR2_X1 U589 ( .A1(n526), .A2(n543), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U591 ( .A(KEYINPUT113), .B(n529), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n555), .A2(n540), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(KEYINPUT114), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U596 ( .A1(n540), .A2(n557), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U598 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n536) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n575), .A2(n540), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(KEYINPUT116), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n562), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n567), .A2(n543), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT119), .B(n544), .Z(n553) );
  NAND2_X1 U610 ( .A1(n553), .A2(n568), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n547) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(KEYINPUT52), .B(n548), .Z(n551) );
  NAND2_X1 U616 ( .A1(n553), .A2(n549), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n575), .A2(n553), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n553), .A2(n562), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n563), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n563), .A2(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT57), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n578), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT125), .Z(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  INV_X1 U643 ( .A(n578), .ZN(n579) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(G218GAT), .B(n583), .Z(G1355GAT) );
endmodule

