

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583;

  INV_X1 U325 ( .A(n418), .ZN(n378) );
  NOR2_X1 U326 ( .A1(n530), .A2(n521), .ZN(n430) );
  XNOR2_X1 U327 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U328 ( .A(n381), .B(n380), .ZN(n382) );
  NOR2_X1 U329 ( .A1(n538), .A2(n456), .ZN(n564) );
  XOR2_X1 U330 ( .A(KEYINPUT41), .B(n575), .Z(n552) );
  XNOR2_X1 U331 ( .A(n457), .B(G176GAT), .ZN(n458) );
  XNOR2_X1 U332 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT90), .B(G190GAT), .Z(n294) );
  XOR2_X1 U334 ( .A(G120GAT), .B(G71GAT), .Z(n377) );
  XOR2_X1 U335 ( .A(G134GAT), .B(KEYINPUT0), .Z(n437) );
  XNOR2_X1 U336 ( .A(n377), .B(n437), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U338 ( .A(n295), .B(G99GAT), .Z(n300) );
  XOR2_X1 U339 ( .A(KEYINPUT19), .B(KEYINPUT91), .Z(n297) );
  XNOR2_X1 U340 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U342 ( .A(G169GAT), .B(n298), .Z(n429) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(n429), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U345 ( .A(G15GAT), .B(G127GAT), .Z(n344) );
  XOR2_X1 U346 ( .A(n344), .B(G176GAT), .Z(n302) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U350 ( .A(G183GAT), .B(KEYINPUT20), .Z(n306) );
  XNOR2_X1 U351 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(n307), .ZN(n308) );
  XOR2_X1 U354 ( .A(n309), .B(n308), .Z(n466) );
  INV_X1 U355 ( .A(n466), .ZN(n538) );
  XOR2_X1 U356 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n311) );
  XNOR2_X1 U357 ( .A(KEYINPUT94), .B(KEYINPUT22), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(n312), .B(KEYINPUT98), .Z(n314) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G155GAT), .Z(n336) );
  XNOR2_X1 U361 ( .A(n336), .B(G106GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n320) );
  XOR2_X1 U363 ( .A(G162GAT), .B(KEYINPUT80), .Z(n316) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(G218GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n394) );
  XOR2_X1 U366 ( .A(KEYINPUT97), .B(n394), .Z(n318) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U369 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U370 ( .A(G78GAT), .B(G148GAT), .Z(n322) );
  XNOR2_X1 U371 ( .A(KEYINPUT76), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n373) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n323), .B(G211GAT), .ZN(n423) );
  XNOR2_X1 U375 ( .A(n373), .B(n423), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U377 ( .A(KEYINPUT96), .B(KEYINPUT2), .Z(n327) );
  XNOR2_X1 U378 ( .A(KEYINPUT3), .B(KEYINPUT95), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U380 ( .A(G141GAT), .B(n328), .Z(n451) );
  XOR2_X1 U381 ( .A(n329), .B(n451), .Z(n471) );
  XOR2_X1 U382 ( .A(KEYINPUT47), .B(KEYINPUT120), .Z(n408) );
  XOR2_X1 U383 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n335) );
  XNOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n330), .B(KEYINPUT74), .ZN(n376) );
  XOR2_X1 U386 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n332) );
  XNOR2_X1 U387 ( .A(G1GAT), .B(KEYINPUT14), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n376), .B(n333), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U391 ( .A(G8GAT), .B(G183GAT), .Z(n417) );
  XOR2_X1 U392 ( .A(n417), .B(n336), .Z(n338) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U395 ( .A(n340), .B(n339), .Z(n346) );
  XOR2_X1 U396 ( .A(G64GAT), .B(G211GAT), .Z(n342) );
  XNOR2_X1 U397 ( .A(G71GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U400 ( .A(n346), .B(n345), .Z(n460) );
  INV_X1 U401 ( .A(n460), .ZN(n578) );
  XOR2_X1 U402 ( .A(G15GAT), .B(G197GAT), .Z(n348) );
  XNOR2_X1 U403 ( .A(G141GAT), .B(G22GAT), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U405 ( .A(n349), .B(G36GAT), .Z(n351) );
  XOR2_X1 U406 ( .A(G113GAT), .B(G1GAT), .Z(n441) );
  XNOR2_X1 U407 ( .A(n441), .B(G50GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n357) );
  XOR2_X1 U409 ( .A(G29GAT), .B(G43GAT), .Z(n353) );
  XNOR2_X1 U410 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n401) );
  XOR2_X1 U412 ( .A(n401), .B(KEYINPUT29), .Z(n355) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(n357), .B(n356), .Z(n365) );
  XOR2_X1 U416 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n359) );
  XNOR2_X1 U417 ( .A(G169GAT), .B(G8GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U419 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n361) );
  XNOR2_X1 U420 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U423 ( .A(n365), .B(n364), .Z(n507) );
  INV_X1 U424 ( .A(n507), .ZN(n570) );
  XOR2_X1 U425 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n367) );
  XNOR2_X1 U426 ( .A(G92GAT), .B(KEYINPUT75), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n383) );
  XOR2_X1 U428 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n369) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U431 ( .A(n370), .B(KEYINPUT33), .Z(n375) );
  XOR2_X1 U432 ( .A(KEYINPUT77), .B(G85GAT), .Z(n372) );
  XNOR2_X1 U433 ( .A(G99GAT), .B(G106GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n400) );
  XNOR2_X1 U435 ( .A(n373), .B(n400), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n379) );
  XOR2_X1 U438 ( .A(G176GAT), .B(G64GAT), .Z(n418) );
  XOR2_X1 U439 ( .A(n383), .B(n382), .Z(n575) );
  NAND2_X1 U440 ( .A1(n570), .A2(n552), .ZN(n384) );
  XOR2_X1 U441 ( .A(KEYINPUT46), .B(n384), .Z(n385) );
  NOR2_X1 U442 ( .A1(n578), .A2(n385), .ZN(n406) );
  XOR2_X1 U443 ( .A(KEYINPUT83), .B(KEYINPUT9), .Z(n387) );
  XNOR2_X1 U444 ( .A(G134GAT), .B(KEYINPUT67), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n389) );
  XNOR2_X1 U447 ( .A(KEYINPUT11), .B(KEYINPUT81), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U449 ( .A(n391), .B(n390), .Z(n396) );
  XOR2_X1 U450 ( .A(KEYINPUT85), .B(G92GAT), .Z(n393) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(G190GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n421) );
  XNOR2_X1 U453 ( .A(n394), .B(n421), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n405) );
  XOR2_X1 U455 ( .A(KEYINPUT82), .B(KEYINPUT65), .Z(n398) );
  NAND2_X1 U456 ( .A1(G232GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U458 ( .A(n399), .B(KEYINPUT84), .Z(n403) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U461 ( .A(n405), .B(n404), .Z(n558) );
  INV_X1 U462 ( .A(n558), .ZN(n409) );
  NAND2_X1 U463 ( .A1(n406), .A2(n409), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n414) );
  XOR2_X1 U465 ( .A(KEYINPUT86), .B(n409), .Z(n565) );
  XNOR2_X1 U466 ( .A(KEYINPUT36), .B(n565), .ZN(n580) );
  NAND2_X1 U467 ( .A1(n580), .A2(n578), .ZN(n410) );
  XOR2_X1 U468 ( .A(KEYINPUT45), .B(n410), .Z(n412) );
  NOR2_X1 U469 ( .A1(n570), .A2(n575), .ZN(n411) );
  NAND2_X1 U470 ( .A1(n412), .A2(n411), .ZN(n413) );
  NAND2_X1 U471 ( .A1(n414), .A2(n413), .ZN(n416) );
  XOR2_X1 U472 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n530) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n427) );
  XOR2_X1 U475 ( .A(G218GAT), .B(KEYINPUT104), .Z(n420) );
  NAND2_X1 U476 ( .A1(G226GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U478 ( .A(n422), .B(n421), .Z(n425) );
  XNOR2_X1 U479 ( .A(G204GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n521) );
  XNOR2_X1 U483 ( .A(n430), .B(KEYINPUT54), .ZN(n454) );
  XOR2_X1 U484 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n432) );
  XNOR2_X1 U485 ( .A(KEYINPUT100), .B(KEYINPUT103), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U487 ( .A(KEYINPUT99), .B(KEYINPUT6), .Z(n434) );
  XNOR2_X1 U488 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(n436), .B(n435), .Z(n443) );
  XOR2_X1 U491 ( .A(n437), .B(KEYINPUT1), .Z(n439) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U496 ( .A(G85GAT), .B(G162GAT), .Z(n445) );
  XNOR2_X1 U497 ( .A(G29GAT), .B(G148GAT), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U499 ( .A(n447), .B(n446), .Z(n453) );
  XOR2_X1 U500 ( .A(G57GAT), .B(G155GAT), .Z(n449) );
  XNOR2_X1 U501 ( .A(G127GAT), .B(G120GAT), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n453), .B(n452), .ZN(n531) );
  NAND2_X1 U505 ( .A1(n454), .A2(n531), .ZN(n568) );
  NOR2_X1 U506 ( .A1(n471), .A2(n568), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n455), .B(KEYINPUT55), .ZN(n456) );
  NAND2_X1 U508 ( .A1(n564), .A2(n552), .ZN(n459) );
  XOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n457) );
  OR2_X1 U510 ( .A1(n507), .A2(n575), .ZN(n495) );
  NOR2_X1 U511 ( .A1(n565), .A2(n460), .ZN(n461) );
  XOR2_X1 U512 ( .A(KEYINPUT89), .B(n461), .Z(n462) );
  XNOR2_X1 U513 ( .A(KEYINPUT16), .B(n462), .ZN(n478) );
  XNOR2_X1 U514 ( .A(KEYINPUT27), .B(KEYINPUT105), .ZN(n463) );
  XOR2_X1 U515 ( .A(n463), .B(n521), .Z(n473) );
  INV_X1 U516 ( .A(n473), .ZN(n532) );
  XOR2_X1 U517 ( .A(n471), .B(KEYINPUT68), .Z(n464) );
  XNOR2_X1 U518 ( .A(KEYINPUT28), .B(n464), .ZN(n535) );
  NAND2_X1 U519 ( .A1(n532), .A2(n535), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U521 ( .A1(n531), .A2(n467), .ZN(n477) );
  NOR2_X1 U522 ( .A1(n538), .A2(n521), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n471), .A2(n468), .ZN(n469) );
  XNOR2_X1 U524 ( .A(KEYINPUT25), .B(n469), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n470), .A2(n531), .ZN(n475) );
  NAND2_X1 U526 ( .A1(n471), .A2(n538), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT26), .ZN(n569) );
  NOR2_X1 U528 ( .A1(n569), .A2(n473), .ZN(n474) );
  NOR2_X1 U529 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U530 ( .A1(n477), .A2(n476), .ZN(n491) );
  NAND2_X1 U531 ( .A1(n478), .A2(n491), .ZN(n479) );
  XNOR2_X1 U532 ( .A(n479), .B(KEYINPUT106), .ZN(n508) );
  NOR2_X1 U533 ( .A1(n495), .A2(n508), .ZN(n480) );
  XNOR2_X1 U534 ( .A(n480), .B(KEYINPUT107), .ZN(n487) );
  NOR2_X1 U535 ( .A1(n531), .A2(n487), .ZN(n481) );
  XOR2_X1 U536 ( .A(KEYINPUT34), .B(n481), .Z(n482) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U538 ( .A1(n521), .A2(n487), .ZN(n483) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  NOR2_X1 U540 ( .A1(n538), .A2(n487), .ZN(n485) );
  XNOR2_X1 U541 ( .A(KEYINPUT108), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n535), .A2(n487), .ZN(n489) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT109), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n490), .ZN(n494) );
  NAND2_X1 U549 ( .A1(n491), .A2(n580), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n578), .A2(n492), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n494), .B(n493), .ZN(n519) );
  NOR2_X1 U552 ( .A1(n519), .A2(n495), .ZN(n497) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT112), .Z(n496) );
  XNOR2_X1 U554 ( .A(n497), .B(n496), .ZN(n504) );
  NOR2_X1 U555 ( .A1(n531), .A2(n504), .ZN(n499) );
  XNOR2_X1 U556 ( .A(KEYINPUT113), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U558 ( .A(G29GAT), .B(n500), .Z(G1328GAT) );
  NOR2_X1 U559 ( .A1(n521), .A2(n504), .ZN(n501) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n501), .Z(G1329GAT) );
  NOR2_X1 U561 ( .A1(n538), .A2(n504), .ZN(n502) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(n502), .Z(n503) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NOR2_X1 U564 ( .A1(n535), .A2(n504), .ZN(n505) );
  XOR2_X1 U565 ( .A(KEYINPUT114), .B(n505), .Z(n506) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  NAND2_X1 U567 ( .A1(n552), .A2(n507), .ZN(n518) );
  NOR2_X1 U568 ( .A1(n518), .A2(n508), .ZN(n509) );
  XNOR2_X1 U569 ( .A(n509), .B(KEYINPUT115), .ZN(n515) );
  NOR2_X1 U570 ( .A1(n531), .A2(n515), .ZN(n510) );
  XOR2_X1 U571 ( .A(KEYINPUT42), .B(n510), .Z(n511) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n521), .A2(n515), .ZN(n512) );
  XOR2_X1 U574 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U575 ( .A1(n538), .A2(n515), .ZN(n513) );
  XOR2_X1 U576 ( .A(KEYINPUT116), .B(n513), .Z(n514) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U578 ( .A1(n535), .A2(n515), .ZN(n517) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  OR2_X1 U581 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U582 ( .A1(n531), .A2(n526), .ZN(n520) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n526), .ZN(n523) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT117), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n538), .A2(n526), .ZN(n524) );
  XOR2_X1 U588 ( .A(KEYINPUT118), .B(n524), .Z(n525) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  NOR2_X1 U590 ( .A1(n535), .A2(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT119), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT122), .ZN(n540) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U597 ( .A(KEYINPUT121), .B(n534), .Z(n549) );
  INV_X1 U598 ( .A(n549), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n570), .A2(n546), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n540), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U604 ( .A1(n546), .A2(n552), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT123), .Z(n544) );
  NAND2_X1 U607 ( .A1(n546), .A2(n578), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U611 ( .A1(n546), .A2(n565), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n569), .A2(n549), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n570), .A2(n559), .ZN(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT124), .B(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U618 ( .A1(n559), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT125), .Z(n557) );
  NAND2_X1 U622 ( .A1(n559), .A2(n578), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT126), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n570), .A2(n564), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n578), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .Z(n572) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n581), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

