//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(G110), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT70), .B(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n190));
  OR2_X1    g004(.A1(new_n190), .A2(KEYINPUT81), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(KEYINPUT81), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT82), .ZN(new_n194));
  OR2_X1    g008(.A1(new_n188), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n187), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n200), .A2(KEYINPUT16), .A3(G140), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(KEYINPUT16), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n203), .B(G146), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n189), .B1(new_n205), .B2(G128), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT24), .B(G110), .Z(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n199), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G953), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(G221), .A3(G234), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT22), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n213), .B(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n196), .A2(new_n187), .A3(new_n198), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n208), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n203), .A2(G146), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n202), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n210), .B(new_n214), .C1(new_n217), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G902), .ZN(new_n223));
  INV_X1    g037(.A(new_n214), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n221), .B1(new_n215), .B2(new_n216), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n199), .A2(new_n209), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n222), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT25), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT80), .B(G217), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(G234), .B2(new_n223), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n222), .A2(new_n227), .A3(new_n233), .A4(new_n223), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n222), .A2(new_n227), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n232), .A2(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT76), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n205), .A2(G116), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n188), .B2(G116), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n243));
  INV_X1    g057(.A(G113), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT2), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT2), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G113), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n242), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT70), .A2(G119), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT70), .A2(G119), .ZN(new_n251));
  OAI21_X1  g065(.A(G116), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n241), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n248), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT72), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n260));
  AOI211_X1 g074(.A(new_n260), .B(new_n257), .C1(new_n249), .C2(new_n255), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G143), .B(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  OR2_X1    g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n263), .A2(new_n264), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT64), .B(G134), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G134), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(KEYINPUT64), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT67), .B(G137), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(KEYINPUT11), .A2(G134), .ZN(new_n280));
  AND2_X1   g094(.A1(KEYINPUT65), .A2(G137), .ZN(new_n281));
  NOR2_X1   g095(.A1(KEYINPUT65), .A2(G137), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT65), .B(G137), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT66), .A3(new_n280), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G131), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n276), .A2(KEYINPUT64), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n274), .A2(G134), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(new_n272), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT11), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n279), .A2(new_n288), .A3(new_n289), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n273), .A2(new_n278), .B1(new_n293), .B2(new_n292), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n289), .B1(new_n297), .B2(new_n288), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n269), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n286), .B2(G134), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n292), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n286), .A2(new_n300), .A3(G134), .ZN(new_n303));
  OAI21_X1  g117(.A(G131), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n305));
  INV_X1    g119(.A(G143), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(G146), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n197), .A2(new_n219), .A3(G143), .ZN(new_n308));
  INV_X1    g122(.A(new_n263), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(new_n305), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n295), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n262), .A2(new_n299), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(KEYINPUT28), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n243), .B1(new_n242), .B2(new_n248), .ZN(new_n315));
  AND4_X1   g129(.A1(new_n243), .A2(new_n252), .A3(new_n248), .A4(new_n253), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n258), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n260), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n256), .A2(KEYINPUT72), .A3(new_n258), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n271), .A2(new_n270), .A3(new_n272), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n290), .A2(new_n291), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT67), .B1(new_n323), .B2(G137), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n294), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n288), .ZN(new_n326));
  OAI21_X1  g140(.A(G131), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n268), .B1(new_n327), .B2(new_n295), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n295), .A2(new_n304), .A3(new_n310), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n320), .B(new_n321), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n299), .A2(new_n311), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n321), .B1(new_n332), .B2(new_n320), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n312), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n314), .B1(new_n334), .B2(KEYINPUT28), .ZN(new_n335));
  INV_X1    g149(.A(G237), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n211), .A3(G210), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n337), .B(KEYINPUT74), .Z(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT26), .B(G101), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n240), .B1(new_n335), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(KEYINPUT69), .A2(KEYINPUT30), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n344), .B(new_n347), .C1(new_n328), .C2(new_n329), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n299), .A2(new_n345), .A3(new_n346), .A4(new_n311), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n320), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n312), .A3(new_n342), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT31), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n313), .B1(new_n350), .B2(new_n320), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT31), .A3(new_n342), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n314), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n320), .B1(new_n328), .B2(new_n329), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT75), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n313), .B1(new_n360), .B2(new_n330), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n342), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT76), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n343), .A2(new_n357), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT32), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT32), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n370), .A3(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n373));
  OR3_X1    g187(.A1(new_n355), .A2(new_n373), .A3(new_n342), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n358), .B(new_n342), .C1(new_n361), .C2(new_n362), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n355), .B2(new_n342), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n223), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n312), .A2(new_n359), .A3(KEYINPUT78), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n332), .A2(new_n381), .A3(new_n320), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(KEYINPUT28), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n358), .A2(new_n383), .A3(new_n384), .ZN(new_n386));
  AOI211_X1 g200(.A(new_n377), .B(new_n364), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G472), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n239), .B1(new_n372), .B2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(G110), .B(G122), .Z(new_n390));
  INV_X1    g204(.A(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(new_n391), .B2(G107), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n393));
  INV_X1    g207(.A(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(G107), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n395), .A3(new_n399), .A4(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n401), .B(new_n402), .C1(KEYINPUT4), .C2(new_n398), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n398), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n400), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n318), .A2(new_n319), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(G113), .C1(KEYINPUT5), .C2(new_n252), .ZN(new_n407));
  INV_X1    g221(.A(new_n396), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n391), .A2(G107), .ZN(new_n409));
  OAI21_X1  g223(.A(G101), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n410), .A2(new_n400), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n407), .A2(new_n256), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n390), .B1(new_n405), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n412), .ZN(new_n414));
  INV_X1    g228(.A(new_n390), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n402), .B1(new_n398), .B2(KEYINPUT4), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n404), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n414), .B(new_n415), .C1(new_n262), .C2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(new_n420), .A3(KEYINPUT6), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n269), .A2(G125), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n310), .A2(new_n200), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n422), .B2(new_n424), .ZN(new_n426));
  INV_X1    g240(.A(G224), .ZN(new_n427));
  OAI22_X1  g241(.A1(new_n425), .A2(new_n426), .B1(new_n427), .B2(G953), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT86), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n427), .A2(G953), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(new_n390), .C1(new_n405), .C2(new_n412), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n421), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT7), .B1(new_n427), .B2(G953), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n429), .B(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n390), .B(KEYINPUT8), .Z(new_n440));
  AOI21_X1  g254(.A(new_n411), .B1(new_n407), .B2(new_n256), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n412), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n420), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n223), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n437), .A2(new_n223), .A3(new_n445), .A4(new_n443), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G214), .B1(G237), .B2(G902), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G221), .ZN(new_n453));
  XOR2_X1   g267(.A(KEYINPUT9), .B(G234), .Z(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n454), .B2(new_n223), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n211), .A2(G227), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT10), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n418), .A2(new_n269), .B1(KEYINPUT84), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n296), .A2(new_n298), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n411), .A2(new_n310), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n461), .A2(KEYINPUT84), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n462), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n460), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT85), .B(new_n460), .C1(new_n467), .C2(new_n468), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n473));
  INV_X1    g287(.A(new_n463), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n411), .B(new_n310), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n474), .A2(KEYINPUT12), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT12), .B1(new_n474), .B2(new_n475), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n473), .B(new_n459), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G469), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n223), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n223), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n467), .A2(new_n468), .A3(new_n460), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n460), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n485), .B2(G469), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n204), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G214), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n490), .A2(G237), .A3(G953), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n306), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT87), .B(G143), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(new_n289), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n289), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(KEYINPUT17), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n204), .A2(new_n488), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n489), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n391), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n496), .A2(KEYINPUT18), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n495), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n202), .B(new_n219), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .A4(new_n499), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n503), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n512));
  NOR2_X1   g326(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n202), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n202), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n515));
  AOI21_X1  g329(.A(G146), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n218), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n518), .A2(KEYINPUT89), .B1(new_n497), .B2(new_n499), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n506), .A2(new_n509), .A3(new_n499), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n508), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n511), .B1(new_n522), .B2(new_n505), .ZN(new_n523));
  INV_X1    g337(.A(G475), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n223), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT20), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n524), .A4(new_n223), .ZN(new_n528));
  INV_X1    g342(.A(new_n511), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n505), .B1(new_n503), .B2(new_n510), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n223), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G475), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n454), .A2(new_n211), .A3(new_n230), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT13), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n306), .A2(KEYINPUT91), .A3(G128), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT91), .B1(new_n306), .B2(G128), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n306), .A2(G128), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n197), .B2(G143), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n306), .A2(KEYINPUT91), .A3(G128), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT13), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n545), .A2(new_n546), .A3(G134), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n546), .B1(new_n545), .B2(G134), .ZN(new_n548));
  XNOR2_X1  g362(.A(G116), .B(G122), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(new_n394), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n542), .A2(new_n543), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n323), .A3(new_n540), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n547), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n540), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n271), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n556), .A2(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n394), .ZN(new_n558));
  INV_X1    g372(.A(new_n549), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT14), .ZN(new_n560));
  INV_X1    g374(.A(G116), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT14), .A3(G122), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G107), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n558), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n534), .B1(new_n554), .B2(new_n565), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n557), .A2(new_n564), .ZN(new_n567));
  INV_X1    g381(.A(new_n534), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n545), .A2(G134), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT92), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n545), .A2(new_n546), .A3(G134), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n567), .B(new_n568), .C1(new_n572), .C2(new_n553), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n573), .A3(KEYINPUT93), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n575), .B(new_n534), .C1(new_n554), .C2(new_n565), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n223), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G478), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT15), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n577), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(G234), .A2(G237), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n581), .A2(G952), .A3(new_n211), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT21), .B(G898), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT94), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n581), .A2(G902), .A3(G953), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n533), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n452), .A2(new_n456), .A3(new_n487), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n389), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND2_X1  g406(.A1(new_n366), .A2(new_n223), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n594), .A2(KEYINPUT95), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n594), .A2(KEYINPUT95), .B1(new_n367), .B2(new_n366), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n239), .A2(new_n455), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n598), .A2(new_n487), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT96), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n574), .A2(new_n603), .A3(new_n576), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n566), .A2(new_n573), .A3(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n223), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G478), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n577), .A2(G478), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n608), .B1(new_n607), .B2(new_n609), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n447), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n437), .A2(new_n223), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n445), .A4(new_n443), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n448), .A2(KEYINPUT97), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n444), .A2(KEYINPUT98), .A3(new_n446), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n615), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n587), .ZN(new_n622));
  AND4_X1   g436(.A1(new_n450), .A2(new_n613), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n602), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n624), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n611), .A2(new_n580), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n450), .A2(new_n621), .A3(new_n622), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n602), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n225), .A2(new_n226), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n636), .B(new_n637), .Z(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n237), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n235), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n595), .A2(new_n596), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT103), .A4(new_n640), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n590), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT37), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n187), .ZN(G12));
  AND3_X1   g461(.A1(new_n366), .A2(new_n370), .A3(new_n367), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n370), .B1(new_n366), .B2(new_n367), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n388), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n621), .A2(new_n450), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n487), .A2(new_n456), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n582), .B1(new_n586), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n628), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n650), .A2(new_n653), .A3(new_n640), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  OR2_X1    g472(.A1(new_n355), .A2(new_n364), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n342), .B1(new_n380), .B2(new_n382), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(G902), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n648), .B2(new_n649), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI211_X1 g480(.A(KEYINPUT104), .B(new_n663), .C1(new_n648), .C2(new_n649), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n655), .B(KEYINPUT39), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT40), .B1(new_n652), .B2(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n533), .A2(new_n450), .A3(new_n580), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n449), .B(KEYINPUT38), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n652), .A2(KEYINPUT40), .A3(new_n669), .ZN(new_n675));
  OR3_X1    g489(.A1(new_n674), .A2(new_n640), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  INV_X1    g491(.A(new_n613), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n655), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n650), .A2(new_n653), .A3(new_n679), .A4(new_n640), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  INV_X1    g495(.A(new_n239), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n479), .A2(new_n480), .A3(new_n223), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n480), .B1(new_n479), .B2(new_n223), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n683), .A2(new_n684), .A3(new_n455), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n650), .A2(new_n623), .A3(new_n682), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT41), .B(G113), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  AND4_X1   g502(.A1(new_n650), .A2(new_n630), .A3(new_n682), .A4(new_n685), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n561), .ZN(G18));
  AND4_X1   g504(.A1(new_n450), .A2(new_n621), .A3(new_n685), .A4(new_n588), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n650), .A2(new_n691), .A3(new_n640), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n650), .A2(new_n691), .A3(KEYINPUT105), .A4(new_n640), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(new_n367), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n385), .A2(new_n364), .A3(new_n386), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n698), .B1(new_n699), .B2(new_n357), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n594), .A2(new_n682), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT106), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n700), .B1(new_n593), .B2(G472), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n682), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n587), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n685), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n621), .A2(new_n671), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n621), .A2(KEYINPUT107), .A3(new_n671), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NOR2_X1   g529(.A1(new_n651), .A2(new_n708), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT108), .B1(new_n704), .B2(new_n640), .ZN(new_n717));
  INV_X1    g531(.A(G472), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n366), .B2(new_n223), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n235), .A2(new_n639), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n719), .A2(new_n720), .A3(new_n700), .A4(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n679), .B(new_n716), .C1(new_n717), .C2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  NAND3_X1  g538(.A1(new_n447), .A2(new_n450), .A3(new_n448), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n652), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n389), .A2(KEYINPUT42), .A3(new_n679), .A4(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n650), .A2(new_n679), .A3(new_n682), .A4(new_n726), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NAND2_X1  g546(.A1(new_n650), .A2(new_n682), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n733), .A2(new_n652), .A3(new_n725), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n656), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  XOR2_X1   g550(.A(new_n485), .B(KEYINPUT45), .Z(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  INV_X1    g552(.A(new_n482), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(G469), .C1(new_n737), .C2(G902), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n481), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n456), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n669), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n725), .B(KEYINPUT110), .Z(new_n746));
  NOR2_X1   g560(.A1(new_n610), .A2(new_n612), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n611), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT109), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT43), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n640), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n597), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n746), .B1(new_n752), .B2(KEYINPUT44), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n755), .B(new_n757), .C1(new_n751), .C2(new_n597), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n745), .B(new_n753), .C1(new_n756), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n744), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n743), .A2(KEYINPUT47), .A3(new_n456), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n679), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(new_n682), .A3(new_n725), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n372), .A3(new_n388), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  NOR2_X1   g583(.A1(new_n708), .A2(new_n725), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT119), .Z(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n582), .A3(new_n750), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n733), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT48), .Z(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(G952), .A3(new_n211), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n750), .A2(new_n582), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n706), .B2(new_n703), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n708), .A2(new_n450), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n673), .B1(new_n778), .B2(KEYINPUT118), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n777), .B(new_n779), .C1(KEYINPUT118), .C2(new_n778), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT50), .Z(new_n781));
  INV_X1    g595(.A(new_n668), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n771), .A2(new_n782), .A3(new_n682), .A4(new_n582), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n533), .A3(new_n747), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n594), .A2(new_n640), .A3(new_n701), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n721), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n704), .A2(KEYINPUT108), .A3(new_n640), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n772), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n746), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n777), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n683), .A2(new_n684), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n455), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n763), .A2(new_n764), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT120), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(KEYINPUT120), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n781), .A2(new_n789), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT51), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n794), .B1(new_n765), .B2(KEYINPUT117), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n765), .A2(KEYINPUT117), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n792), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n781), .A2(new_n803), .A3(new_n789), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n775), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n777), .A2(new_n716), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n629), .A2(KEYINPUT113), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n629), .A2(KEYINPUT113), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n678), .A3(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n811), .A2(new_n452), .A3(new_n622), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n597), .A3(new_n599), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n645), .A2(new_n591), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n389), .A2(new_n630), .A3(new_n685), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n720), .B1(new_n372), .B2(new_n388), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT105), .B1(new_n816), .B2(new_n691), .ZN(new_n817));
  INV_X1    g631(.A(new_n695), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n389), .A2(new_n623), .A3(new_n685), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n705), .B1(new_n704), .B2(new_n682), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n719), .A2(KEYINPUT106), .A3(new_n700), .A4(new_n239), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n622), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n713), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT112), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n686), .B1(new_n707), .B2(new_n713), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n689), .B1(new_n694), .B2(new_n695), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n814), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n766), .B1(new_n786), .B2(new_n787), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n533), .A2(new_n580), .ZN(new_n833));
  INV_X1    g647(.A(new_n655), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n650), .A2(new_n833), .A3(new_n640), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n726), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n731), .A3(new_n735), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n711), .A2(new_n712), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n652), .A2(new_n640), .A3(new_n655), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n668), .A2(new_n839), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n723), .A2(new_n657), .A3(new_n680), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n668), .A2(new_n839), .A3(new_n842), .A4(new_n843), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n657), .A2(new_n680), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT52), .A4(new_n723), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n837), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n831), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT53), .B1(new_n831), .B2(new_n850), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT54), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n846), .A2(new_n849), .ZN(new_n856));
  INV_X1    g670(.A(new_n837), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n814), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n819), .A2(new_n825), .A3(KEYINPUT112), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n829), .B1(new_n827), .B2(new_n828), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n852), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n827), .A2(new_n828), .A3(KEYINPUT116), .A4(new_n731), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT53), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n827), .A2(new_n828), .A3(new_n731), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n836), .A2(new_n735), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n870), .A2(new_n856), .A3(new_n872), .A4(new_n859), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n854), .A2(KEYINPUT115), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n865), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI221_X1 g689(.A(new_n855), .B1(new_n678), .B2(new_n783), .C1(new_n875), .C2(KEYINPUT54), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n808), .A2(new_n876), .B1(G952), .B2(G953), .ZN(new_n877));
  INV_X1    g691(.A(new_n793), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n878), .A2(KEYINPUT49), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(KEYINPUT49), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n879), .A2(new_n880), .A3(new_n673), .A4(new_n748), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n450), .A3(new_n598), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n877), .B1(new_n668), .B2(new_n882), .ZN(G75));
  NAND2_X1  g697(.A1(new_n421), .A2(new_n436), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(new_n434), .Z(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n875), .A2(G210), .A3(G902), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n211), .A2(G952), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT123), .Z(new_n892));
  OR2_X1    g706(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n886), .B1(KEYINPUT121), .B2(KEYINPUT56), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n888), .A2(new_n897), .A3(new_n893), .A4(new_n894), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n890), .B(new_n892), .C1(new_n896), .C2(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n739), .A2(KEYINPUT57), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT115), .B1(new_n851), .B2(new_n852), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n864), .B(KEYINPUT53), .C1(new_n831), .C2(new_n850), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n901), .B1(new_n904), .B2(new_n873), .ZN(new_n905));
  AND4_X1   g719(.A1(new_n901), .A2(new_n865), .A3(new_n874), .A4(new_n873), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n739), .A2(KEYINPUT57), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n479), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n223), .B1(new_n904), .B2(new_n873), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(G469), .A3(new_n737), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n891), .B1(new_n909), .B2(new_n911), .ZN(G54));
  NAND3_X1  g726(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  INV_X1    g727(.A(new_n523), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n891), .ZN(G60));
  NAND2_X1  g731(.A1(new_n604), .A2(new_n605), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT59), .Z(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n905), .B2(new_n906), .ZN(new_n922));
  INV_X1    g736(.A(new_n892), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n855), .B1(new_n875), .B2(KEYINPUT54), .ZN(new_n925));
  INV_X1    g739(.A(new_n920), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n925), .A2(new_n926), .B1(new_n604), .B2(new_n605), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT124), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n926), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n918), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n930), .A2(new_n931), .A3(new_n923), .A4(new_n922), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT60), .Z(new_n935));
  XNOR2_X1  g749(.A(new_n638), .B(KEYINPUT125), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n875), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n875), .A2(new_n935), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n923), .B(new_n937), .C1(new_n938), .C2(new_n236), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G66));
  OAI21_X1  g755(.A(G953), .B1(new_n585), .B2(new_n427), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n831), .B2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n884), .B1(G898), .B2(new_n211), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT126), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G69));
  NAND3_X1  g760(.A1(new_n745), .A2(new_n389), .A3(new_n839), .ZN(new_n947));
  INV_X1    g761(.A(new_n845), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n948), .A2(new_n731), .A3(new_n735), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n760), .A2(new_n768), .A3(new_n947), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n211), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(G900), .B2(new_n211), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n514), .A2(new_n515), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n350), .B(new_n954), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n951), .B(new_n957), .C1(G900), .C2(new_n211), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n760), .A2(new_n768), .ZN(new_n960));
  INV_X1    g774(.A(new_n669), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n734), .A2(new_n961), .A3(new_n811), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT62), .B1(new_n676), .B2(new_n948), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n676), .A2(KEYINPUT62), .A3(new_n948), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n960), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n955), .B1(new_n966), .B2(G953), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n211), .B1(G227), .B2(G900), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n959), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n959), .B2(new_n967), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G72));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n965), .B2(new_n862), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n891), .B1(new_n974), .B2(new_n660), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n950), .B2(new_n862), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n355), .A3(new_n364), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n374), .A2(new_n352), .A3(new_n376), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n973), .B(new_n978), .C1(new_n853), .C2(new_n854), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n975), .A2(new_n977), .A3(new_n979), .ZN(G57));
endmodule


