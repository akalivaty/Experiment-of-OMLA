//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  AND2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G244), .ZN(new_n213));
  AND2_X1   g0013(.A1(new_n213), .A2(G77), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n209), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G20), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n212), .B1(new_n220), .B2(KEYINPUT1), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G50), .B(G68), .Z(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  INV_X1    g0041(.A(G1), .ZN(new_n242));
  OAI21_X1  g0042(.A(new_n242), .B1(G41), .B2(G45), .ZN(new_n243));
  INV_X1    g0043(.A(G274), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n243), .A2(KEYINPUT66), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n222), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT66), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n250), .B(new_n242), .C1(G41), .C2(G45), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n246), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n261), .A2(G223), .B1(new_n264), .B2(G77), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G222), .A3(new_n256), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n221), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n255), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n273), .A2(G179), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(new_n209), .B2(new_n258), .ZN(new_n276));
  NAND4_X1  g0076(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n221), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G20), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n203), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT8), .B(G58), .Z(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n278), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G20), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n278), .B1(new_n242), .B2(G20), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G50), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n273), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n274), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n288), .A2(KEYINPUT9), .A3(new_n294), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n273), .A2(G200), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n255), .A2(new_n271), .A3(G190), .A4(new_n272), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n306), .A3(new_n302), .ZN(new_n308));
  INV_X1    g0108(.A(new_n305), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n299), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n283), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(G20), .B2(G77), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n281), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n291), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n319), .A2(new_n278), .B1(new_n204), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n293), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n204), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n261), .A2(G238), .B1(new_n264), .B2(G107), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n266), .A2(G232), .A3(new_n256), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n270), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n245), .B1(new_n328), .B2(new_n213), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI211_X1 g0132(.A(new_n323), .B(new_n332), .C1(G200), .C2(new_n330), .ZN(new_n333));
  INV_X1    g0133(.A(new_n330), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n323), .B1(G169), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT70), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(new_n334), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n335), .A2(new_n336), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n311), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT75), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT18), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n282), .A2(new_n291), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n293), .B2(new_n282), .ZN(new_n345));
  AND2_X1   g0145(.A1(G58), .A2(G68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G58), .A2(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n285), .A2(G159), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n259), .A2(new_n279), .A3(new_n260), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT7), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n259), .A2(new_n356), .A3(new_n279), .A4(new_n260), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(G68), .A3(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n348), .A2(new_n350), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n278), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n353), .B1(new_n359), .B2(new_n358), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n345), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n247), .A2(new_n249), .A3(G232), .A4(new_n251), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G223), .A2(G1698), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n253), .B2(G1698), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n266), .B1(G33), .B2(G87), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n364), .B(new_n246), .C1(new_n367), .C2(new_n249), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G169), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n253), .A2(G1698), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(G223), .B2(G1698), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n372), .B2(new_n264), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n245), .B1(new_n373), .B2(new_n270), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(G179), .A3(new_n364), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n343), .B1(new_n363), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n363), .A2(new_n343), .A3(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT17), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n368), .A2(G190), .ZN(new_n382));
  AOI21_X1  g0182(.A(G200), .B1(new_n374), .B2(new_n364), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n363), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n358), .A2(new_n359), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n352), .A3(new_n351), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n278), .A3(new_n360), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n368), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G190), .B2(new_n368), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT17), .A4(new_n345), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT74), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n385), .A2(KEYINPUT74), .A3(new_n392), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n380), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G68), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n290), .A2(G20), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g0201(.A(new_n401), .B(KEYINPUT12), .Z(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n322), .B2(new_n398), .ZN(new_n403));
  INV_X1    g0203(.A(G50), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n286), .A2(new_n404), .B1(new_n279), .B2(G68), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n283), .A2(new_n204), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n278), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g0207(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n408));
  XNOR2_X1  g0208(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n266), .A2(G232), .A3(G1698), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n266), .A2(G226), .A3(new_n256), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n270), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n245), .B1(new_n328), .B2(G238), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n418), .B1(new_n416), .B2(new_n417), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT14), .B1(new_n421), .B2(new_n296), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(G179), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n421), .A2(KEYINPUT14), .A3(new_n296), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n411), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n421), .A2(G190), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n410), .C1(new_n389), .C2(new_n421), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n341), .A2(new_n342), .A3(new_n397), .A4(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n311), .A2(new_n426), .A3(new_n340), .A4(new_n428), .ZN(new_n431));
  INV_X1    g0231(.A(new_n379), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n377), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n385), .A2(KEYINPUT74), .A3(new_n392), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT74), .B1(new_n385), .B2(new_n392), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT75), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n242), .A2(G45), .ZN(new_n439));
  OR2_X1    g0239(.A1(KEYINPUT5), .A2(G41), .ZN(new_n440));
  NAND2_X1  g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(G274), .A4(new_n249), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  INV_X1    g0246(.A(new_n441), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(G274), .B1(new_n269), .B2(new_n221), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT76), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n442), .A2(new_n270), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G264), .ZN(new_n454));
  OAI211_X1 g0254(.A(G250), .B(new_n256), .C1(new_n262), .C2(new_n263), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G294), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n261), .A2(KEYINPUT85), .A3(G257), .ZN(new_n458));
  OAI211_X1 g0258(.A(G257), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n452), .B(new_n454), .C1(new_n462), .C2(new_n249), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n296), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n455), .A2(new_n456), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT85), .B1(new_n261), .B2(G257), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n459), .A2(new_n460), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n468), .A2(new_n270), .B1(G264), .B2(new_n453), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(new_n337), .A3(new_n452), .ZN(new_n470));
  INV_X1    g0270(.A(new_n278), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT23), .B1(new_n279), .B2(G107), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT23), .ZN(new_n473));
  INV_X1    g0273(.A(G107), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(G20), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n279), .A2(G33), .A3(G116), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT83), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n477), .B(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n279), .B(G87), .C1(new_n262), .C2(new_n263), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n480), .B(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT24), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n477), .B(KEYINPUT83), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(new_n481), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n480), .A2(new_n481), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n471), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n291), .A2(G107), .ZN(new_n490));
  XOR2_X1   g0290(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n491));
  XNOR2_X1  g0291(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n290), .A2(G20), .B1(new_n242), .B2(G33), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n471), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n494), .B2(new_n474), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n464), .B(new_n470), .C1(new_n489), .C2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(G244), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n497));
  OAI211_X1 g0297(.A(G238), .B(new_n256), .C1(new_n262), .C2(new_n263), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G116), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n270), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT78), .B1(new_n445), .B2(G1), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT78), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n242), .A3(G45), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G250), .B1(new_n269), .B2(new_n221), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n505), .A2(new_n506), .B1(new_n244), .B2(new_n439), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT79), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n501), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n337), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n266), .A2(new_n279), .A3(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n279), .B1(new_n414), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G87), .B2(new_n207), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n283), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n278), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n320), .A2(new_n312), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n494), .C2(new_n312), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n501), .A2(new_n508), .A3(new_n511), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n511), .B1(new_n501), .B2(new_n508), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n513), .B(new_n523), .C1(new_n526), .C2(G169), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n510), .A2(G190), .A3(new_n512), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n471), .A2(G87), .A3(new_n493), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n521), .A2(new_n530), .A3(new_n522), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n496), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(G244), .B(new_n256), .C1(new_n262), .C2(new_n263), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n256), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n270), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n444), .A2(new_n451), .B1(new_n453), .B2(G257), .ZN(new_n542));
  AOI21_X1  g0342(.A(G169), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n277), .A2(new_n221), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n493), .A2(new_n544), .A3(G97), .A4(new_n276), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n320), .A2(new_n518), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n286), .A2(new_n204), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  AND2_X1   g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n206), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n474), .A2(KEYINPUT6), .A3(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n548), .B1(new_n553), .B2(G20), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n355), .A2(G107), .A3(new_n357), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n547), .B1(new_n556), .B2(new_n278), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n543), .A2(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n541), .A2(new_n337), .A3(new_n542), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n389), .B1(new_n541), .B2(new_n542), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT77), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n541), .A2(new_n542), .A3(G190), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n557), .B(new_n566), .C1(new_n562), .C2(new_n563), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n561), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n533), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT86), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n469), .A2(new_n570), .A3(new_n331), .A4(new_n452), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT86), .B1(new_n463), .B2(G190), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n463), .A2(new_n389), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n489), .A2(new_n495), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n290), .A2(G20), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n493), .A2(new_n544), .A3(G116), .A4(new_n276), .ZN(new_n579));
  AOI21_X1  g0379(.A(G20), .B1(G33), .B2(G283), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n258), .A2(G97), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n580), .A2(new_n581), .B1(G20), .B2(new_n577), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n278), .A2(KEYINPUT20), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT20), .B1(new_n278), .B2(new_n582), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n578), .B(new_n579), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G264), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(new_n256), .C1(new_n262), .C2(new_n263), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n259), .A2(G303), .A3(new_n260), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n270), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n453), .A2(G270), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n452), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n585), .A2(new_n592), .A3(G169), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT80), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n585), .A2(new_n592), .A3(KEYINPUT80), .A4(G169), .ZN(new_n596));
  XOR2_X1   g0396(.A(KEYINPUT81), .B(KEYINPUT21), .Z(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n592), .A2(KEYINPUT21), .A3(G169), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n592), .A2(new_n337), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n585), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n585), .B1(G200), .B2(new_n592), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n331), .B2(new_n592), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n598), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n576), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n438), .A2(new_n569), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT87), .ZN(G372));
  AND2_X1   g0407(.A1(new_n339), .A2(new_n338), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n428), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(new_n426), .B1(new_n395), .B2(new_n396), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n610), .A2(new_n380), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n307), .A2(new_n310), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n299), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n559), .A2(new_n543), .A3(new_n557), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n527), .A2(new_n532), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n615), .A2(KEYINPUT26), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n507), .B1(new_n270), .B2(new_n500), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT88), .B1(new_n617), .B2(G169), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n509), .A2(new_n619), .A3(new_n296), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(new_n513), .A3(new_n523), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n509), .A2(G200), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n529), .A2(new_n531), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n614), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(KEYINPUT26), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n616), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n496), .A2(new_n598), .A3(new_n601), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n541), .A2(new_n542), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n563), .B1(new_n629), .B2(G200), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n566), .A2(new_n557), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n614), .B1(new_n632), .B2(new_n564), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n622), .A2(new_n624), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n574), .A2(new_n575), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n628), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n627), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n438), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n613), .A2(new_n638), .ZN(G369));
  NAND2_X1  g0439(.A1(new_n598), .A2(new_n601), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n289), .A2(G20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n242), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT89), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT27), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(G213), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G343), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n640), .A2(new_n585), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n585), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n604), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n575), .A2(new_n649), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n496), .B1(new_n576), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n650), .A2(new_n496), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n650), .B1(new_n598), .B2(new_n601), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n659), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n210), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n224), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  AOI211_X1 g0474(.A(KEYINPUT29), .B(new_n650), .C1(new_n627), .C2(new_n636), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n625), .A2(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n527), .A2(new_n532), .A3(new_n614), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n622), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT91), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT91), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n676), .A2(new_n682), .A3(new_n622), .A4(new_n679), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n636), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n622), .A2(new_n624), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n568), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(KEYINPUT92), .A3(new_n635), .A4(new_n628), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n649), .B1(new_n684), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n675), .B1(new_n691), .B2(KEYINPUT29), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n605), .A2(new_n569), .A3(new_n649), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n454), .B1(new_n462), .B2(new_n249), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n629), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n526), .A3(new_n600), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n629), .A2(new_n463), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n617), .A2(G179), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n700), .A2(new_n701), .A3(new_n592), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n700), .B2(new_n592), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n695), .A2(new_n526), .A3(KEYINPUT30), .A4(new_n600), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n650), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n650), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n693), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n692), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n674), .B1(new_n717), .B2(G1), .ZN(G364));
  AOI21_X1  g0518(.A(new_n242), .B1(new_n641), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n669), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT94), .Z(new_n726));
  OR2_X1    g0526(.A1(new_n654), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n279), .A2(new_n331), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n337), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n279), .A2(G190), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(G58), .A2(new_n731), .B1(new_n734), .B2(G77), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n337), .A2(new_n389), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n728), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n404), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT96), .Z(new_n739));
  NAND2_X1  g0539(.A1(new_n337), .A2(G200), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT97), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n742), .A2(new_n279), .A3(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G107), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n742), .A2(new_n279), .A3(new_n331), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G87), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n736), .A2(new_n732), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n266), .B1(new_n747), .B2(new_n398), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n279), .B1(new_n749), .B2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n748), .B1(G97), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n732), .A2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(G159), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT32), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n744), .A2(new_n746), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n747), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT33), .B(G317), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n758), .A2(new_n759), .B1(new_n731), .B2(G322), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT98), .Z(new_n761));
  AOI22_X1  g0561(.A1(G283), .A2(new_n743), .B1(new_n745), .B2(G303), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n751), .A2(G294), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n266), .B1(new_n734), .B2(G311), .ZN(new_n764));
  INV_X1    g0564(.A(new_n737), .ZN(new_n765));
  INV_X1    g0565(.A(new_n753), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n765), .A2(G326), .B1(new_n766), .B2(G329), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n739), .A2(new_n757), .B1(new_n761), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n221), .B1(G20), .B2(new_n296), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n726), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n773), .ZN(new_n775));
  XOR2_X1   g0575(.A(G355), .B(KEYINPUT93), .Z(new_n776));
  NOR2_X1   g0576(.A1(new_n668), .A2(new_n264), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n776), .A2(new_n777), .B1(new_n577), .B2(new_n668), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n224), .A2(G45), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n668), .A2(new_n266), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(new_n237), .C2(new_n445), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n769), .A2(new_n773), .B1(new_n775), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n722), .B1(new_n727), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n654), .B(G330), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(new_n722), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT99), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  AOI21_X1  g0588(.A(new_n650), .B1(new_n627), .B2(new_n636), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n650), .A2(new_n323), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n340), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n339), .A2(new_n338), .A3(new_n323), .A4(new_n650), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n789), .B(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n715), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n721), .B1(new_n715), .B2(new_n794), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n773), .A2(new_n723), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n722), .B1(new_n798), .B2(new_n204), .ZN(new_n799));
  INV_X1    g0599(.A(new_n773), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n264), .B1(new_n737), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G294), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n730), .A2(new_n803), .B1(new_n753), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n802), .B(new_n805), .C1(G97), .C2(new_n751), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n745), .A2(G107), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n747), .A2(new_n808), .B1(new_n733), .B2(new_n577), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT100), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n743), .A2(G87), .ZN(new_n811));
  AND4_X1   g0611(.A1(new_n806), .A2(new_n807), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G143), .A2(new_n731), .B1(new_n734), .B2(G159), .ZN(new_n813));
  INV_X1    g0613(.A(G137), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n814), .B2(new_n737), .C1(new_n284), .C2(new_n747), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT34), .ZN(new_n816));
  INV_X1    g0616(.A(G58), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n266), .B1(new_n750), .B2(new_n817), .C1(new_n818), .C2(new_n753), .ZN(new_n819));
  INV_X1    g0619(.A(new_n743), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n398), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(G50), .C2(new_n745), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n812), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n799), .B1(new_n800), .B2(new_n823), .C1(new_n793), .C2(new_n724), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT101), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n797), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  OAI21_X1  g0627(.A(G77), .B1(new_n817), .B2(new_n398), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n828), .A2(new_n224), .B1(G50), .B2(new_n398), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n829), .A2(G1), .A3(new_n289), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT102), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n577), .B(new_n223), .C1(new_n553), .C2(KEYINPUT35), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(KEYINPUT35), .B2(new_n553), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT36), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n608), .A2(new_n649), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n789), .B2(new_n793), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n650), .A2(new_n411), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n426), .A2(new_n428), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n411), .B(new_n650), .C1(new_n424), .C2(new_n425), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n388), .A2(new_n391), .A3(new_n345), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n471), .B1(new_n386), .B2(new_n352), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n322), .A2(new_n281), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n846), .A2(new_n847), .B1(new_n848), .B2(new_n344), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n845), .B1(new_n647), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n369), .B2(new_n375), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT37), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n648), .A2(new_n363), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n363), .A2(new_n376), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n853), .A2(new_n845), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n849), .A2(new_n647), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n857), .B1(new_n397), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(KEYINPUT38), .B(new_n857), .C1(new_n397), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n844), .A2(new_n864), .B1(new_n380), .B2(new_n647), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n426), .A2(new_n650), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n862), .B2(new_n863), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n853), .A2(new_n845), .A3(new_n854), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(new_n855), .ZN(new_n871));
  INV_X1    g0671(.A(new_n393), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n853), .B1(new_n872), .B2(new_n433), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n861), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n863), .A2(new_n874), .A3(new_n868), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT103), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n863), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n436), .A2(new_n858), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n878), .B2(new_n857), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT39), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n863), .A2(new_n874), .A3(new_n868), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n867), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n866), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n613), .ZN(new_n886));
  INV_X1    g0686(.A(new_n692), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n438), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n885), .B(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n711), .A2(new_n842), .A3(new_n793), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n863), .A2(new_n874), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT40), .B1(new_n862), .B2(new_n863), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n892), .A2(KEYINPUT40), .B1(new_n893), .B2(new_n890), .ZN(new_n894));
  INV_X1    g0694(.A(new_n438), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n894), .B1(new_n895), .B2(new_n712), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n890), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n863), .A2(new_n874), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n711), .A2(new_n842), .A3(new_n793), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT40), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n438), .A3(new_n711), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n896), .A2(G330), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n889), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n242), .B2(new_n641), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n889), .A2(new_n903), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n836), .B1(new_n905), .B2(new_n906), .ZN(G367));
  AND2_X1   g0707(.A1(new_n233), .A2(new_n780), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n775), .B1(new_n210), .B2(new_n312), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT46), .ZN(new_n910));
  INV_X1    g0710(.A(new_n745), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n577), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n743), .A2(G97), .ZN(new_n913));
  OAI221_X1 g0713(.A(new_n264), .B1(new_n750), .B2(new_n474), .C1(new_n737), .C2(new_n804), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n803), .A2(new_n747), .B1(new_n730), .B2(new_n801), .ZN(new_n915));
  INV_X1    g0715(.A(G317), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n733), .A2(new_n808), .B1(new_n753), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n745), .A2(KEYINPUT46), .A3(G116), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n912), .A2(new_n913), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n820), .A2(new_n204), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n264), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT109), .ZN(new_n923));
  INV_X1    g0723(.A(G143), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n737), .A2(new_n924), .B1(new_n730), .B2(new_n284), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n750), .A2(new_n398), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT108), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n745), .A2(G58), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n747), .A2(new_n754), .B1(new_n733), .B2(new_n404), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(G137), .B2(new_n766), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n929), .A2(new_n930), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n920), .B1(new_n923), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT47), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n773), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n721), .B1(new_n908), .B2(new_n909), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT110), .Z(new_n940));
  OR2_X1    g0740(.A1(new_n649), .A2(new_n531), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n634), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n622), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n940), .B1(new_n726), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT104), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(KEYINPUT43), .B2(new_n943), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT42), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n661), .A2(new_n665), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n633), .B1(new_n557), .B2(new_n649), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT105), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n650), .A2(new_n614), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n950), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n561), .B1(new_n955), .B2(new_n496), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n649), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n957), .A3(new_n950), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(KEYINPUT106), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n949), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n955), .A2(new_n956), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n664), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n960), .A2(new_n962), .A3(new_n964), .A4(new_n948), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n968), .B1(new_n966), .B2(new_n969), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  INV_X1    g0775(.A(new_n666), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n957), .A2(KEYINPUT45), .A3(new_n666), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n967), .A2(KEYINPUT44), .A3(new_n976), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n957), .B2(new_n666), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(KEYINPUT107), .A3(new_n663), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n663), .A2(KEYINPUT107), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n661), .B(new_n665), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n656), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n717), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n669), .B(KEYINPUT41), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n720), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n944), .B1(new_n974), .B2(new_n994), .ZN(G387));
  OR2_X1    g0795(.A1(new_n716), .A2(new_n990), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n716), .A2(new_n990), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n669), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n990), .A2(new_n719), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n230), .A2(new_n445), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n281), .A2(new_n404), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT50), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n671), .B(new_n445), .C1(new_n398), .C2(new_n204), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n780), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1000), .B1(KEYINPUT111), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(KEYINPUT111), .B2(new_n1004), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n777), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(G107), .B2(new_n210), .C1(new_n671), .C2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n722), .B1(new_n1008), .B2(new_n775), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n750), .A2(new_n312), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G50), .B2(new_n731), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT112), .Z(new_n1012));
  OAI21_X1  g0812(.A(new_n266), .B1(new_n753), .B2(new_n284), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n747), .A2(new_n282), .B1(new_n733), .B2(new_n398), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G159), .C2(new_n765), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n745), .A2(G77), .ZN(new_n1016));
  AND4_X1   g0816(.A1(new_n913), .A2(new_n1012), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n745), .A2(G294), .B1(G283), .B2(new_n751), .ZN(new_n1018));
  INV_X1    g0818(.A(G322), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n737), .A2(new_n1019), .B1(new_n747), .B2(new_n804), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n730), .A2(new_n916), .B1(new_n733), .B2(new_n801), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1020), .B1(KEYINPUT113), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT113), .B2(new_n1021), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1018), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n266), .B1(new_n766), .B2(G326), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n820), .B2(new_n577), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n1026), .B2(KEYINPUT49), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1017), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1009), .B1(new_n1031), .B2(new_n800), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n662), .B2(new_n774), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n999), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n998), .A2(new_n1034), .ZN(G393));
  NOR2_X1   g0835(.A1(new_n984), .A2(new_n663), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n664), .B1(new_n979), .B2(new_n983), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n996), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n669), .C1(new_n996), .C2(new_n988), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n967), .A2(new_n774), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n775), .B1(new_n518), .B2(new_n210), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n240), .A2(new_n668), .A3(new_n266), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n721), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n737), .A2(new_n916), .B1(new_n730), .B2(new_n804), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT52), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n743), .A2(G107), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1045), .C1(new_n808), .C2(new_n911), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G294), .A2(new_n734), .B1(new_n766), .B2(G322), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n266), .B1(new_n758), .B2(G303), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n577), .C2(new_n750), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G50), .A2(new_n758), .B1(new_n766), .B2(G143), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n264), .B1(new_n734), .B2(new_n281), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n204), .C2(new_n750), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n737), .A2(new_n284), .B1(new_n730), .B2(new_n754), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT51), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n745), .A2(G68), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n811), .C1(new_n1056), .C2(new_n1055), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1048), .A2(new_n1051), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1044), .B1(new_n1059), .B2(new_n773), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1040), .A2(new_n720), .B1(new_n1041), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1039), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT114), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT114), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1039), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(G390));
  NAND3_X1  g0866(.A1(new_n711), .A2(G330), .A3(new_n793), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n843), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n711), .A2(new_n793), .A3(G330), .A4(new_n842), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n838), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n686), .A2(new_n689), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n681), .A2(new_n683), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n650), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n837), .B1(new_n1073), .B2(new_n793), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n438), .A2(new_n714), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n613), .B(new_n1077), .C1(new_n692), .C2(new_n895), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n867), .B1(new_n838), .B2(new_n843), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n876), .A2(new_n883), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n867), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n898), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1074), .B2(new_n843), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1069), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n1082), .A2(new_n1085), .A3(new_n1069), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1080), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1069), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1082), .A2(new_n1085), .A3(new_n1069), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1079), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n669), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1087), .A2(new_n1086), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n876), .A2(new_n883), .A3(new_n723), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n798), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n721), .B1(new_n1097), .B2(new_n281), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n747), .A2(new_n474), .B1(new_n753), .B2(new_n803), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n746), .B1(new_n820), .B2(new_n398), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n737), .A2(new_n808), .B1(new_n733), .B2(new_n518), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n264), .B1(new_n750), .B2(new_n204), .C1(new_n577), .C2(new_n730), .ZN(new_n1102));
  OR4_X1    g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(G125), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n266), .B1(new_n1104), .B2(new_n753), .C1(new_n820), .C2(new_n404), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT116), .Z(new_n1106));
  NOR2_X1   g0906(.A1(new_n747), .A2(new_n814), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n737), .A2(new_n1108), .B1(new_n730), .B2(new_n818), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1107), .B(new_n1109), .C1(G159), .C2(new_n751), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT115), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n745), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT53), .B1(new_n745), .B2(G150), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1110), .B1(new_n733), .B2(new_n1113), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1103), .B1(new_n1106), .B2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1117), .A2(KEYINPUT117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(new_n773), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(KEYINPUT117), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1098), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1095), .A2(new_n720), .B1(new_n1096), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1094), .A2(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(KEYINPUT119), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1078), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n612), .A2(new_n298), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n648), .A2(new_n295), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n311), .A2(new_n1129), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1127), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n311), .A2(new_n1129), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n1126), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n713), .B(new_n1137), .C1(new_n897), .C2(new_n900), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1137), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n901), .B2(G330), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1138), .A2(new_n1140), .B1(new_n884), .B2(new_n866), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1137), .B1(new_n894), .B2(new_n713), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n901), .A2(G330), .A3(new_n1139), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n876), .A2(new_n883), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1083), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .A4(new_n865), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1093), .A2(new_n1125), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1124), .B1(new_n1147), .B2(KEYINPUT57), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT57), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1078), .B1(new_n1095), .B2(new_n1079), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1151));
  OAI211_X1 g0951(.A(KEYINPUT119), .B(new_n1149), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1093), .A2(new_n1125), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT118), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1141), .A2(new_n1146), .A3(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(KEYINPUT118), .B1(new_n866), .B2(new_n884), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(KEYINPUT57), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1148), .A2(new_n1152), .A3(new_n669), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1151), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1137), .A2(new_n723), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n721), .B1(new_n1097), .B2(G50), .ZN(new_n1161));
  INV_X1    g0961(.A(G41), .ZN(new_n1162));
  AOI21_X1  g0962(.A(G50), .B1(new_n260), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G58), .A2(new_n743), .B1(new_n745), .B2(G77), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n765), .A2(G116), .B1(new_n766), .B2(G283), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G107), .A2(new_n731), .B1(new_n734), .B2(new_n313), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1162), .B(new_n264), .C1(new_n747), .C2(new_n518), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(new_n926), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT58), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1163), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n747), .A2(new_n818), .B1(new_n733), .B2(new_n814), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n737), .A2(new_n1104), .B1(new_n730), .B2(new_n1108), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(G150), .C2(new_n751), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n911), .B2(new_n1113), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n743), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1171), .B1(new_n1170), .B2(new_n1169), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1161), .B1(new_n1181), .B2(new_n773), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1159), .A2(new_n720), .B1(new_n1160), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1158), .A2(new_n1183), .ZN(G375));
  NOR2_X1   g0984(.A1(new_n1076), .A2(new_n719), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT120), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT120), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n722), .B1(new_n798), .B2(new_n398), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n745), .A2(G97), .B1(G303), .B2(new_n766), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT121), .Z(new_n1190));
  AOI22_X1  g0990(.A1(G283), .A2(new_n731), .B1(new_n734), .B2(G107), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n577), .B2(new_n747), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n264), .B1(new_n737), .B2(new_n803), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n921), .A2(new_n1192), .A3(new_n1010), .A4(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n817), .A2(new_n820), .B1(new_n911), .B2(new_n754), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n758), .B2(new_n1112), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n730), .A2(new_n814), .B1(new_n753), .B2(new_n1108), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n266), .B1(new_n750), .B2(new_n404), .C1(new_n284), .C2(new_n733), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(G132), .C2(new_n765), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1190), .A2(new_n1194), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1188), .B1(new_n800), .B2(new_n1200), .C1(new_n842), .C2(new_n724), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1186), .A2(new_n1187), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1080), .A2(new_n993), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(G381));
  AND2_X1   g1006(.A1(new_n991), .A2(new_n993), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n973), .B1(new_n1207), .B2(new_n720), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1208), .A2(new_n1063), .A3(new_n944), .A4(new_n1065), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n998), .A2(new_n787), .A3(new_n1034), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1209), .A2(G384), .A3(G381), .A4(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G378), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1158), .A2(new_n1212), .A3(new_n1183), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT122), .ZN(G407));
  OAI211_X1 g1016(.A(G407), .B(G213), .C1(G343), .C2(new_n1213), .ZN(G409));
  NAND2_X1  g1017(.A1(G390), .A2(G387), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(G393), .B(new_n787), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1218), .A2(new_n1209), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1218), .B2(new_n1209), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1155), .A2(new_n720), .A3(new_n1156), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1160), .A2(new_n1182), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1223), .A2(new_n1094), .A3(new_n1122), .A4(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1150), .A2(new_n1151), .A3(new_n992), .ZN(new_n1226));
  INV_X1    g1026(.A(G213), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1225), .A2(new_n1226), .B1(new_n1227), .B2(G343), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G375), .B2(G378), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1230));
  OR2_X1    g1030(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT60), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1204), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1078), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n669), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT123), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1233), .A2(new_n1237), .A3(new_n669), .A4(new_n1234), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(G384), .B1(new_n1239), .B2(new_n1203), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n826), .B(new_n1202), .C1(new_n1236), .C2(new_n1238), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  INV_X1    g1044(.A(G2897), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G343), .B(new_n1227), .C1(KEYINPUT124), .C2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(KEYINPUT124), .B2(new_n1245), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1242), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1212), .B1(new_n1158), .B2(new_n1183), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n1228), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1227), .A2(new_n1245), .A3(G343), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT125), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1254), .B(new_n1251), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1243), .B(new_n1244), .C1(new_n1250), .C2(new_n1256), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(new_n1249), .A2(new_n1228), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1230), .B1(new_n1258), .B2(new_n1231), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1222), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT63), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1229), .A2(new_n1242), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1222), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1229), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1264), .A2(new_n1248), .A3(new_n1253), .A4(new_n1255), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1258), .A2(KEYINPUT63), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1263), .A2(new_n1244), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1260), .A2(new_n1267), .ZN(G405));
  INV_X1    g1068(.A(new_n1249), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1242), .A2(KEYINPUT127), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1213), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT127), .B(new_n1242), .C1(new_n1214), .C2(new_n1249), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1273), .B(new_n1222), .Z(G402));
endmodule


