//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  OR2_X1    g0017(.A1(KEYINPUT65), .A2(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(KEYINPUT65), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n220), .A2(G1), .A3(G13), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n214), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n217), .B1(new_n221), .B2(new_n222), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G68), .Z(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G232), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G1698), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n251), .B1(G226), .B2(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT69), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n254), .A2(new_n261), .A3(new_n255), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT13), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT66), .A2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n211), .B(G274), .C1(new_n258), .C2(new_n259), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  OAI211_X1 g0074(.A(G1), .B(G13), .C1(new_n274), .C2(new_n266), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n271), .A2(new_n273), .B1(new_n278), .B2(G238), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n263), .A2(new_n264), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n264), .B1(new_n263), .B2(new_n279), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G190), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n263), .A2(new_n279), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n263), .A2(new_n264), .A3(new_n279), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G200), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n259), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n211), .B2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G68), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT70), .ZN(new_n293));
  INV_X1    g0093(.A(new_n290), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n220), .A2(new_n274), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G77), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n224), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n293), .B1(KEYINPUT11), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT11), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n224), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT12), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n283), .A2(new_n288), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT14), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(G169), .C1(new_n280), .C2(new_n281), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT71), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n287), .A2(KEYINPUT71), .A3(new_n310), .A4(G169), .ZN(new_n314));
  OAI21_X1  g0114(.A(G169), .B1(new_n280), .B2(new_n281), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n282), .A2(G179), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n313), .A2(new_n314), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n307), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n309), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(KEYINPUT67), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n295), .A3(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n297), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n294), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n303), .A2(new_n202), .ZN(new_n327));
  INV_X1    g0127(.A(new_n291), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n202), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT9), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n252), .A2(new_n253), .ZN(new_n332));
  INV_X1    g0132(.A(G1698), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G223), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT3), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n274), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G222), .A3(new_n333), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n332), .A2(G77), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n260), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n271), .A2(new_n273), .B1(new_n278), .B2(G226), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G200), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(G190), .A3(new_n344), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT9), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n326), .B2(new_n329), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n331), .A2(new_n346), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT10), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n349), .A2(new_n347), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT10), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(new_n331), .A4(new_n346), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n330), .B1(new_n356), .B2(new_n345), .ZN(new_n357));
  INV_X1    g0157(.A(G179), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n343), .A2(new_n358), .A3(new_n344), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G77), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n303), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n328), .B2(new_n361), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n295), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(KEYINPUT65), .A2(G20), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT65), .A2(G20), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n297), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n366), .B1(new_n361), .B2(new_n369), .C1(new_n370), .C2(new_n321), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n363), .B1(new_n371), .B2(new_n290), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G232), .A2(G1698), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n225), .B2(G1698), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n332), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n260), .B1(new_n339), .B2(G107), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G244), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n270), .A2(new_n272), .B1(new_n277), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT68), .ZN(new_n380));
  OR3_X1    g0180(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n377), .B2(new_n379), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n372), .B1(new_n383), .B2(new_n358), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n356), .A3(new_n382), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(G200), .A3(new_n382), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n387), .A2(new_n372), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n383), .A2(G190), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AND4_X1   g0190(.A1(new_n355), .A2(new_n360), .A3(new_n386), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n322), .A2(new_n323), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n302), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT67), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n321), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n328), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n275), .A2(G232), .A3(new_n276), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(new_n270), .C2(new_n272), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(G223), .A2(G1698), .ZN(new_n402));
  INV_X1    g0202(.A(G226), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n339), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT73), .A3(new_n260), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n404), .A2(new_n339), .B1(G33), .B2(G87), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n275), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n401), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G200), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n275), .B1(new_n405), .B2(new_n406), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n398), .B1(new_n270), .B2(new_n272), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT16), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n369), .B2(new_n332), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT7), .A4(G20), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n420), .A2(new_n421), .A3(new_n224), .ZN(new_n422));
  AND2_X1   g0222(.A1(G58), .A2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(G20), .B1(new_n423), .B2(new_n201), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n297), .A2(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n418), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n290), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n369), .A2(new_n332), .A3(new_n419), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n337), .A2(new_n212), .A3(new_n338), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT7), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n431), .A3(G68), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n424), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n432), .B2(new_n434), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n397), .B(new_n417), .C1(new_n428), .C2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n397), .B1(new_n428), .B2(new_n437), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n398), .B(new_n358), .C1(new_n270), .C2(new_n272), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(new_n408), .A3(new_n411), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n356), .B1(new_n414), .B2(new_n415), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n441), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n397), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n432), .A2(new_n434), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT72), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT7), .B1(new_n220), .B2(new_n339), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n332), .A2(new_n419), .A3(new_n212), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(G68), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n426), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n294), .B1(new_n459), .B2(new_n418), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n450), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n461), .A2(KEYINPUT18), .A3(new_n447), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT74), .B1(new_n449), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n442), .A2(new_n441), .A3(new_n448), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT18), .B1(new_n461), .B2(new_n447), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT74), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n440), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n320), .A2(new_n391), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT5), .B1(new_n267), .B2(new_n268), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n211), .B(G45), .C1(new_n472), .C2(G41), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(G274), .A3(new_n275), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(new_n275), .C1(new_n471), .C2(new_n473), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(G244), .B(new_n333), .C1(new_n252), .C2(new_n253), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT77), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n334), .A2(G250), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n479), .A2(new_n480), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n482), .A2(new_n483), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n487), .A2(KEYINPUT78), .A3(new_n260), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT78), .B1(new_n487), .B2(new_n260), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G200), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n211), .A2(G33), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n302), .A2(new_n492), .A3(new_n259), .A4(new_n289), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT76), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G97), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n303), .A2(new_n205), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g0300(.A(G97), .B(G107), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n502), .A2(new_n205), .A3(G107), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(new_n220), .B1(G77), .B2(new_n297), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n455), .A2(G107), .A3(new_n456), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n294), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n420), .A2(new_n421), .A3(new_n206), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n504), .B1(new_n502), .B2(new_n501), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n512), .A2(new_n369), .B1(new_n361), .B2(new_n370), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n290), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT75), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n500), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n477), .B1(new_n487), .B2(new_n260), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n491), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n498), .A2(new_n499), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n522));
  AOI211_X1 g0322(.A(new_n515), .B(new_n294), .C1(new_n507), .C2(new_n508), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n518), .A2(G169), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n526), .C1(new_n490), .C2(G179), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n520), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT19), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n255), .A2(new_n529), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n220), .A2(new_n530), .B1(G87), .B2(new_n207), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n218), .A2(G33), .A3(G97), .A4(new_n219), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n529), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n339), .A2(new_n369), .A3(G68), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n290), .B1(new_n303), .B2(new_n364), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n495), .A2(G87), .A3(new_n496), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G45), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n227), .B1(new_n539), .B2(G1), .ZN(new_n540));
  INV_X1    g0340(.A(G274), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n211), .A2(new_n541), .A3(G45), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n275), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n339), .A2(G238), .A3(new_n333), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n548), .B2(new_n260), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G190), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT79), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT79), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n552), .A3(G190), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n260), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n543), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n538), .A2(new_n551), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n495), .A2(new_n496), .A3(new_n365), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n536), .A2(new_n558), .B1(new_n549), .B2(new_n358), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G169), .B2(new_n549), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n339), .A2(G257), .A3(G1698), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n339), .A2(G250), .A3(new_n333), .ZN(new_n563));
  XNOR2_X1  g0363(.A(KEYINPUT84), .B(G294), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G33), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n260), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n471), .A2(new_n473), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G264), .A3(new_n275), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n569), .A3(new_n475), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n356), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n567), .A2(new_n569), .A3(new_n358), .A4(new_n475), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT83), .ZN(new_n575));
  AOI211_X1 g0375(.A(KEYINPUT23), .B(G107), .C1(new_n218), .C2(new_n219), .ZN(new_n576));
  NAND2_X1  g0376(.A1(KEYINPUT23), .A2(G107), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(G20), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n575), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n220), .A2(new_n581), .A3(new_n206), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n578), .A2(G20), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n582), .A2(KEYINPUT83), .A3(new_n583), .A4(new_n577), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n339), .A2(new_n369), .A3(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT22), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT22), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n339), .A2(new_n369), .A3(new_n588), .A4(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g0391(.A(KEYINPUT82), .B(KEYINPUT24), .Z(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n592), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n585), .A2(new_n594), .A3(new_n590), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n294), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n497), .A2(G107), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n303), .A2(new_n206), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT25), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n574), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n595), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n594), .B1(new_n585), .B2(new_n590), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n290), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n570), .A2(new_n413), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G190), .B2(new_n570), .ZN(new_n607));
  INV_X1    g0407(.A(new_n601), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n561), .A2(new_n602), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n369), .B(new_n483), .C1(G33), .C2(new_n205), .ZN(new_n612));
  INV_X1    g0412(.A(G116), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n289), .A2(new_n259), .B1(G20), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(KEYINPUT20), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT81), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n612), .A2(KEYINPUT81), .A3(KEYINPUT20), .A4(new_n614), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n612), .A2(new_n614), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n617), .B(new_n618), .C1(KEYINPUT20), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT80), .ZN(new_n621));
  OR3_X1    g0421(.A1(new_n493), .A2(new_n621), .A3(new_n613), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n493), .B2(new_n613), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(new_n613), .B2(new_n303), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n339), .A2(G264), .A3(G1698), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n339), .A2(G257), .A3(new_n333), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n332), .A2(G303), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n260), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n568), .A2(G270), .A3(new_n275), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n475), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G169), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n611), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(G200), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n632), .A2(new_n399), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n625), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n620), .A2(new_n624), .ZN(new_n638));
  AND4_X1   g0438(.A1(G179), .A2(new_n630), .A3(new_n475), .A4(new_n631), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n638), .A2(KEYINPUT21), .A3(G169), .A4(new_n632), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n634), .A2(new_n637), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n528), .A2(new_n610), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n470), .A2(new_n643), .ZN(G372));
  INV_X1    g0444(.A(KEYINPUT86), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n449), .B2(new_n462), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT86), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n318), .A2(new_n319), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(new_n386), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n438), .B(KEYINPUT17), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n308), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n648), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n653), .A2(new_n355), .B1(new_n359), .B2(new_n357), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n555), .A2(KEYINPUT85), .A3(new_n356), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT85), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n549), .B2(G169), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n559), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n538), .A2(new_n550), .A3(new_n556), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n520), .A2(new_n662), .A3(new_n527), .A4(new_n609), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n573), .B1(new_n605), .B2(new_n608), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n659), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n527), .B2(new_n661), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n517), .A2(new_n525), .ZN(new_n670));
  INV_X1    g0470(.A(new_n489), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n487), .A2(KEYINPUT78), .A3(new_n260), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n477), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n358), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n561), .A2(new_n670), .A3(KEYINPUT26), .A4(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n470), .B1(new_n667), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n654), .A2(new_n677), .ZN(G369));
  NAND3_X1  g0478(.A1(new_n369), .A2(new_n211), .A3(G13), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n625), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n664), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n642), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n609), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n665), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n684), .B1(new_n596), .B2(new_n601), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n665), .A2(new_n684), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n690), .A2(KEYINPUT87), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT87), .ZN(new_n698));
  INV_X1    g0498(.A(new_n696), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n689), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n664), .A2(new_n685), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n702), .A2(new_n692), .B1(new_n665), .B2(new_n685), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(KEYINPUT89), .ZN(new_n705));
  INV_X1    g0505(.A(new_n215), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n269), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n215), .A2(KEYINPUT89), .A3(new_n267), .A4(new_n268), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT88), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n222), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n557), .A2(new_n560), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n691), .A2(new_n665), .A3(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n519), .B(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n718), .A2(new_n491), .B1(new_n670), .B2(new_n674), .ZN(new_n719));
  INV_X1    g0519(.A(new_n642), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n716), .A2(new_n719), .A3(new_n720), .A4(new_n685), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n685), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n549), .A2(new_n569), .A3(new_n567), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n639), .A2(new_n724), .A3(KEYINPUT30), .A4(new_n518), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n632), .A2(new_n570), .A3(new_n358), .A4(new_n555), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n639), .A2(new_n724), .A3(new_n518), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT90), .B(KEYINPUT30), .Z(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n490), .A2(new_n727), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT91), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n725), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n727), .A2(new_n490), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n728), .A2(new_n730), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n734), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n723), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n725), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n684), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n722), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n721), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n685), .B1(new_n667), .B2(new_n676), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(KEYINPUT92), .B(new_n668), .C1(new_n527), .C2(new_n715), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n662), .A2(KEYINPUT26), .A3(new_n674), .A4(new_n670), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n561), .A2(new_n670), .A3(new_n674), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT92), .B1(new_n749), .B2(new_n668), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT29), .B(new_n685), .C1(new_n751), .C2(new_n667), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n742), .B1(new_n745), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n714), .B1(new_n753), .B2(G1), .ZN(G364));
  INV_X1    g0554(.A(new_n709), .ZN(new_n755));
  INV_X1    g0555(.A(G13), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n220), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n211), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n259), .B1(G20), .B2(new_n356), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n369), .A2(new_n358), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(new_n399), .A3(new_n413), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(KEYINPUT95), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n369), .B1(G190), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n564), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n765), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n413), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G326), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n770), .A2(G311), .B1(new_n779), .B2(KEYINPUT97), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n765), .A2(new_n399), .A3(G200), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n413), .A2(G179), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT96), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n212), .A2(new_n399), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n339), .B1(new_n788), .B2(G303), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n369), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(new_n771), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n792), .A2(G283), .B1(new_n794), .B2(G329), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n783), .A2(new_n789), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n775), .A2(G200), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(G322), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n780), .B(new_n798), .C1(KEYINPUT97), .C2(new_n779), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n792), .A2(G107), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n788), .A2(G87), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n773), .A2(G97), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n800), .A2(new_n801), .A3(new_n339), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n794), .A2(G159), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT32), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n805), .C1(G50), .C2(new_n776), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n797), .A2(G58), .B1(new_n781), .B2(G68), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(new_n361), .C2(new_n769), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n763), .B1(new_n799), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n762), .ZN(new_n813));
  AND2_X1   g0613(.A1(G355), .A2(KEYINPUT93), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G355), .A2(KEYINPUT93), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n215), .A2(new_n339), .ZN(new_n816));
  OR3_X1    g0616(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n248), .A2(new_n539), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n706), .A2(new_n339), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(G45), .B2(new_n222), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n817), .B1(G116), .B2(new_n215), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n761), .B(new_n809), .C1(new_n813), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n812), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n688), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n690), .A2(new_n760), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G330), .B2(new_n688), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  OAI21_X1  g0628(.A(new_n390), .B1(new_n372), .B2(new_n685), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n386), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n384), .A2(new_n385), .A3(new_n685), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n743), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n742), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT98), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT98), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n834), .A2(new_n837), .A3(new_n742), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n761), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT99), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n836), .A2(KEYINPUT99), .A3(new_n761), .A4(new_n838), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(new_n742), .C2(new_n834), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G137), .A2(new_n776), .B1(new_n797), .B2(G143), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  INV_X1    g0645(.A(new_n781), .ZN(new_n846));
  INV_X1    g0646(.A(G159), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n844), .B1(new_n845), .B2(new_n846), .C1(new_n769), .C2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT34), .Z(new_n849));
  OAI21_X1  g0649(.A(new_n339), .B1(new_n787), .B2(new_n202), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n792), .A2(G68), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n794), .A2(G132), .ZN(new_n852));
  INV_X1    g0652(.A(G58), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n772), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n797), .A2(G294), .B1(new_n781), .B2(G283), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n802), .A2(new_n332), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n226), .A2(new_n791), .B1(new_n787), .B2(new_n206), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(G311), .C2(new_n794), .ZN(new_n859));
  INV_X1    g0659(.A(G303), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n856), .B(new_n859), .C1(new_n860), .C2(new_n777), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G116), .B2(new_n770), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n762), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n762), .A2(new_n810), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n761), .B1(new_n361), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n863), .B(new_n865), .C1(new_n811), .C2(new_n833), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n843), .A2(new_n866), .ZN(G384));
  NAND2_X1  g0667(.A1(new_n442), .A2(new_n448), .ZN(new_n868));
  INV_X1    g0668(.A(new_n682), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n442), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .A4(new_n438), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n432), .A2(new_n458), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n418), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(KEYINPUT101), .A3(new_n290), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT101), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT16), .B1(new_n432), .B2(new_n458), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n294), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n454), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n682), .B1(new_n879), .B2(new_n397), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n447), .B1(new_n879), .B2(new_n397), .ZN(new_n881));
  INV_X1    g0681(.A(new_n438), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n872), .B1(new_n883), .B2(new_n871), .ZN(new_n884));
  INV_X1    g0684(.A(new_n880), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n468), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n884), .B(KEYINPUT38), .C1(new_n468), .C2(new_n885), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n440), .B1(new_n646), .B2(new_n647), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n870), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n438), .B1(new_n461), .B2(new_n447), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n461), .A2(new_n682), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT102), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(new_n872), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT102), .B(KEYINPUT37), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT86), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT86), .B1(new_n464), .B2(new_n465), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n651), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(KEYINPUT103), .A3(new_n896), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n894), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n887), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n889), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n891), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n649), .A2(new_n684), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n648), .A2(new_n869), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n319), .A2(new_n684), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n649), .A2(new_n308), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n319), .B(new_n684), .C1(new_n309), .C2(new_n318), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n833), .B(new_n685), .C1(new_n667), .C2(new_n676), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n831), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n888), .A2(new_n889), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n912), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n745), .A2(new_n752), .A3(new_n470), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n654), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n889), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n906), .B2(new_n887), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n832), .B1(new_n915), .B2(new_n916), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n685), .B1(new_n731), .B2(new_n725), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT104), .B1(new_n930), .B2(KEYINPUT31), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n738), .A2(new_n723), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n739), .A2(new_n933), .A3(new_n722), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n721), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n929), .A2(new_n935), .A3(KEYINPUT40), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT105), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT105), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n929), .A2(new_n935), .A3(KEYINPUT40), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n899), .A2(new_n900), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n870), .B1(new_n648), .B2(new_n651), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n940), .B1(new_n941), .B2(KEYINPUT103), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n942), .B2(new_n894), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n938), .B(new_n939), .C1(new_n943), .C2(new_n927), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n921), .A2(new_n935), .A3(new_n929), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n932), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n643), .B2(new_n685), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n931), .A2(new_n934), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n469), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(G330), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n949), .B2(new_n954), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n926), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n926), .A2(new_n956), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(new_n211), .C2(new_n757), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n613), .B(new_n221), .C1(new_n506), .C2(KEYINPUT35), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(KEYINPUT35), .B2(new_n506), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT36), .ZN(new_n962));
  OAI21_X1  g0762(.A(G77), .B1(new_n853), .B2(new_n224), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n963), .A2(new_n222), .B1(G50), .B2(new_n224), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(G1), .A3(new_n756), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT100), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n959), .A2(new_n967), .ZN(G367));
  AOI21_X1  g0768(.A(new_n602), .B1(new_n718), .B2(new_n491), .ZN(new_n969));
  INV_X1    g0769(.A(new_n527), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n685), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n685), .A2(new_n538), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n559), .A3(new_n658), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n661), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n524), .A2(new_n684), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n520), .A2(new_n527), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n670), .A2(new_n674), .A3(new_n684), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AND4_X1   g0779(.A1(KEYINPUT42), .A2(new_n979), .A3(new_n692), .A4(new_n702), .ZN(new_n980));
  AND4_X1   g0780(.A1(new_n664), .A2(new_n602), .A3(new_n609), .A4(new_n685), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT42), .B1(new_n981), .B2(new_n979), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n971), .B(new_n975), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT106), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n971), .B1(new_n980), .B2(new_n982), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n974), .B(KEYINPUT43), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT107), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT107), .B1(new_n987), .B2(new_n988), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n985), .B(new_n986), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n979), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n701), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT108), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n991), .A2(new_n992), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n986), .A2(new_n985), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT108), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n995), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n993), .A2(new_n996), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n703), .B2(new_n979), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n692), .A2(new_n664), .A3(new_n685), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n665), .A2(new_n685), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1004), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n994), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1005), .A2(KEYINPUT110), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT110), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1012), .B(new_n1004), .C1(new_n703), .C2(new_n979), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1008), .B2(new_n994), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1011), .A2(new_n1013), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n701), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n696), .A2(new_n702), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n1006), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(new_n690), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n701), .A2(new_n1011), .A3(new_n1013), .A4(new_n1017), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1023), .A3(new_n753), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n753), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n709), .B(KEYINPUT41), .Z(new_n1027));
  AOI21_X1  g0827(.A(new_n759), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n819), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n813), .B1(new_n215), .B2(new_n364), .C1(new_n1029), .C2(new_n241), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n760), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n788), .A2(G116), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT46), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n339), .B1(new_n792), .B2(G97), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n794), .A2(G317), .B1(new_n773), .B2(G107), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G303), .B2(new_n797), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n776), .A2(G311), .B1(new_n781), .B2(new_n564), .ZN(new_n1038));
  INV_X1    g0838(.A(G283), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1037), .B(new_n1038), .C1(new_n1039), .C2(new_n769), .ZN(new_n1040));
  INV_X1    g0840(.A(G137), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n339), .B1(new_n793), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n773), .A2(G68), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n787), .B2(new_n853), .C1(new_n361), .C2(new_n791), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(G159), .C2(new_n781), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G143), .A2(new_n776), .B1(new_n797), .B2(G150), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n202), .C2(new_n769), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1040), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT47), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1031), .B1(new_n1049), .B2(new_n762), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT111), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n974), .A2(new_n823), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1003), .A2(new_n1028), .B1(new_n1051), .B2(new_n1052), .ZN(G387));
  NAND2_X1  g0853(.A1(new_n797), .A2(G317), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(KEYINPUT113), .B(G322), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n776), .A2(new_n1056), .B1(new_n781), .B2(G311), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1054), .B(new_n1057), .C1(new_n769), .C2(new_n860), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n788), .A2(new_n564), .B1(new_n773), .B2(G283), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT49), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT114), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n332), .B1(new_n793), .B2(new_n778), .C1(new_n791), .C2(new_n613), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n788), .A2(G77), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n773), .A2(new_n365), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n845), .C2(new_n793), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n332), .B(new_n1072), .C1(G97), .C2(new_n792), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n797), .A2(G50), .B1(new_n781), .B2(new_n395), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n847), .C2(new_n777), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G68), .B2(new_n770), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n762), .B1(new_n1069), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n696), .A2(new_n823), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n711), .A2(new_n816), .B1(G107), .B2(new_n215), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT112), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n321), .A2(G50), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT50), .ZN(new_n1082));
  AOI21_X1  g0882(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n711), .A3(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n819), .C1(new_n238), .C2(new_n539), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n761), .B(new_n1078), .C1(new_n813), .C2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1077), .A2(new_n1087), .B1(new_n759), .B2(new_n1023), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n709), .B1(new_n1023), .B2(new_n753), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n753), .B2(new_n1023), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(G393));
  NAND2_X1  g0891(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1023), .A2(new_n753), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n1025), .A3(new_n755), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1020), .A2(new_n759), .A3(new_n1024), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n813), .B1(new_n205), .B2(new_n215), .C1(new_n1029), .C2(new_n245), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n760), .A2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G311), .A2(new_n797), .B1(new_n776), .B2(G317), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT52), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n793), .A2(new_n1055), .B1(new_n772), .B2(new_n613), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G283), .B2(new_n788), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1102), .A2(new_n332), .A3(new_n800), .ZN(new_n1103));
  INV_X1    g0903(.A(G294), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1103), .B1(new_n860), .B2(new_n846), .C1(new_n769), .C2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G150), .A2(new_n776), .B1(new_n797), .B2(G159), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT51), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n339), .B1(new_n791), .B2(new_n226), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n794), .A2(G143), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n773), .A2(G77), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n224), .C2(new_n787), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1108), .B(new_n1111), .C1(new_n781), .C2(G50), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n321), .B2(new_n769), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1100), .A2(new_n1105), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1098), .B1(new_n1114), .B2(new_n762), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n823), .B2(new_n979), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1096), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1095), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT115), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT115), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1095), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(G390));
  OAI211_X1 g0922(.A(new_n685), .B(new_n830), .C1(new_n751), .C2(new_n667), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n831), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n917), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n911), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n908), .ZN(new_n1127));
  INV_X1    g0927(.A(G330), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n832), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n741), .A2(new_n917), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n920), .A2(new_n911), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1127), .B(new_n1131), .C1(new_n910), .C2(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n920), .A2(new_n911), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n890), .B1(new_n928), .B2(KEYINPUT39), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n928), .A2(new_n911), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1134), .A2(new_n1135), .B1(new_n1125), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n935), .A2(new_n917), .A3(new_n1129), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1133), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(new_n758), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n864), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n776), .A2(G128), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n781), .A2(G137), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n332), .B1(new_n792), .B2(G50), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n787), .A2(new_n845), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n794), .A2(G125), .B1(new_n773), .B2(G159), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1142), .B(new_n1148), .C1(G132), .C2(new_n797), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n770), .A2(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n777), .A2(new_n1039), .B1(new_n846), .B2(new_n206), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n797), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n613), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n801), .A2(new_n332), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n851), .B(new_n1110), .C1(new_n1104), .C2(new_n793), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n770), .A2(G97), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1149), .A2(new_n1152), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n760), .B1(new_n395), .B2(new_n1141), .C1(new_n1160), .C2(new_n763), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1135), .B2(new_n810), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT117), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1140), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1124), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n917), .B1(new_n935), .B2(new_n1129), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1130), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n741), .A2(new_n1129), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n918), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1138), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n919), .A2(new_n831), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1165), .A2(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT116), .B1(new_n953), .B2(G330), .ZN(new_n1173));
  AND4_X1   g0973(.A1(KEYINPUT116), .A2(new_n470), .A3(G330), .A4(new_n935), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n654), .B(new_n924), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1139), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1176), .B(new_n1133), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n755), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1164), .A2(new_n1180), .ZN(G378));
  AOI21_X1  g0981(.A(new_n1128), .B1(new_n946), .B2(new_n947), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n355), .A2(new_n360), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n330), .A2(new_n682), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1183), .B(new_n1184), .Z(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1185), .B(new_n1186), .Z(new_n1187));
  AND3_X1   g0987(.A1(new_n945), .A2(new_n1182), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n945), .B2(new_n1182), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n923), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n938), .B1(new_n908), .B2(new_n939), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n928), .A2(KEYINPUT105), .A3(new_n936), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1182), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1187), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n912), .A2(new_n922), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n945), .A2(new_n1182), .A3(new_n1187), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1190), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1187), .A2(new_n810), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n760), .B1(G50), .B2(new_n1141), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n339), .A2(new_n269), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G50), .B(new_n1202), .C1(new_n274), .C2(new_n266), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1154), .A2(new_n206), .B1(new_n846), .B2(new_n205), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G116), .B2(new_n776), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT118), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1070), .A2(new_n1206), .A3(new_n1202), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n792), .A2(G58), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1043), .C1(new_n1039), .C2(new_n793), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1206), .B1(new_n1070), .B2(new_n1202), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1205), .B(new_n1211), .C1(new_n364), .C2(new_n769), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT58), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1203), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT119), .B(G124), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n274), .B(new_n266), .C1(new_n793), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G159), .B2(new_n792), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n776), .A2(G125), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n797), .A2(G128), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n788), .A2(new_n1151), .B1(new_n773), .B2(G150), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n781), .A2(G132), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G137), .B2(new_n770), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT59), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1223), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1214), .B1(new_n1213), .B2(new_n1212), .C1(new_n1225), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1201), .B1(new_n1228), .B2(new_n762), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1199), .A2(new_n759), .B1(new_n1200), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1175), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1190), .A2(new_n1198), .B1(new_n1179), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n755), .B1(new_n1232), .B2(KEYINPUT57), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT120), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1190), .A2(new_n1198), .A3(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n923), .B(KEYINPUT120), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT57), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1179), .B2(new_n1231), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1230), .B1(new_n1233), .B2(new_n1239), .ZN(G375));
  NAND2_X1  g1040(.A1(new_n1167), .A2(new_n1165), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1231), .A2(new_n1243), .A3(KEYINPUT121), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT121), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n1027), .A3(new_n1177), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1243), .A2(new_n759), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n760), .B1(G68), .B2(new_n1141), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1071), .B1(new_n793), .B2(new_n860), .C1(new_n787), .C2(new_n205), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n339), .B(new_n1251), .C1(G77), .C2(new_n792), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G283), .A2(new_n797), .B1(new_n776), .B2(G294), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(new_n613), .C2(new_n846), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n769), .A2(new_n206), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1208), .A2(KEYINPUT122), .A3(new_n339), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n794), .A2(G128), .B1(new_n773), .B2(G50), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n847), .B2(new_n787), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT122), .B1(new_n1208), .B2(new_n339), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1256), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G132), .A2(new_n776), .B1(new_n797), .B2(G137), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n846), .C2(new_n1150), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n769), .A2(new_n845), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n1254), .A2(new_n1255), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1250), .B1(new_n1264), .B2(new_n762), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n917), .B2(new_n811), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1248), .A2(new_n1268), .ZN(G381));
  NOR2_X1   g1069(.A1(G381), .A2(G390), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n843), .A2(new_n866), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n997), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1028), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1270), .A2(new_n1271), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  OR3_X1    g1077(.A1(new_n1277), .A2(G375), .A3(G378), .ZN(G407));
  INV_X1    g1078(.A(G378), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n683), .A2(G213), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G407), .B(G213), .C1(G375), .C2(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(KEYINPUT123), .ZN(G409));
  OAI211_X1 g1084(.A(G378), .B(new_n1230), .C1(new_n1233), .C2(new_n1239), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1235), .A2(new_n759), .A3(new_n1236), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1200), .A2(new_n1229), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1179), .A2(new_n1231), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1199), .A2(new_n1027), .A3(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1279), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1285), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1172), .A2(new_n1175), .A3(KEYINPUT60), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n755), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1177), .A2(KEYINPUT60), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1247), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1271), .B1(new_n1267), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1247), .A2(new_n1295), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1294), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(G384), .A3(new_n1268), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1292), .A2(new_n1280), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT125), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1281), .B1(new_n1285), .B2(new_n1291), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(KEYINPUT125), .A3(new_n1304), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1275), .A2(G390), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(G387), .A2(new_n1121), .A3(new_n1119), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n827), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1276), .A2(new_n1314), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(G2897), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1280), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1302), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1320), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1297), .A2(new_n1301), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1311), .B(new_n1318), .C1(new_n1308), .C2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1302), .ZN(new_n1327));
  AOI211_X1 g1127(.A(KEYINPUT124), .B(KEYINPUT63), .C1(new_n1308), .C2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT124), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1292), .A2(new_n1280), .A3(new_n1327), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(new_n1303), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1310), .B(new_n1326), .C1(new_n1328), .C2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1292), .A2(new_n1280), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1323), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1322), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1333), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1308), .A2(new_n1338), .A3(new_n1327), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1330), .A2(KEYINPUT62), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1337), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT126), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1342), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1315), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1346), .A2(KEYINPUT126), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT127), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1343), .A2(new_n1348), .A3(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1349), .B1(new_n1343), .B2(new_n1348), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1341), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1332), .A2(new_n1353), .ZN(G405));
  AND2_X1   g1154(.A1(G375), .A2(new_n1279), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1285), .ZN(new_n1356));
  OR3_X1    g1156(.A1(new_n1355), .A2(new_n1356), .A3(new_n1327), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1327), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1343), .A2(new_n1348), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1357), .A2(new_n1348), .A3(new_n1343), .A4(new_n1358), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(G402));
endmodule


