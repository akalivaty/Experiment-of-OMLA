

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  BUF_X1 U553 ( .A(n696), .Z(n697) );
  INV_X1 U554 ( .A(KEYINPUT28), .ZN(n597) );
  AND2_X1 U555 ( .A1(n686), .A2(n685), .ZN(n691) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n695) );
  XNOR2_X2 U557 ( .A(KEYINPUT66), .B(n534), .ZN(n607) );
  XOR2_X1 U558 ( .A(KEYINPUT29), .B(n637), .Z(n515) );
  INV_X1 U559 ( .A(n648), .ZN(n639) );
  INV_X1 U560 ( .A(n924), .ZN(n681) );
  NOR2_X1 U561 ( .A1(n681), .A2(n735), .ZN(n682) );
  NAND2_X2 U562 ( .A1(n695), .A2(n693), .ZN(n648) );
  INV_X1 U563 ( .A(KEYINPUT33), .ZN(n685) );
  NOR2_X1 U564 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U565 ( .A1(n784), .A2(G54), .ZN(n601) );
  NAND2_X1 U566 ( .A1(n866), .A2(G138), .ZN(n590) );
  INV_X1 U567 ( .A(KEYINPUT17), .ZN(n516) );
  NOR2_X2 U568 ( .A1(n563), .A2(G651), .ZN(n784) );
  NAND2_X1 U569 ( .A1(n617), .A2(n616), .ZN(n931) );
  XNOR2_X2 U570 ( .A(n517), .B(n516), .ZN(n866) );
  NAND2_X1 U571 ( .A1(n866), .A2(G137), .ZN(n526) );
  INV_X1 U572 ( .A(G2105), .ZN(n518) );
  AND2_X1 U573 ( .A1(n518), .A2(G2104), .ZN(n696) );
  NAND2_X1 U574 ( .A1(G101), .A2(n696), .ZN(n519) );
  XNOR2_X1 U575 ( .A(KEYINPUT23), .B(n519), .ZN(n524) );
  INV_X1 U576 ( .A(G2104), .ZN(n586) );
  AND2_X1 U577 ( .A1(n586), .A2(G125), .ZN(n520) );
  NAND2_X1 U578 ( .A1(G2105), .A2(n520), .ZN(n522) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n870) );
  NAND2_X1 U580 ( .A1(G113), .A2(n870), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n524), .A2(n523), .ZN(n525) );
  AND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(G160) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n787) );
  NAND2_X1 U585 ( .A1(G91), .A2(n787), .ZN(n528) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n563) );
  INV_X1 U587 ( .A(G651), .ZN(n532) );
  NOR2_X2 U588 ( .A1(n563), .A2(n532), .ZN(n788) );
  NAND2_X1 U589 ( .A1(G78), .A2(n788), .ZN(n527) );
  NAND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n784), .A2(G53), .ZN(n529) );
  XOR2_X1 U592 ( .A(KEYINPUT68), .B(n529), .Z(n530) );
  NOR2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n536) );
  NOR2_X1 U594 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n533), .Z(n534) );
  NAND2_X1 U596 ( .A1(G65), .A2(n607), .ZN(n535) );
  NAND2_X1 U597 ( .A1(n536), .A2(n535), .ZN(G299) );
  NAND2_X1 U598 ( .A1(n784), .A2(G52), .ZN(n538) );
  NAND2_X1 U599 ( .A1(G64), .A2(n607), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G90), .A2(n787), .ZN(n540) );
  NAND2_X1 U602 ( .A1(G77), .A2(n788), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(KEYINPUT9), .B(n541), .ZN(n542) );
  XNOR2_X1 U605 ( .A(KEYINPUT67), .B(n542), .ZN(n543) );
  NOR2_X1 U606 ( .A1(n544), .A2(n543), .ZN(G171) );
  NAND2_X1 U607 ( .A1(G88), .A2(n787), .ZN(n546) );
  NAND2_X1 U608 ( .A1(G75), .A2(n788), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G62), .A2(n607), .ZN(n547) );
  XNOR2_X1 U611 ( .A(KEYINPUT79), .B(n547), .ZN(n548) );
  NOR2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n784), .A2(G50), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(G303) );
  NAND2_X1 U615 ( .A1(n784), .A2(G51), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G63), .A2(n607), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT6), .B(n554), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n787), .A2(G89), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U621 ( .A1(G76), .A2(n788), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(KEYINPUT5), .B(n558), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT73), .B(n559), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U626 ( .A(KEYINPUT7), .B(n562), .Z(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G87), .A2(n563), .ZN(n570) );
  NAND2_X1 U629 ( .A1(G651), .A2(G74), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G49), .A2(n784), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n607), .A2(n567), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT77), .B(n568), .Z(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT78), .ZN(G288) );
  NAND2_X1 U637 ( .A1(n787), .A2(G86), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G61), .A2(n607), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n788), .A2(G73), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n784), .A2(G48), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(G305) );
  AND2_X1 U645 ( .A1(G60), .A2(n607), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G85), .A2(n787), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G72), .A2(n788), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n784), .A2(G47), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(G290) );
  NAND2_X1 U652 ( .A1(n696), .A2(G102), .ZN(n585) );
  XOR2_X1 U653 ( .A(n585), .B(KEYINPUT82), .Z(n592) );
  AND2_X1 U654 ( .A1(n586), .A2(G2105), .ZN(n869) );
  NAND2_X1 U655 ( .A1(G126), .A2(n869), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G114), .A2(n870), .ZN(n587) );
  AND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U659 ( .A1(n592), .A2(n591), .ZN(G164) );
  AND2_X1 U660 ( .A1(G160), .A2(G40), .ZN(n693) );
  NAND2_X1 U661 ( .A1(n639), .A2(G2072), .ZN(n593) );
  XOR2_X1 U662 ( .A(KEYINPUT27), .B(n593), .Z(n595) );
  NAND2_X1 U663 ( .A1(n648), .A2(G1956), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT91), .ZN(n632) );
  INV_X1 U666 ( .A(G299), .ZN(n798) );
  NOR2_X1 U667 ( .A1(n632), .A2(n798), .ZN(n598) );
  XNOR2_X1 U668 ( .A(n598), .B(n597), .ZN(n636) );
  NAND2_X1 U669 ( .A1(G79), .A2(n788), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n787), .A2(G92), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G66), .A2(n607), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT72), .B(n601), .Z(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X2 U676 ( .A(n606), .B(KEYINPUT15), .ZN(n916) );
  NAND2_X1 U677 ( .A1(G56), .A2(n607), .ZN(n608) );
  XNOR2_X1 U678 ( .A(KEYINPUT14), .B(n608), .ZN(n614) );
  NAND2_X1 U679 ( .A1(G68), .A2(n788), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n787), .A2(G81), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n612), .B(KEYINPUT13), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n615), .B(KEYINPUT69), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n784), .A2(G43), .ZN(n616) );
  INV_X1 U687 ( .A(G1996), .ZN(n1003) );
  NOR2_X1 U688 ( .A1(n648), .A2(n1003), .ZN(n620) );
  XNOR2_X1 U689 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n618), .B(KEYINPUT65), .ZN(n619) );
  XNOR2_X1 U691 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n648), .A2(G1341), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U694 ( .A1(n931), .A2(n623), .ZN(n624) );
  OR2_X1 U695 ( .A1(n916), .A2(n624), .ZN(n631) );
  NAND2_X1 U696 ( .A1(n916), .A2(n624), .ZN(n629) );
  INV_X1 U697 ( .A(G2067), .ZN(n1004) );
  NOR2_X1 U698 ( .A1(n648), .A2(n1004), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT93), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n648), .A2(G1348), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n798), .A2(n632), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U707 ( .A(G2078), .B(KEYINPUT25), .Z(n638) );
  XNOR2_X1 U708 ( .A(KEYINPUT89), .B(n638), .ZN(n995) );
  NAND2_X1 U709 ( .A1(n639), .A2(n995), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n640), .B(KEYINPUT90), .ZN(n642) );
  XOR2_X1 U711 ( .A(G1961), .B(KEYINPUT88), .Z(n952) );
  NAND2_X1 U712 ( .A1(n952), .A2(n648), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n654) );
  NAND2_X1 U714 ( .A1(G171), .A2(n654), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n515), .A2(n643), .ZN(n667) );
  NAND2_X1 U716 ( .A1(G8), .A2(n648), .ZN(n735) );
  NOR2_X1 U717 ( .A1(G1971), .A2(n735), .ZN(n645) );
  NOR2_X1 U718 ( .A1(G2090), .A2(n648), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n646), .A2(G303), .ZN(n660) );
  AND2_X1 U721 ( .A1(n667), .A2(n660), .ZN(n659) );
  NOR2_X1 U722 ( .A1(n735), .A2(G1966), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n647), .B(KEYINPUT87), .ZN(n669) );
  INV_X1 U724 ( .A(G8), .ZN(n649) );
  NOR2_X1 U725 ( .A1(G2084), .A2(n648), .ZN(n668) );
  NOR2_X1 U726 ( .A1(n649), .A2(n668), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n669), .A2(n650), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n651), .B(KEYINPUT30), .ZN(n652) );
  NOR2_X1 U729 ( .A1(G168), .A2(n652), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(KEYINPUT94), .ZN(n656) );
  NOR2_X1 U731 ( .A1(n654), .A2(G171), .ZN(n655) );
  NOR2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n658) );
  INV_X1 U733 ( .A(KEYINPUT31), .ZN(n657) );
  XNOR2_X1 U734 ( .A(n658), .B(n657), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n659), .A2(n666), .ZN(n664) );
  INV_X1 U736 ( .A(n660), .ZN(n661) );
  OR2_X1 U737 ( .A1(n661), .A2(G286), .ZN(n662) );
  AND2_X1 U738 ( .A1(G8), .A2(n662), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(KEYINPUT32), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n673) );
  AND2_X1 U742 ( .A1(G8), .A2(n668), .ZN(n671) );
  INV_X1 U743 ( .A(n669), .ZN(n670) );
  NOR2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  AND2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n674), .B(KEYINPUT95), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n729) );
  NOR2_X1 U748 ( .A1(G288), .A2(G1976), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT96), .ZN(n687) );
  NOR2_X1 U750 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U751 ( .A1(n687), .A2(n678), .ZN(n925) );
  XOR2_X1 U752 ( .A(n925), .B(KEYINPUT97), .Z(n679) );
  NAND2_X1 U753 ( .A1(n729), .A2(n679), .ZN(n680) );
  XNOR2_X1 U754 ( .A(n680), .B(KEYINPUT98), .ZN(n683) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n924) );
  AND2_X1 U756 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U757 ( .A(n684), .B(KEYINPUT64), .ZN(n686) );
  INV_X1 U758 ( .A(n687), .ZN(n688) );
  NOR2_X1 U759 ( .A1(n735), .A2(n688), .ZN(n689) );
  NOR2_X1 U760 ( .A1(n685), .A2(n689), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT99), .ZN(n728) );
  XOR2_X1 U762 ( .A(G1981), .B(G305), .Z(n913) );
  INV_X1 U763 ( .A(n693), .ZN(n694) );
  NOR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n755) );
  NAND2_X1 U765 ( .A1(n697), .A2(G104), .ZN(n698) );
  XOR2_X1 U766 ( .A(KEYINPUT83), .B(n698), .Z(n700) );
  NAND2_X1 U767 ( .A1(n866), .A2(G140), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(KEYINPUT34), .B(n701), .ZN(n706) );
  NAND2_X1 U770 ( .A1(G128), .A2(n869), .ZN(n703) );
  NAND2_X1 U771 ( .A1(G116), .A2(n870), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U773 ( .A(KEYINPUT35), .B(n704), .Z(n705) );
  NOR2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U775 ( .A(KEYINPUT36), .B(n707), .ZN(n888) );
  XNOR2_X1 U776 ( .A(KEYINPUT37), .B(G2067), .ZN(n753) );
  NOR2_X1 U777 ( .A1(n888), .A2(n753), .ZN(n985) );
  NAND2_X1 U778 ( .A1(n755), .A2(n985), .ZN(n751) );
  NAND2_X1 U779 ( .A1(n697), .A2(G105), .ZN(n709) );
  XNOR2_X1 U780 ( .A(KEYINPUT84), .B(KEYINPUT38), .ZN(n708) );
  XNOR2_X1 U781 ( .A(n709), .B(n708), .ZN(n716) );
  NAND2_X1 U782 ( .A1(G129), .A2(n869), .ZN(n711) );
  NAND2_X1 U783 ( .A1(G117), .A2(n870), .ZN(n710) );
  NAND2_X1 U784 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U785 ( .A1(G141), .A2(n866), .ZN(n712) );
  XNOR2_X1 U786 ( .A(KEYINPUT85), .B(n712), .ZN(n713) );
  NOR2_X1 U787 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U788 ( .A1(n716), .A2(n715), .ZN(n855) );
  AND2_X1 U789 ( .A1(n855), .A2(G1996), .ZN(n724) );
  NAND2_X1 U790 ( .A1(G95), .A2(n697), .ZN(n718) );
  NAND2_X1 U791 ( .A1(G131), .A2(n866), .ZN(n717) );
  NAND2_X1 U792 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U793 ( .A1(G119), .A2(n869), .ZN(n720) );
  NAND2_X1 U794 ( .A1(G107), .A2(n870), .ZN(n719) );
  NAND2_X1 U795 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U796 ( .A1(n722), .A2(n721), .ZN(n877) );
  INV_X1 U797 ( .A(G1991), .ZN(n996) );
  NOR2_X1 U798 ( .A1(n877), .A2(n996), .ZN(n723) );
  NOR2_X1 U799 ( .A1(n724), .A2(n723), .ZN(n979) );
  XOR2_X1 U800 ( .A(n755), .B(KEYINPUT86), .Z(n725) );
  NOR2_X1 U801 ( .A1(n979), .A2(n725), .ZN(n747) );
  INV_X1 U802 ( .A(n747), .ZN(n726) );
  AND2_X1 U803 ( .A1(n751), .A2(n726), .ZN(n739) );
  AND2_X1 U804 ( .A1(n913), .A2(n739), .ZN(n727) );
  NAND2_X1 U805 ( .A1(n728), .A2(n727), .ZN(n741) );
  NOR2_X1 U806 ( .A1(G2090), .A2(G303), .ZN(n730) );
  NAND2_X1 U807 ( .A1(G8), .A2(n730), .ZN(n731) );
  NAND2_X1 U808 ( .A1(n729), .A2(n731), .ZN(n732) );
  NAND2_X1 U809 ( .A1(n732), .A2(n735), .ZN(n737) );
  NOR2_X1 U810 ( .A1(G1981), .A2(G305), .ZN(n733) );
  XOR2_X1 U811 ( .A(n733), .B(KEYINPUT24), .Z(n734) );
  OR2_X1 U812 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U813 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U816 ( .A(n742), .B(KEYINPUT100), .ZN(n744) );
  XNOR2_X1 U817 ( .A(G1986), .B(G290), .ZN(n919) );
  NAND2_X1 U818 ( .A1(n919), .A2(n755), .ZN(n743) );
  NAND2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n758) );
  NOR2_X1 U820 ( .A1(G1996), .A2(n855), .ZN(n967) );
  NOR2_X1 U821 ( .A1(G1986), .A2(G290), .ZN(n745) );
  AND2_X1 U822 ( .A1(n996), .A2(n877), .ZN(n976) );
  NOR2_X1 U823 ( .A1(n745), .A2(n976), .ZN(n746) );
  NOR2_X1 U824 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U825 ( .A(KEYINPUT101), .B(n748), .Z(n749) );
  NOR2_X1 U826 ( .A1(n967), .A2(n749), .ZN(n750) );
  XNOR2_X1 U827 ( .A(n750), .B(KEYINPUT39), .ZN(n752) );
  NAND2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U829 ( .A1(n888), .A2(n753), .ZN(n987) );
  NAND2_X1 U830 ( .A1(n754), .A2(n987), .ZN(n756) );
  NAND2_X1 U831 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U832 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U833 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U835 ( .A(G69), .ZN(G235) );
  INV_X1 U836 ( .A(G57), .ZN(G237) );
  NAND2_X1 U837 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U838 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U839 ( .A(G223), .ZN(n823) );
  NAND2_X1 U840 ( .A1(n823), .A2(G567), .ZN(n762) );
  XOR2_X1 U841 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  INV_X1 U842 ( .A(G860), .ZN(n768) );
  OR2_X1 U843 ( .A1(n931), .A2(n768), .ZN(n763) );
  XNOR2_X1 U844 ( .A(KEYINPUT70), .B(n763), .ZN(G153) );
  XNOR2_X1 U845 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U846 ( .A1(G868), .A2(G301), .ZN(n765) );
  OR2_X1 U847 ( .A1(n916), .A2(G868), .ZN(n764) );
  NAND2_X1 U848 ( .A1(n765), .A2(n764), .ZN(G284) );
  INV_X1 U849 ( .A(G868), .ZN(n805) );
  NOR2_X1 U850 ( .A1(G286), .A2(n805), .ZN(n767) );
  NOR2_X1 U851 ( .A1(G868), .A2(G299), .ZN(n766) );
  NOR2_X1 U852 ( .A1(n767), .A2(n766), .ZN(G297) );
  NAND2_X1 U853 ( .A1(n768), .A2(G559), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n769), .A2(n916), .ZN(n770) );
  XNOR2_X1 U855 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U856 ( .A1(G868), .A2(n931), .ZN(n771) );
  XNOR2_X1 U857 ( .A(KEYINPUT74), .B(n771), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G868), .A2(n916), .ZN(n772) );
  NOR2_X1 U859 ( .A1(G559), .A2(n772), .ZN(n773) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(G282) );
  NAND2_X1 U861 ( .A1(G123), .A2(n869), .ZN(n775) );
  XNOR2_X1 U862 ( .A(n775), .B(KEYINPUT18), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n697), .A2(G99), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U865 ( .A1(G135), .A2(n866), .ZN(n779) );
  NAND2_X1 U866 ( .A1(G111), .A2(n870), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n975) );
  XNOR2_X1 U869 ( .A(G2096), .B(n975), .ZN(n783) );
  INV_X1 U870 ( .A(G2100), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(G156) );
  NAND2_X1 U872 ( .A1(n784), .A2(G55), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G67), .A2(n607), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G93), .A2(n787), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G80), .A2(n788), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  OR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n806) );
  NAND2_X1 U879 ( .A1(G559), .A2(n916), .ZN(n793) );
  XNOR2_X1 U880 ( .A(n793), .B(KEYINPUT75), .ZN(n803) );
  XOR2_X1 U881 ( .A(n803), .B(n931), .Z(n794) );
  NOR2_X1 U882 ( .A1(G860), .A2(n794), .ZN(n795) );
  XOR2_X1 U883 ( .A(n806), .B(n795), .Z(G145) );
  XNOR2_X1 U884 ( .A(KEYINPUT19), .B(n806), .ZN(n796) );
  XNOR2_X1 U885 ( .A(G305), .B(n796), .ZN(n797) );
  XNOR2_X1 U886 ( .A(n797), .B(G290), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n798), .B(G288), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n799), .B(G303), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n801), .B(n800), .ZN(n802) );
  XNOR2_X1 U890 ( .A(n802), .B(n931), .ZN(n893) );
  XOR2_X1 U891 ( .A(n893), .B(n803), .Z(n804) );
  NOR2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n808) );
  NOR2_X1 U893 ( .A1(G868), .A2(n806), .ZN(n807) );
  NOR2_X1 U894 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U895 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U897 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U898 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n812), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U901 ( .A1(G237), .A2(G235), .ZN(n813) );
  NAND2_X1 U902 ( .A1(G120), .A2(n813), .ZN(n814) );
  XNOR2_X1 U903 ( .A(KEYINPUT81), .B(n814), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n815), .A2(G108), .ZN(n910) );
  NAND2_X1 U905 ( .A1(n910), .A2(G567), .ZN(n821) );
  NAND2_X1 U906 ( .A1(G132), .A2(G82), .ZN(n816) );
  XNOR2_X1 U907 ( .A(n816), .B(KEYINPUT80), .ZN(n817) );
  XNOR2_X1 U908 ( .A(n817), .B(KEYINPUT22), .ZN(n818) );
  NOR2_X1 U909 ( .A1(G218), .A2(n818), .ZN(n819) );
  NAND2_X1 U910 ( .A1(G96), .A2(n819), .ZN(n911) );
  NAND2_X1 U911 ( .A1(n911), .A2(G2106), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n827) );
  NAND2_X1 U913 ( .A1(G483), .A2(G661), .ZN(n822) );
  NOR2_X1 U914 ( .A1(n827), .A2(n822), .ZN(n826) );
  NAND2_X1 U915 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U918 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(G188) );
  XOR2_X1 U921 ( .A(G120), .B(KEYINPUT102), .Z(G236) );
  XNOR2_X1 U922 ( .A(G96), .B(KEYINPUT103), .ZN(G221) );
  INV_X1 U923 ( .A(n827), .ZN(G319) );
  XOR2_X1 U924 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n829) );
  XNOR2_X1 U925 ( .A(G2678), .B(G2096), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U927 ( .A(n830), .B(KEYINPUT105), .Z(n832) );
  XNOR2_X1 U928 ( .A(G2067), .B(G2072), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U930 ( .A(G2100), .B(G2090), .Z(n834) );
  XNOR2_X1 U931 ( .A(G2078), .B(G2084), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U934 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U936 ( .A(G1981), .B(G1961), .Z(n840) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1966), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U939 ( .A(n841), .B(G2474), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1971), .B(G1976), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(KEYINPUT41), .B(G1956), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G124), .A2(n869), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U948 ( .A1(n697), .A2(G100), .ZN(n849) );
  NAND2_X1 U949 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U950 ( .A1(G136), .A2(n866), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G112), .A2(n870), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U953 ( .A1(n854), .A2(n853), .ZN(G162) );
  XOR2_X1 U954 ( .A(G160), .B(n855), .Z(n887) );
  XNOR2_X1 U955 ( .A(G164), .B(G162), .ZN(n865) );
  NAND2_X1 U956 ( .A1(G130), .A2(n869), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G118), .A2(n870), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U959 ( .A1(n697), .A2(G106), .ZN(n858) );
  XOR2_X1 U960 ( .A(KEYINPUT107), .B(n858), .Z(n860) );
  NAND2_X1 U961 ( .A1(n866), .A2(G142), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT45), .B(n861), .Z(n862) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n880) );
  NAND2_X1 U966 ( .A1(G103), .A2(n697), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G139), .A2(n866), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G127), .A2(n869), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G115), .A2(n870), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(KEYINPUT108), .B(n873), .Z(n874) );
  XNOR2_X1 U973 ( .A(KEYINPUT47), .B(n874), .ZN(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n969) );
  XNOR2_X1 U975 ( .A(n877), .B(n969), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n878), .B(n975), .ZN(n879) );
  XOR2_X1 U977 ( .A(n880), .B(n879), .Z(n885) );
  XOR2_X1 U978 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(KEYINPUT109), .B(n883), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U985 ( .A1(G37), .A2(n890), .ZN(G395) );
  XOR2_X1 U986 ( .A(KEYINPUT112), .B(G286), .Z(n892) );
  XNOR2_X1 U987 ( .A(G171), .B(n916), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2451), .B(G2430), .Z(n897) );
  XNOR2_X1 U992 ( .A(G2438), .B(G2443), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n903) );
  XOR2_X1 U994 ( .A(G2435), .B(G2454), .Z(n899) );
  XNOR2_X1 U995 ( .A(G1348), .B(G1341), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U997 ( .A(G2446), .B(G2427), .Z(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U999 ( .A(n903), .B(n902), .Z(n904) );
  NAND2_X1 U1000 ( .A1(G14), .A2(n904), .ZN(n912) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n912), .ZN(n907) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(G225) );
  XNOR2_X1 U1007 ( .A(KEYINPUT113), .B(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G132), .ZN(G219) );
  INV_X1 U1010 ( .A(G108), .ZN(G238) );
  INV_X1 U1011 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(G325) );
  INV_X1 U1013 ( .A(G325), .ZN(G261) );
  INV_X1 U1014 ( .A(G303), .ZN(G166) );
  INV_X1 U1015 ( .A(n912), .ZN(G401) );
  XNOR2_X1 U1016 ( .A(G16), .B(KEYINPUT56), .ZN(n937) );
  XNOR2_X1 U1017 ( .A(G1966), .B(G168), .ZN(n914) );
  NAND2_X1 U1018 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1019 ( .A(n915), .B(KEYINPUT57), .ZN(n935) );
  XNOR2_X1 U1020 ( .A(n916), .B(G1348), .ZN(n917) );
  XNOR2_X1 U1021 ( .A(n917), .B(KEYINPUT122), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G1956), .B(G299), .ZN(n918) );
  NOR2_X1 U1023 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n923) );
  XOR2_X1 U1025 ( .A(G171), .B(G1961), .Z(n922) );
  NOR2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n927) );
  AND2_X1 U1028 ( .A1(G303), .A2(G1971), .ZN(n926) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1030 ( .A(KEYINPUT123), .B(n928), .Z(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(G1341), .B(n931), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n965) );
  INV_X1 U1036 ( .A(G16), .ZN(n963) );
  XOR2_X1 U1037 ( .A(G1986), .B(G24), .Z(n940) );
  XNOR2_X1 U1038 ( .A(G23), .B(KEYINPUT125), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n938), .B(G1976), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G22), .B(G1971), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1043 ( .A(KEYINPUT58), .B(n943), .Z(n959) );
  XNOR2_X1 U1044 ( .A(G1348), .B(KEYINPUT59), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(n944), .B(G4), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(G1981), .B(G6), .ZN(n945) );
  NOR2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(G20), .B(G1956), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(KEYINPUT60), .B(n951), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(n952), .B(G5), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(G21), .B(G1966), .ZN(n955) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1057 ( .A(KEYINPUT124), .B(n957), .Z(n958) );
  NOR2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1059 ( .A(n960), .B(KEYINPUT61), .ZN(n961) );
  XNOR2_X1 U1060 ( .A(n961), .B(KEYINPUT126), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n994) );
  XOR2_X1 U1063 ( .A(G2090), .B(G162), .Z(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT51), .B(n968), .ZN(n974) );
  XOR2_X1 U1066 ( .A(G2072), .B(n969), .Z(n971) );
  XOR2_X1 U1067 ( .A(G164), .B(G2078), .Z(n970) );
  NOR2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1069 ( .A(KEYINPUT50), .B(n972), .Z(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n983) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n977), .B(KEYINPUT114), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n981) );
  XOR2_X1 U1074 ( .A(G160), .B(G2084), .Z(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n988), .B(KEYINPUT115), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(KEYINPUT52), .B(n989), .ZN(n990) );
  XOR2_X1 U1081 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n1017) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n1017), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(G29), .A2(n991), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(KEYINPUT117), .B(n992), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1024) );
  INV_X1 U1086 ( .A(G29), .ZN(n1020) );
  XOR2_X1 U1087 ( .A(G2090), .B(G35), .Z(n1012) );
  XNOR2_X1 U1088 ( .A(G27), .B(n995), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G25), .B(n996), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n997), .A2(G28), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(KEYINPUT118), .B(G2072), .ZN(n998) );
  XNOR2_X1 U1092 ( .A(G33), .B(n998), .ZN(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(n1003), .B(G32), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1004), .B(G26), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(KEYINPUT119), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT53), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G34), .B(G2084), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT54), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(KEYINPUT120), .ZN(n1018) );
  XOR2_X1 U1106 ( .A(n1018), .B(n1017), .Z(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(G11), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(n1022), .B(KEYINPUT121), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

