//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT65), .B(G68), .ZN(new_n208));
  AND2_X1   g0008(.A1(new_n208), .A2(G238), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G58), .A2(G232), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n207), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT66), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n207), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(G58), .A2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n201), .B1(new_n227), .B2(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n228), .B1(KEYINPUT64), .B2(new_n227), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n222), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  AND3_X1   g0031(.A1(new_n218), .A2(new_n219), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n251), .A2(G77), .B1(new_n252), .B2(G50), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(new_n224), .B2(new_n208), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(new_n223), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n255), .A3(new_n223), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT11), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n254), .A2(KEYINPUT11), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT76), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(KEYINPUT76), .A3(new_n264), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G13), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n224), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n256), .A2(new_n223), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n224), .A2(G1), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n274), .A2(new_n203), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G13), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT12), .B1(new_n279), .B2(new_n208), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n280), .B(KEYINPUT77), .ZN(new_n281));
  OR3_X1    g0081(.A1(new_n279), .A2(KEYINPUT12), .A3(G68), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n267), .A2(new_n268), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n287), .A2(new_n289), .A3(G232), .A4(G1698), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n287), .A2(new_n289), .A3(G226), .A4(new_n291), .ZN(new_n292));
  AND3_X1   g0092(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT75), .B1(G33), .B2(G97), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n290), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(G1), .A3(G13), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT13), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  AOI21_X1  g0105(.A(G1), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G274), .ZN(new_n307));
  INV_X1    g0107(.A(new_n223), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n297), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n303), .A2(G238), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n300), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n301), .B1(new_n300), .B2(new_n310), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n286), .B(G169), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT78), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n300), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n300), .A2(new_n301), .A3(new_n310), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n319), .A2(KEYINPUT78), .A3(new_n286), .A4(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(G169), .B1(new_n311), .B2(new_n312), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n311), .A2(new_n312), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n322), .A2(KEYINPUT14), .B1(new_n323), .B2(G179), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n285), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n319), .A2(new_n328), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n327), .A2(new_n284), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n288), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n333));
  OAI21_X1  g0133(.A(G77), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n287), .A2(new_n289), .A3(G222), .A4(new_n291), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n287), .A2(new_n289), .A3(G223), .A4(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n299), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n306), .A2(new_n298), .A3(G274), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n298), .A2(G226), .A3(new_n302), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(G179), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT69), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n275), .A2(new_n201), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n258), .A2(new_n346), .A3(new_n279), .A4(new_n259), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n279), .A2(G50), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n224), .A2(G33), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT8), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G58), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n224), .B1(new_n226), .B2(new_n201), .ZN(new_n355));
  INV_X1    g0155(.A(G150), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n356), .A2(G20), .A3(G33), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n259), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n257), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n347), .B(new_n349), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(new_n343), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n345), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n351), .A2(new_n353), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n350), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n272), .ZN(new_n370));
  INV_X1    g0170(.A(G77), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n275), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n273), .A2(new_n372), .B1(new_n371), .B2(new_n271), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n303), .A2(G244), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n339), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT3), .B(G33), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(G232), .A3(new_n291), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(G238), .A3(G1698), .ZN(new_n379));
  INV_X1    g0179(.A(G107), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT70), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT70), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G107), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n378), .B(new_n379), .C1(new_n377), .C2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n376), .B1(new_n299), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n374), .B1(new_n386), .B2(G190), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n326), .B2(new_n386), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n374), .B1(new_n386), .B2(G169), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n365), .A2(new_n388), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT10), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n361), .A2(new_n396), .A3(KEYINPUT9), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n204), .A2(G20), .ZN(new_n398));
  INV_X1    g0198(.A(new_n357), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT8), .B(G58), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n398), .B(new_n399), .C1(new_n400), .C2(new_n350), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n348), .B1(new_n401), .B2(new_n260), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n396), .A2(KEYINPUT9), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n396), .A2(KEYINPUT9), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n402), .A2(new_n347), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n328), .B(new_n341), .C1(new_n299), .C2(new_n337), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n326), .B1(new_n338), .B2(new_n342), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n395), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n411));
  XOR2_X1   g0211(.A(KEYINPUT73), .B(KEYINPUT10), .Z(new_n412));
  NOR3_X1   g0212(.A1(new_n407), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n397), .A2(new_n414), .A3(new_n405), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n397), .B2(new_n405), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n410), .A2(KEYINPUT74), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n331), .B(new_n394), .C1(new_n411), .C2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(new_n208), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n377), .B2(G20), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n287), .A2(new_n289), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n252), .A2(G159), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n226), .B1(new_n208), .B2(G58), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(new_n224), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n420), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT7), .B1(new_n424), .B2(new_n224), .ZN(new_n431));
  AOI211_X1 g0231(.A(new_n422), .B(G20), .C1(new_n287), .C2(new_n289), .ZN(new_n432));
  OAI21_X1  g0232(.A(G68), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(KEYINPUT65), .A2(G68), .ZN(new_n434));
  NOR2_X1   g0234(.A1(KEYINPUT65), .A2(G68), .ZN(new_n435));
  OAI21_X1  g0235(.A(G58), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n227), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(G20), .B1(G159), .B2(new_n252), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n433), .A2(KEYINPUT16), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n430), .A2(new_n439), .A3(new_n272), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n260), .A2(new_n271), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n400), .A2(new_n275), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n441), .A2(new_n442), .B1(new_n271), .B2(new_n400), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n287), .A2(new_n289), .A3(G226), .A4(G1698), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n287), .A2(new_n289), .A3(G223), .A4(new_n291), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G87), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n299), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n303), .A2(G232), .B1(new_n306), .B2(new_n309), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT80), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n451), .A2(new_n455), .A3(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n457), .A2(new_n363), .B1(new_n389), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n440), .A2(KEYINPUT79), .A3(new_n443), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n446), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(G200), .B1(new_n454), .B2(new_n456), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n453), .A2(G190), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n443), .B(new_n440), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n443), .ZN(new_n470));
  INV_X1    g0270(.A(new_n272), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n203), .B1(new_n423), .B2(new_n425), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n429), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n473), .B2(KEYINPUT16), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n470), .B1(new_n474), .B2(new_n430), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n451), .A2(new_n455), .A3(new_n452), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n455), .B1(new_n451), .B2(new_n452), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n326), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n466), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n475), .A2(new_n480), .A3(KEYINPUT17), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n463), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n446), .A2(new_n459), .A3(new_n460), .A4(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n464), .A2(new_n469), .A3(new_n481), .A4(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n419), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n305), .A2(G1), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n309), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(G270), .A3(new_n298), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n287), .A2(new_n289), .A3(G264), .A4(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n287), .A2(new_n289), .A3(G257), .A4(new_n291), .ZN(new_n496));
  INV_X1    g0296(.A(G303), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n377), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n299), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n269), .A2(G33), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G116), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n224), .A2(G116), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n273), .A2(new_n503), .B1(new_n278), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n223), .B2(new_n256), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n507), .B(new_n224), .C1(G33), .C2(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n506), .A2(KEYINPUT20), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT20), .B1(new_n506), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n500), .A2(new_n512), .A3(G169), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n500), .A2(G200), .ZN(new_n516));
  INV_X1    g0316(.A(new_n512), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n494), .A2(new_n499), .A3(G190), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n500), .A2(new_n389), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n512), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n500), .A2(new_n512), .A3(KEYINPUT21), .A4(G169), .ZN(new_n522));
  AND4_X1   g0322(.A1(new_n515), .A2(new_n519), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n287), .A2(new_n289), .A3(new_n224), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n377), .A2(new_n526), .A3(new_n224), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT23), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n380), .A3(G20), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n350), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n381), .A2(new_n383), .A3(G20), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(KEYINPUT23), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n528), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n471), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n258), .A2(new_n279), .A3(new_n259), .A4(new_n501), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n380), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n278), .A2(G20), .A3(new_n380), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT25), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT87), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n538), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n537), .B1(new_n528), .B2(new_n534), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n272), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT87), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n544), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n287), .A2(new_n289), .A3(G257), .A4(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n287), .A2(new_n289), .A3(G250), .A4(new_n291), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G294), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n487), .A2(new_n488), .B1(new_n308), .B2(new_n297), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n555), .A2(new_n299), .B1(new_n556), .B2(G264), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n489), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G169), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n389), .B2(new_n558), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n546), .A2(new_n551), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n309), .A2(new_n488), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n298), .B(G250), .C1(G1), .C2(new_n305), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n287), .A2(new_n289), .A3(G244), .A4(G1698), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G116), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n377), .A2(new_n569), .A3(G238), .A4(new_n291), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n287), .A2(new_n289), .A3(G238), .A4(new_n291), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT84), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n565), .B1(new_n573), .B2(new_n298), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G190), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(G200), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n271), .A2(new_n368), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT19), .B1(new_n293), .B2(new_n294), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n224), .ZN(new_n581));
  NOR2_X1   g0381(.A1(G87), .A2(G97), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n384), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n377), .A2(KEYINPUT85), .A3(new_n224), .A4(G68), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n287), .A2(new_n289), .A3(new_n224), .A4(G68), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT85), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n251), .A2(G97), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n586), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n584), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n579), .B1(new_n591), .B2(new_n272), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n441), .A2(G87), .A3(new_n501), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n576), .A2(new_n577), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n572), .A2(new_n570), .ZN(new_n595));
  INV_X1    g0395(.A(new_n568), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n298), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n363), .B1(new_n597), .B2(new_n564), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n389), .B(new_n565), .C1(new_n573), .C2(new_n298), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT86), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n590), .A2(new_n585), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n224), .A2(new_n580), .B1(new_n384), .B2(new_n582), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n272), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n540), .A2(new_n368), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n601), .A2(new_n604), .A3(new_n578), .A4(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n601), .B1(new_n592), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n523), .A2(new_n561), .A3(new_n594), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n492), .A2(G257), .A3(new_n298), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT82), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n287), .A2(new_n289), .A3(G244), .A4(new_n291), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT4), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n377), .A2(KEYINPUT4), .A3(G244), .A4(new_n291), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n377), .A2(G250), .A3(G1698), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n507), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n299), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n611), .A2(new_n618), .A3(new_n489), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT83), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n611), .A2(new_n618), .A3(KEYINPUT83), .A4(new_n489), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(G200), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n271), .A2(new_n508), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n540), .B2(new_n508), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT6), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n508), .A2(new_n380), .ZN(new_n627));
  NOR2_X1   g0427(.A1(G97), .A2(G107), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n380), .A2(KEYINPUT6), .A3(G97), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(G20), .B1(G77), .B2(new_n252), .ZN(new_n632));
  INV_X1    g0432(.A(new_n384), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n431), .B2(new_n432), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n625), .B1(new_n635), .B2(new_n272), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n611), .A2(new_n618), .A3(G190), .A4(new_n489), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n623), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n636), .B1(new_n363), .B2(new_n619), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n611), .A2(new_n618), .A3(new_n389), .A4(new_n489), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n558), .A2(G200), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n557), .A2(G190), .A3(new_n489), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n549), .A2(new_n643), .A3(new_n544), .A4(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n639), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n609), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n486), .A2(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n469), .A2(new_n481), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n330), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n325), .B2(new_n392), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n363), .B1(new_n476), .B2(new_n477), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n458), .A2(new_n389), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n444), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT18), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT18), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n459), .A2(new_n656), .A3(new_n444), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n651), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT90), .B1(new_n418), .B2(new_n411), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT74), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n406), .A2(new_n409), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n395), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT90), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n666));
  INV_X1    g0466(.A(new_n417), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n415), .A3(new_n413), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n664), .A2(new_n665), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n660), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n365), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n608), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT88), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n595), .A2(new_n596), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n299), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n326), .B1(new_n678), .B2(new_n565), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n604), .A2(new_n593), .A3(new_n578), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n577), .A2(new_n592), .A3(KEYINPUT88), .A4(new_n593), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n576), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n608), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n646), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n515), .A2(new_n521), .A3(new_n522), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n560), .B1(new_n539), .B2(new_n545), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n675), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n619), .A2(new_n363), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n635), .A2(new_n272), .ZN(new_n691));
  INV_X1    g0491(.A(new_n625), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n690), .A2(new_n693), .A3(new_n641), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n683), .A2(new_n694), .A3(new_n608), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT26), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n608), .A2(new_n694), .A3(KEYINPUT26), .A4(new_n594), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT89), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n604), .A2(new_n578), .A3(new_n605), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT86), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n592), .A2(new_n601), .A3(new_n605), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n679), .A2(new_n680), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n704), .A2(new_n600), .B1(new_n705), .B2(new_n576), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n694), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n697), .A2(new_n700), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n689), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n486), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n674), .A2(new_n710), .ZN(G369));
  INV_X1    g0511(.A(new_n686), .ZN(new_n712));
  OR3_X1    g0512(.A1(new_n270), .A2(KEYINPUT27), .A3(G20), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT27), .B1(new_n270), .B2(G20), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G213), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G343), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n517), .A2(new_n718), .ZN(new_n719));
  MUX2_X1   g0519(.A(new_n523), .B(new_n712), .S(new_n719), .Z(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n546), .A2(new_n551), .A3(new_n560), .A4(new_n717), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n546), .A2(new_n551), .A3(new_n717), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n561), .A2(new_n727), .A3(new_n645), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n712), .A2(new_n718), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n726), .B2(new_n728), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n687), .A2(new_n717), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(G399));
  NOR2_X1   g0535(.A1(new_n583), .A2(G116), .ZN(new_n736));
  INV_X1    g0536(.A(new_n220), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G41), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(G1), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n741), .A2(KEYINPUT92), .B1(new_n230), .B2(new_n738), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(KEYINPUT92), .B2(new_n741), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT94), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n717), .B1(new_n689), .B2(new_n708), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(KEYINPUT29), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n697), .A2(new_n700), .A3(new_n707), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n577), .A2(new_n592), .A3(new_n593), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n749), .A2(new_n676), .B1(G190), .B2(new_n575), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n750), .A2(new_n682), .B1(new_n704), .B2(new_n600), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n694), .B1(new_n623), .B2(new_n638), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n751), .A2(new_n752), .A3(new_n645), .A4(new_n688), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n608), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n718), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(KEYINPUT94), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n639), .A2(new_n642), .A3(new_n645), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n561), .A2(KEYINPUT95), .A3(new_n686), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT95), .B1(new_n561), .B2(new_n686), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n759), .B(new_n751), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT96), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n685), .B(KEYINPUT96), .C1(new_n761), .C2(new_n760), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n695), .A2(KEYINPUT26), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n706), .A2(new_n696), .A3(new_n694), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n766), .A2(new_n608), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n764), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT29), .A3(new_n718), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n523), .A2(new_n561), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n759), .A2(new_n771), .A3(new_n706), .A4(new_n718), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n557), .B(new_n565), .C1(new_n573), .C2(new_n298), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT93), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n611), .A2(new_n618), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n678), .A2(KEYINPUT93), .A3(new_n557), .A4(new_n565), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n775), .A2(new_n777), .A3(new_n778), .A4(new_n520), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT30), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n776), .A2(new_n389), .A3(new_n500), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n782), .A2(KEYINPUT30), .A3(new_n778), .A4(new_n775), .ZN(new_n783));
  AOI21_X1  g0583(.A(G179), .B1(new_n494), .B2(new_n499), .ZN(new_n784));
  AND4_X1   g0584(.A1(new_n619), .A2(new_n558), .A3(new_n574), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n781), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n717), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT31), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n785), .B1(new_n779), .B2(new_n780), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n718), .B1(new_n791), .B2(new_n783), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT31), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n772), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n758), .A2(new_n770), .B1(G330), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n744), .B1(new_n795), .B2(G1), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT97), .Z(G364));
  NOR2_X1   g0597(.A1(new_n277), .A2(G20), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n269), .B1(new_n798), .B2(G45), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n739), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n723), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G330), .B2(new_n720), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n377), .A2(new_n220), .ZN(new_n804));
  INV_X1    g0604(.A(G355), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n805), .B1(G116), .B2(new_n220), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n245), .A2(new_n305), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT98), .Z(new_n808));
  NOR2_X1   g0608(.A1(new_n737), .A2(new_n377), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n230), .B2(new_n305), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n806), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G13), .A2(G33), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n223), .B1(G20), .B2(new_n363), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n801), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n389), .A2(G200), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(G20), .A3(G190), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n224), .A2(G190), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n822), .A2(G58), .B1(new_n825), .B2(G77), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n328), .A2(new_n326), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n224), .A2(G179), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G87), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n377), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n827), .A2(KEYINPUT99), .B1(new_n833), .B2(KEYINPUT100), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n326), .A2(G190), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n380), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n224), .A2(new_n389), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n837), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n839), .B1(G68), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n828), .A2(new_n840), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n201), .B2(new_n844), .C1(new_n827), .C2(KEYINPUT99), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT32), .ZN(new_n846));
  NOR2_X1   g0646(.A1(G179), .A2(G200), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n823), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n849), .B2(G159), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n846), .A3(G159), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n224), .B1(new_n847), .B2(G190), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(G97), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  OR4_X1    g0655(.A1(new_n836), .A2(new_n845), .A3(new_n850), .A4(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(KEYINPUT101), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G303), .A2(new_n831), .B1(new_n825), .B2(G311), .ZN(new_n858));
  INV_X1    g0658(.A(G326), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(new_n424), .C1(new_n859), .C2(new_n844), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n822), .A2(G322), .B1(new_n849), .B2(G329), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  XOR2_X1   g0662(.A(KEYINPUT33), .B(G317), .Z(new_n863));
  OAI221_X1 g0663(.A(new_n861), .B1(new_n862), .B2(new_n838), .C1(new_n841), .C2(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n860), .B(new_n864), .C1(G294), .C2(new_n853), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n856), .B2(KEYINPUT101), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n857), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n819), .B1(new_n867), .B2(new_n816), .ZN(new_n868));
  INV_X1    g0668(.A(new_n815), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n720), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n803), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(G396));
  NAND3_X1  g0672(.A1(new_n393), .A2(new_n388), .A3(new_n718), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n748), .B2(new_n754), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n393), .A2(new_n717), .ZN(new_n876));
  INV_X1    g0676(.A(new_n374), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n388), .B1(new_n877), .B2(new_n718), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n393), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n875), .B1(new_n746), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n794), .A2(G330), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n801), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n816), .A2(new_n813), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n801), .B1(G77), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT102), .ZN(new_n887));
  INV_X1    g0687(.A(new_n816), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n841), .A2(new_n356), .ZN(new_n889));
  INV_X1    g0689(.A(G143), .ZN(new_n890));
  INV_X1    g0690(.A(G159), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n821), .A2(new_n890), .B1(new_n824), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n844), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n889), .B(new_n892), .C1(G137), .C2(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(KEYINPUT34), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n377), .B1(new_n838), .B2(new_n203), .ZN(new_n896));
  INV_X1    g0696(.A(G132), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n830), .A2(new_n201), .B1(new_n848), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n896), .B(new_n898), .C1(G58), .C2(new_n853), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n894), .A2(KEYINPUT34), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n895), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n838), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(G87), .ZN(new_n903));
  INV_X1    g0703(.A(G311), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n848), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n377), .B(new_n905), .C1(G303), .C2(new_n893), .ZN(new_n906));
  AOI22_X1  g0706(.A1(G294), .A2(new_n822), .B1(new_n842), .B2(G283), .ZN(new_n907));
  AOI22_X1  g0707(.A1(G107), .A2(new_n831), .B1(new_n825), .B2(G116), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n906), .A2(new_n854), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n887), .B1(new_n888), .B2(new_n910), .C1(new_n879), .C2(new_n814), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n883), .A2(new_n911), .ZN(G384));
  NOR2_X1   g0712(.A1(new_n798), .A2(new_n269), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n440), .A2(KEYINPUT79), .A3(new_n443), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT79), .B1(new_n440), .B2(new_n443), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n914), .A2(new_n915), .A3(new_n715), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n467), .A2(new_n654), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n715), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n446), .A2(new_n460), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT37), .B1(new_n475), .B2(new_n480), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n461), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n916), .B1(new_n649), .B2(new_n658), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n420), .B1(new_n472), .B2(new_n429), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n439), .A3(new_n260), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n443), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n919), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n652), .A3(new_n653), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n467), .A2(new_n931), .A3(new_n929), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT37), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n485), .A2(new_n930), .B1(new_n933), .B2(new_n922), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n925), .B1(KEYINPUT38), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n876), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n878), .A2(new_n393), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n284), .A2(new_n717), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n331), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n939), .B1(new_n321), .B2(new_n324), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n938), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT105), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n789), .B1(new_n792), .B2(new_n944), .ZN(new_n945));
  AOI211_X1 g0745(.A(KEYINPUT105), .B(new_n718), .C1(new_n791), .C2(new_n783), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n772), .A2(new_n793), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT40), .B1(new_n935), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n652), .A2(new_n653), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n914), .A2(new_n915), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n484), .B1(new_n952), .B2(new_n462), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n930), .B1(new_n953), .B2(new_n649), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n933), .A2(new_n922), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT38), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n934), .A2(KEYINPUT38), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT40), .ZN(new_n961));
  INV_X1    g0761(.A(new_n939), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n325), .A2(new_n330), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n879), .B1(new_n963), .B2(new_n941), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n788), .A2(KEYINPUT105), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n792), .A2(new_n944), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n966), .A3(new_n789), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n647), .A2(new_n718), .B1(KEYINPUT31), .B2(new_n792), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n960), .A2(new_n961), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n950), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT106), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n967), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(new_n486), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n722), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n972), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT39), .ZN(new_n977));
  AOI221_X4 g0777(.A(new_n957), .B1(new_n933), .B2(new_n922), .C1(new_n485), .C2(new_n930), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n978), .B2(new_n925), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT39), .ZN(new_n980));
  INV_X1    g0780(.A(new_n325), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n717), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n875), .A2(new_n936), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n963), .A2(new_n941), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n960), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n659), .A2(new_n919), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n983), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT104), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT104), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n983), .A2(new_n987), .A3(new_n992), .A4(new_n989), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n486), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n766), .A2(new_n608), .A3(new_n767), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n763), .B2(new_n762), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n717), .B1(new_n997), .B2(new_n765), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n995), .B1(new_n998), .B2(KEYINPUT29), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n673), .B1(new_n999), .B2(new_n758), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n994), .B(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n913), .B1(new_n976), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n976), .B2(new_n1001), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n631), .B(KEYINPUT103), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT35), .ZN(new_n1005));
  OAI211_X1 g0805(.A(G116), .B(new_n225), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n1005), .B2(new_n1004), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT36), .Z(new_n1008));
  NAND3_X1  g0808(.A1(new_n230), .A2(G77), .A3(new_n436), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(G50), .B2(new_n203), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(G1), .A3(new_n277), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1003), .A2(new_n1008), .A3(new_n1011), .ZN(G367));
  INV_X1    g0812(.A(KEYINPUT108), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n680), .A2(new_n717), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n608), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n751), .B2(new_n1014), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT42), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n732), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n639), .B(new_n642), .C1(new_n636), .C2(new_n718), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n694), .A2(new_n717), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1018), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n732), .A2(KEYINPUT42), .A3(new_n1022), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n642), .B1(new_n1020), .B2(new_n561), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(KEYINPUT107), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n718), .B1(new_n1027), .B2(KEYINPUT107), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1013), .B(new_n1017), .C1(new_n1026), .C2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1030), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1016), .B1(new_n1032), .B2(KEYINPUT108), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT43), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n730), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1031), .A2(new_n1033), .A3(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1022), .A4(new_n1039), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1031), .A2(new_n1033), .A3(new_n1038), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT43), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1041), .A2(new_n1042), .B1(new_n730), .B2(new_n1023), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n738), .B(KEYINPUT41), .Z(new_n1044));
  INV_X1    g0844(.A(new_n734), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT44), .B1(new_n1045), .B2(new_n1023), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT44), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n734), .A2(new_n1047), .A3(new_n1022), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT45), .B1(new_n734), .B2(new_n1022), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT45), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n732), .A2(new_n1050), .A3(new_n1023), .A4(new_n733), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1046), .A2(new_n1048), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n1037), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n730), .B1(new_n1049), .B2(new_n1051), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n729), .B(new_n731), .Z(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(new_n723), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n795), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1044), .B1(new_n1057), .B2(new_n795), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n799), .B(KEYINPUT109), .Z(new_n1059));
  OAI211_X1 g0859(.A(new_n1040), .B(new_n1043), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n237), .A2(new_n810), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n817), .B1(new_n220), .B2(new_n368), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n801), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n844), .A2(new_n890), .B1(new_n838), .B2(new_n371), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n424), .B(new_n1064), .C1(G150), .C2(new_n822), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G159), .A2(new_n842), .B1(new_n849), .B2(G137), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G58), .A2(new_n831), .B1(new_n825), .B2(G50), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n852), .A2(new_n203), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n830), .A2(new_n531), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(KEYINPUT46), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1072), .A2(KEYINPUT112), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n838), .A2(new_n508), .ZN(new_n1074));
  INV_X1    g0874(.A(G294), .ZN(new_n1075));
  INV_X1    g0875(.A(G317), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n841), .A2(new_n1075), .B1(new_n848), .B2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(KEYINPUT112), .B2(new_n1072), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(KEYINPUT110), .B(G311), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n844), .A2(new_n1080), .B1(new_n821), .B2(new_n497), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT111), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n424), .B1(new_n824), .B2(new_n862), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n633), .B2(new_n853), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(KEYINPUT46), .C2(new_n1071), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1070), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT47), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1063), .B1(new_n1087), .B2(new_n816), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1017), .B2(new_n869), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1060), .A2(new_n1089), .ZN(G387));
  NAND2_X1  g0890(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n809), .B1(new_n241), .B2(new_n305), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n736), .B2(new_n804), .ZN(new_n1093));
  OR3_X1    g0893(.A1(new_n400), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1094));
  AOI21_X1  g0894(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT50), .B1(new_n400), .B2(G50), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n736), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1093), .A2(new_n1097), .B1(new_n380), .B2(new_n737), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n801), .B1(new_n1098), .B2(new_n818), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n822), .A2(G317), .B1(new_n825), .B2(G303), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n893), .A2(G322), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n841), .C2(new_n1080), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT48), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n830), .A2(new_n1075), .B1(new_n852), .B2(new_n862), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(KEYINPUT49), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n377), .B1(new_n902), .B2(G116), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n859), .C2(new_n848), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT49), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n841), .A2(new_n400), .B1(new_n824), .B2(new_n203), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT113), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n893), .A2(G159), .B1(new_n849), .B2(G150), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n201), .B2(new_n821), .C1(new_n371), .C2(new_n830), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n852), .A2(new_n368), .ZN(new_n1115));
  OR4_X1    g0915(.A1(new_n424), .A2(new_n1114), .A3(new_n1074), .A4(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1109), .A2(new_n1110), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1117), .A2(KEYINPUT114), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n888), .B1(new_n1117), .B2(KEYINPUT114), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1099), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n729), .B2(new_n869), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n795), .A2(new_n1056), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n738), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n795), .A2(new_n1056), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1091), .B(new_n1121), .C1(new_n1123), .C2(new_n1124), .ZN(G393));
  NAND3_X1  g0925(.A1(new_n1053), .A2(new_n1054), .A3(new_n1059), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n844), .A2(new_n1076), .B1(new_n821), .B2(new_n904), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT52), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G283), .A2(new_n831), .B1(new_n842), .B2(G303), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n825), .A2(G294), .B1(new_n849), .B2(G322), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n377), .B(new_n839), .C1(G116), .C2(new_n853), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n853), .A2(G77), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n201), .B2(new_n841), .C1(new_n400), .C2(new_n824), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT115), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n844), .A2(new_n356), .B1(new_n821), .B2(new_n891), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT51), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n208), .A2(new_n831), .B1(new_n849), .B2(G143), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1137), .A2(new_n377), .A3(new_n903), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1132), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n816), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n818), .B1(G97), .B2(new_n737), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n248), .A2(new_n809), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n800), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1141), .B(new_n1144), .C1(new_n1022), .C2(new_n869), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1146), .A2(new_n1122), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1057), .A2(new_n738), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1126), .B(new_n1145), .C1(new_n1147), .C2(new_n1148), .ZN(G390));
  NAND3_X1  g0949(.A1(new_n973), .A2(G330), .A3(new_n943), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n982), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n978), .B2(new_n925), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n769), .A2(new_n718), .A3(new_n937), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n936), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n1155), .B2(new_n986), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n873), .B1(new_n689), .B2(new_n708), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n986), .B1(new_n1157), .B2(new_n876), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n979), .A2(new_n980), .B1(new_n1158), .B2(new_n1152), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1151), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1152), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n979), .A2(new_n980), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n986), .A2(new_n794), .A3(G330), .A4(new_n879), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n985), .B1(new_n1154), .B2(new_n936), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1163), .B(new_n1164), .C1(new_n1165), .C2(new_n1153), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n722), .B1(new_n968), .B2(new_n967), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1167), .A2(new_n486), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n673), .B(new_n1168), .C1(new_n999), .C2(new_n758), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n985), .B1(new_n881), .B2(new_n938), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1170), .A2(new_n1150), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1157), .A2(new_n876), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1154), .A2(new_n936), .A3(new_n1164), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n986), .B1(new_n1167), .B2(new_n879), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1171), .A2(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1160), .A2(new_n1166), .A3(new_n1169), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT116), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(new_n1177), .A3(new_n738), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1176), .A2(new_n738), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT116), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1160), .A2(new_n1166), .A3(new_n1059), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1162), .A2(new_n813), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n801), .B1(new_n366), .B2(new_n885), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n821), .A2(new_n897), .B1(new_n838), .B2(new_n201), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G128), .B2(new_n893), .ZN(new_n1189));
  INV_X1    g0989(.A(G137), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT54), .B(G143), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n841), .A2(new_n1190), .B1(new_n824), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT117), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1189), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n830), .A2(KEYINPUT53), .A3(new_n356), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n424), .B1(new_n849), .B2(G125), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT53), .B1(new_n830), .B2(new_n356), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n853), .A2(G159), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n822), .A2(G116), .B1(new_n825), .B2(G97), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n862), .B2(new_n844), .C1(new_n384), .C2(new_n841), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n902), .A2(G68), .B1(new_n849), .B2(G294), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1204), .A2(new_n424), .A3(new_n832), .A4(new_n1133), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1196), .A2(new_n1201), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1187), .B1(new_n1206), .B2(new_n816), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1186), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1185), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT118), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1185), .A2(KEYINPUT118), .A3(new_n1208), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1182), .A2(new_n1184), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(G378));
  NAND2_X1  g1014(.A1(new_n971), .A2(G330), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n661), .A2(new_n365), .A3(new_n669), .ZN(new_n1216));
  XOR2_X1   g1016(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n661), .A2(new_n669), .A3(new_n365), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n362), .A2(new_n715), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1222), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1218), .A2(new_n1225), .A3(new_n1220), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1224), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1218), .A2(new_n1225), .A3(new_n1220), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1215), .A2(new_n1227), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1227), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n971), .A2(new_n1233), .A3(G330), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n994), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n971), .A2(new_n1233), .A3(G330), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(G330), .B2(new_n971), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n993), .B(new_n991), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1235), .A2(new_n1238), .B1(new_n1176), .B2(new_n1169), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n739), .B1(new_n1239), .B2(KEYINPUT57), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1176), .A2(new_n1169), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT57), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1231), .A2(new_n1227), .A3(new_n813), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n893), .A2(G125), .B1(new_n853), .B2(G150), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT119), .Z(new_n1249));
  NOR2_X1   g1049(.A1(new_n824), .A2(new_n1190), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n897), .A2(new_n841), .B1(new_n830), .B2(new_n1191), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(G128), .C2(new_n822), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1253), .A2(KEYINPUT59), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(KEYINPUT59), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n849), .A2(G124), .ZN(new_n1256));
  AOI211_X1 g1056(.A(G33), .B(G41), .C1(new_n902), .C2(G159), .ZN(new_n1257));
  AND4_X1   g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G116), .A2(new_n893), .B1(new_n822), .B2(G107), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n862), .B2(new_n848), .C1(new_n368), .C2(new_n824), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n304), .B(new_n424), .C1(new_n830), .C2(new_n371), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n902), .A2(G58), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n508), .B2(new_n841), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(new_n1260), .A2(new_n1068), .A3(new_n1261), .A4(new_n1263), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1264), .A2(KEYINPUT58), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(KEYINPUT58), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G50), .B1(new_n250), .B2(new_n304), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n377), .B2(G41), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n816), .B1(new_n1258), .B2(new_n1269), .ZN(new_n1270));
  XOR2_X1   g1070(.A(new_n1270), .B(KEYINPUT120), .Z(new_n1271));
  AOI211_X1 g1071(.A(new_n800), .B(new_n1271), .C1(new_n201), .C2(new_n884), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1241), .A2(new_n1059), .B1(new_n1247), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1246), .A2(new_n1273), .ZN(G375));
  AOI21_X1  g1074(.A(new_n377), .B1(new_n902), .B2(G77), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n508), .B2(new_n830), .C1(new_n531), .C2(new_n841), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n844), .A2(new_n1075), .B1(new_n848), .B2(new_n497), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n384), .A2(new_n824), .B1(new_n821), .B2(new_n862), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(new_n1276), .A2(new_n1115), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n831), .A2(G159), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n849), .A2(G128), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1262), .A3(new_n1281), .A4(new_n377), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n824), .A2(new_n356), .B1(new_n852), .B2(new_n201), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(KEYINPUT123), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(KEYINPUT123), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1282), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1288), .A2(KEYINPUT124), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n822), .A2(G137), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n1290), .B1(new_n897), .B2(new_n844), .C1(new_n841), .C2(new_n1191), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1288), .B2(KEYINPUT124), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1279), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n801), .B1(G68), .B2(new_n885), .C1(new_n1293), .C2(new_n888), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n985), .B2(new_n813), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1175), .B2(new_n1059), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1044), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1180), .A2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1296), .B1(new_n1298), .B2(new_n1299), .ZN(G381));
  NAND2_X1  g1100(.A1(new_n1241), .A2(new_n1059), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1272), .A2(new_n1247), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1213), .ZN(new_n1305));
  OR2_X1    g1105(.A1(G393), .A2(G396), .ZN(new_n1306));
  OR4_X1    g1106(.A1(G384), .A2(new_n1306), .A3(G390), .A4(G381), .ZN(new_n1307));
  OR3_X1    g1107(.A1(new_n1305), .A2(new_n1307), .A3(G387), .ZN(G407));
  OAI211_X1 g1108(.A(G407), .B(G213), .C1(G343), .C2(new_n1305), .ZN(G409));
  NAND2_X1  g1109(.A1(new_n716), .A2(G213), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1184), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1239), .A2(new_n1297), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1273), .A4(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1310), .B(new_n1314), .C1(new_n1304), .C2(new_n1213), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1172), .B1(new_n1170), .B2(new_n1150), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1154), .A2(new_n936), .A3(new_n1164), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1174), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1316), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1168), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n747), .A2(new_n757), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n770), .A2(new_n486), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n674), .B(new_n1320), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1319), .A2(new_n1323), .A3(KEYINPUT60), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT125), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1319), .A2(new_n1323), .A3(KEYINPUT125), .A4(KEYINPUT60), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT60), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n739), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1326), .A2(new_n1327), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT126), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n883), .A2(new_n1332), .A3(new_n911), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1331), .A2(new_n1296), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1333), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1337), .B1(new_n1331), .B2(new_n1296), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1334), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(KEYINPUT62), .B1(new_n1315), .B2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n716), .A2(G213), .A3(G2897), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1343), .B1(new_n1334), .B2(new_n1338), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1331), .A2(new_n1296), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1336), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1331), .A2(new_n1296), .A3(new_n1333), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1346), .A2(new_n1347), .A3(new_n1342), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1344), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT61), .B1(new_n1315), .B2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(G375), .A2(G378), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1314), .A2(new_n1310), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1351), .A2(new_n1352), .A3(new_n1353), .A4(new_n1339), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1341), .A2(new_n1350), .A3(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT127), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1060), .A2(new_n1089), .A3(G390), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(G390), .B1(new_n1060), .B2(new_n1089), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(G393), .B(G396), .ZN(new_n1360));
  NOR3_X1   g1160(.A1(new_n1358), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1360), .ZN(new_n1362));
  INV_X1    g1162(.A(G390), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(G387), .A2(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1362), .B1(new_n1364), .B2(new_n1357), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1356), .B1(new_n1361), .B2(new_n1365), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1360), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1364), .A2(new_n1362), .A3(new_n1357), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1367), .A2(KEYINPUT127), .A3(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1366), .A2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1355), .A2(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT63), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1372), .B1(new_n1315), .B2(new_n1340), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1361), .A2(new_n1365), .ZN(new_n1374));
  NAND4_X1  g1174(.A1(new_n1351), .A2(new_n1352), .A3(KEYINPUT63), .A4(new_n1339), .ZN(new_n1375));
  NAND4_X1  g1175(.A1(new_n1373), .A2(new_n1350), .A3(new_n1374), .A4(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1371), .A2(new_n1376), .ZN(G405));
  AND3_X1   g1177(.A1(new_n1351), .A2(new_n1305), .A3(new_n1340), .ZN(new_n1378));
  AOI21_X1  g1178(.A(new_n1340), .B1(new_n1351), .B2(new_n1305), .ZN(new_n1379));
  NOR3_X1   g1179(.A1(new_n1370), .A2(new_n1378), .A3(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1351), .A2(new_n1305), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1381), .A2(new_n1339), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1351), .A2(new_n1305), .A3(new_n1340), .ZN(new_n1383));
  AOI22_X1  g1183(.A1(new_n1382), .A2(new_n1383), .B1(new_n1369), .B2(new_n1366), .ZN(new_n1384));
  NOR2_X1   g1184(.A1(new_n1380), .A2(new_n1384), .ZN(G402));
endmodule


