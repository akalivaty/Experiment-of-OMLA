

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587;

  XNOR2_X1 U321 ( .A(n381), .B(n380), .ZN(n534) );
  AND2_X1 U322 ( .A1(n378), .A2(n377), .ZN(n381) );
  XNOR2_X1 U323 ( .A(n342), .B(n289), .ZN(n343) );
  XNOR2_X1 U324 ( .A(n477), .B(n476), .ZN(n520) );
  XOR2_X1 U325 ( .A(n451), .B(n398), .Z(n525) );
  XOR2_X1 U326 ( .A(n341), .B(n340), .Z(n289) );
  INV_X1 U327 ( .A(KEYINPUT95), .ZN(n387) );
  NOR2_X1 U328 ( .A1(n534), .A2(n503), .ZN(n399) );
  INV_X1 U329 ( .A(KEYINPUT37), .ZN(n475) );
  XNOR2_X1 U330 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U331 ( .A(n379), .B(KEYINPUT48), .ZN(n380) );
  XNOR2_X1 U332 ( .A(n475), .B(KEYINPUT100), .ZN(n476) );
  XNOR2_X1 U333 ( .A(n431), .B(n389), .ZN(n393) );
  XNOR2_X1 U334 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U335 ( .A(n329), .B(n328), .ZN(n372) );
  XNOR2_X1 U336 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U337 ( .A(n451), .B(n450), .Z(n527) );
  INV_X1 U338 ( .A(G43GAT), .ZN(n480) );
  XNOR2_X1 U339 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U340 ( .A(n480), .B(KEYINPUT40), .ZN(n481) );
  XNOR2_X1 U341 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n482), .B(n481), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT87), .B(KEYINPUT84), .Z(n291) );
  XNOR2_X1 U344 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n290) );
  XNOR2_X1 U345 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U346 ( .A(G22GAT), .B(G155GAT), .Z(n423) );
  XOR2_X1 U347 ( .A(n423), .B(G78GAT), .Z(n293) );
  XOR2_X1 U348 ( .A(G15GAT), .B(G1GAT), .Z(n332) );
  XNOR2_X1 U349 ( .A(n332), .B(G127GAT), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U351 ( .A(n295), .B(n294), .Z(n297) );
  NAND2_X1 U352 ( .A1(G231GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U354 ( .A(KEYINPUT15), .B(KEYINPUT85), .Z(n299) );
  XNOR2_X1 U355 ( .A(KEYINPUT86), .B(G64GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(n301), .B(n300), .Z(n306) );
  XNOR2_X1 U358 ( .A(G8GAT), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n302), .B(G211GAT), .ZN(n395) );
  XOR2_X1 U360 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n304) );
  XNOR2_X1 U361 ( .A(G71GAT), .B(G57GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n326) );
  XNOR2_X1 U363 ( .A(n395), .B(n326), .ZN(n305) );
  XOR2_X1 U364 ( .A(n306), .B(n305), .Z(n487) );
  XNOR2_X1 U365 ( .A(KEYINPUT109), .B(n487), .ZN(n564) );
  XOR2_X1 U366 ( .A(G64GAT), .B(KEYINPUT77), .Z(n308) );
  XNOR2_X1 U367 ( .A(G176GAT), .B(G204GAT), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n394) );
  XNOR2_X1 U369 ( .A(n394), .B(KEYINPUT33), .ZN(n312) );
  INV_X1 U370 ( .A(n312), .ZN(n310) );
  XOR2_X1 U371 ( .A(G120GAT), .B(KEYINPUT74), .Z(n311) );
  INV_X1 U372 ( .A(n311), .ZN(n309) );
  NAND2_X1 U373 ( .A1(n310), .A2(n309), .ZN(n314) );
  NAND2_X1 U374 ( .A1(n312), .A2(n311), .ZN(n313) );
  NAND2_X1 U375 ( .A1(n314), .A2(n313), .ZN(n316) );
  INV_X1 U376 ( .A(KEYINPUT32), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n318) );
  NAND2_X1 U379 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U381 ( .A(KEYINPUT72), .B(n319), .Z(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n329) );
  XNOR2_X1 U383 ( .A(G106GAT), .B(G78GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n322), .B(G148GAT), .ZN(n422) );
  XOR2_X1 U385 ( .A(KEYINPUT76), .B(G92GAT), .Z(n324) );
  XNOR2_X1 U386 ( .A(G99GAT), .B(KEYINPUT75), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U388 ( .A(G85GAT), .B(n325), .Z(n357) );
  XNOR2_X1 U389 ( .A(n422), .B(n357), .ZN(n327) );
  XOR2_X1 U390 ( .A(KEYINPUT41), .B(n372), .Z(n554) );
  XOR2_X1 U391 ( .A(G22GAT), .B(G197GAT), .Z(n331) );
  XNOR2_X1 U392 ( .A(G169GAT), .B(G141GAT), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n346) );
  XOR2_X1 U394 ( .A(n332), .B(G50GAT), .Z(n336) );
  XOR2_X1 U395 ( .A(G29GAT), .B(G43GAT), .Z(n334) );
  XNOR2_X1 U396 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n365) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(n365), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n344) );
  XOR2_X1 U400 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n338) );
  XNOR2_X1 U401 ( .A(G113GAT), .B(G8GAT), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n339), .B(KEYINPUT29), .ZN(n342) );
  XOR2_X1 U404 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n341) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n569) );
  INV_X1 U407 ( .A(n569), .ZN(n538) );
  AND2_X1 U408 ( .A1(n554), .A2(n538), .ZN(n348) );
  XNOR2_X1 U409 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n349) );
  NOR2_X1 U411 ( .A1(n564), .A2(n349), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n350), .B(KEYINPUT111), .ZN(n370) );
  XOR2_X1 U413 ( .A(G36GAT), .B(G190GAT), .Z(n390) );
  XOR2_X1 U414 ( .A(KEYINPUT10), .B(KEYINPUT81), .Z(n352) );
  XNOR2_X1 U415 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U417 ( .A(n390), .B(n353), .Z(n355) );
  NAND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n369) );
  XOR2_X1 U421 ( .A(KEYINPUT82), .B(KEYINPUT9), .Z(n359) );
  XNOR2_X1 U422 ( .A(G134GAT), .B(G106GAT), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U424 ( .A(KEYINPUT83), .B(KEYINPUT66), .Z(n361) );
  XNOR2_X1 U425 ( .A(KEYINPUT80), .B(KEYINPUT67), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U427 ( .A(n363), .B(n362), .Z(n367) );
  XNOR2_X1 U428 ( .A(G50GAT), .B(KEYINPUT79), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n364), .B(G162GAT), .ZN(n426) );
  XNOR2_X1 U430 ( .A(n365), .B(n426), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n561) );
  NOR2_X1 U433 ( .A1(n370), .A2(n561), .ZN(n371) );
  XNOR2_X1 U434 ( .A(KEYINPUT47), .B(n371), .ZN(n378) );
  BUF_X1 U435 ( .A(n372), .Z(n575) );
  XOR2_X1 U436 ( .A(KEYINPUT36), .B(n561), .Z(n585) );
  NOR2_X1 U437 ( .A1(n585), .A2(n487), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n373), .B(KEYINPUT45), .ZN(n374) );
  NAND2_X1 U439 ( .A1(n374), .A2(n569), .ZN(n375) );
  NOR2_X1 U440 ( .A1(n575), .A2(n375), .ZN(n376) );
  XOR2_X1 U441 ( .A(KEYINPUT112), .B(n376), .Z(n377) );
  XOR2_X1 U442 ( .A(KEYINPUT64), .B(KEYINPUT113), .Z(n379) );
  XOR2_X1 U443 ( .A(KEYINPUT89), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U444 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U446 ( .A(G169GAT), .B(n384), .Z(n451) );
  XOR2_X1 U447 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n386) );
  XNOR2_X1 U448 ( .A(G197GAT), .B(G218GAT), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n431) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U451 ( .A(G92GAT), .B(n390), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n391), .B(KEYINPUT94), .ZN(n392) );
  XOR2_X1 U453 ( .A(n393), .B(n392), .Z(n397) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  INV_X1 U456 ( .A(n525), .ZN(n503) );
  XNOR2_X1 U457 ( .A(n399), .B(KEYINPUT54), .ZN(n418) );
  XOR2_X1 U458 ( .A(G57GAT), .B(KEYINPUT6), .Z(n401) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n409) );
  XOR2_X1 U461 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n407) );
  XOR2_X1 U462 ( .A(G127GAT), .B(G134GAT), .Z(n403) );
  XNOR2_X1 U463 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U465 ( .A(G113GAT), .B(n404), .Z(n442) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n405), .B(KEYINPUT2), .ZN(n432) );
  XNOR2_X1 U468 ( .A(n442), .B(n432), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n417) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XOR2_X1 U472 ( .A(KEYINPUT93), .B(G85GAT), .Z(n411) );
  XNOR2_X1 U473 ( .A(G148GAT), .B(G155GAT), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n413) );
  XOR2_X1 U475 ( .A(G29GAT), .B(G162GAT), .Z(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U478 ( .A(n417), .B(n416), .Z(n522) );
  INV_X1 U479 ( .A(n522), .ZN(n500) );
  NAND2_X1 U480 ( .A1(n418), .A2(n500), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n419), .B(KEYINPUT65), .ZN(n568) );
  XOR2_X1 U482 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n421) );
  XNOR2_X1 U483 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n436) );
  XOR2_X1 U485 ( .A(n423), .B(n422), .Z(n425) );
  XNOR2_X1 U486 ( .A(G211GAT), .B(G204GAT), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n430) );
  XOR2_X1 U488 ( .A(n426), .B(KEYINPUT24), .Z(n428) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U491 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U494 ( .A(n436), .B(n435), .Z(n465) );
  NAND2_X1 U495 ( .A1(n568), .A2(n465), .ZN(n438) );
  XOR2_X1 U496 ( .A(KEYINPUT118), .B(KEYINPUT55), .Z(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n452) );
  XOR2_X1 U498 ( .A(KEYINPUT88), .B(G176GAT), .Z(n440) );
  XNOR2_X1 U499 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n449) );
  XOR2_X1 U502 ( .A(G71GAT), .B(G99GAT), .Z(n444) );
  XNOR2_X1 U503 ( .A(G43GAT), .B(G190GAT), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U505 ( .A(G183GAT), .B(n445), .Z(n447) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U509 ( .A(n527), .ZN(n537) );
  NOR2_X1 U510 ( .A1(n452), .A2(n537), .ZN(n454) );
  INV_X1 U511 ( .A(KEYINPUT119), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n565) );
  NAND2_X1 U513 ( .A1(n565), .A2(n538), .ZN(n456) );
  XNOR2_X1 U514 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(G1348GAT) );
  NAND2_X1 U516 ( .A1(n565), .A2(n561), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n575), .A2(n569), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT78), .B(n459), .Z(n491) );
  XNOR2_X1 U519 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n460) );
  XOR2_X1 U520 ( .A(n460), .B(n525), .Z(n467) );
  NOR2_X1 U521 ( .A1(n467), .A2(n500), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT97), .ZN(n533) );
  XOR2_X1 U523 ( .A(n465), .B(KEYINPUT28), .Z(n530) );
  INV_X1 U524 ( .A(n530), .ZN(n535) );
  NAND2_X1 U525 ( .A1(n537), .A2(n535), .ZN(n462) );
  NOR2_X1 U526 ( .A1(n533), .A2(n462), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n527), .A2(n525), .ZN(n463) );
  NAND2_X1 U528 ( .A1(n465), .A2(n463), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n464), .B(KEYINPUT25), .ZN(n469) );
  NOR2_X1 U530 ( .A1(n465), .A2(n527), .ZN(n466) );
  XOR2_X1 U531 ( .A(n466), .B(KEYINPUT26), .Z(n550) );
  NOR2_X1 U532 ( .A1(n467), .A2(n550), .ZN(n468) );
  NOR2_X1 U533 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U534 ( .A1(n522), .A2(n470), .ZN(n471) );
  NOR2_X1 U535 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U536 ( .A(KEYINPUT98), .B(n473), .Z(n489) );
  INV_X1 U537 ( .A(n487), .ZN(n578) );
  NOR2_X1 U538 ( .A1(n578), .A2(n585), .ZN(n474) );
  NAND2_X1 U539 ( .A1(n489), .A2(n474), .ZN(n477) );
  NOR2_X1 U540 ( .A1(n491), .A2(n520), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n478), .B(KEYINPUT101), .ZN(n479) );
  XNOR2_X1 U542 ( .A(KEYINPUT38), .B(n479), .ZN(n505) );
  NOR2_X1 U543 ( .A1(n505), .A2(n537), .ZN(n482) );
  XOR2_X1 U544 ( .A(n554), .B(KEYINPUT103), .Z(n540) );
  NAND2_X1 U545 ( .A1(n540), .A2(n565), .ZN(n486) );
  XOR2_X1 U546 ( .A(G176GAT), .B(KEYINPUT57), .Z(n484) );
  XOR2_X1 U547 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n483) );
  XNOR2_X1 U548 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(G1349GAT) );
  NOR2_X1 U550 ( .A1(n561), .A2(n487), .ZN(n488) );
  XNOR2_X1 U551 ( .A(KEYINPUT16), .B(n488), .ZN(n490) );
  NAND2_X1 U552 ( .A1(n490), .A2(n489), .ZN(n507) );
  NOR2_X1 U553 ( .A1(n491), .A2(n507), .ZN(n498) );
  NAND2_X1 U554 ( .A1(n498), .A2(n522), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(KEYINPUT34), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  NAND2_X1 U557 ( .A1(n498), .A2(n525), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n496) );
  NAND2_X1 U560 ( .A1(n498), .A2(n527), .ZN(n495) );
  XNOR2_X1 U561 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U562 ( .A(G15GAT), .B(n497), .Z(G1326GAT) );
  NAND2_X1 U563 ( .A1(n498), .A2(n530), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U565 ( .A1(n505), .A2(n500), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n505), .A2(n503), .ZN(n504) );
  XOR2_X1 U569 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U570 ( .A1(n505), .A2(n535), .ZN(n506) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  XOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT102), .Z(n509) );
  NAND2_X1 U573 ( .A1(n540), .A2(n569), .ZN(n519) );
  NOR2_X1 U574 ( .A1(n519), .A2(n507), .ZN(n515) );
  NAND2_X1 U575 ( .A1(n515), .A2(n522), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U577 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n525), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT105), .Z(n514) );
  NAND2_X1 U582 ( .A1(n515), .A2(n527), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U585 ( .A1(n515), .A2(n530), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n524) );
  NOR2_X1 U589 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U590 ( .A(KEYINPUT107), .B(n521), .Z(n529) );
  NAND2_X1 U591 ( .A1(n522), .A2(n529), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n525), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n529), .A2(n527), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n532) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n551), .A2(n535), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n538), .A2(n546), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U606 ( .A1(n546), .A2(n540), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n544) );
  NAND2_X1 U609 ( .A1(n546), .A2(n564), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n545), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n561), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n549), .Z(G1343GAT) );
  INV_X1 U616 ( .A(n550), .ZN(n567) );
  NAND2_X1 U617 ( .A1(n551), .A2(n567), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n569), .A2(n553), .ZN(n552) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n556) );
  INV_X1 U621 ( .A(n553), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n562), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(n557), .B(KEYINPUT52), .Z(n559) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n578), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n584) );
  NOR2_X1 U634 ( .A1(n569), .A2(n584), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT122), .B(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U641 ( .A(n584), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT124), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n583) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

