//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G77), .A2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n215), .B(new_n219), .C1(G116), .C2(G270), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G50), .A2(G226), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  INV_X1    g0032(.A(G13), .ZN(new_n233));
  OAI21_X1  g0033(.A(KEYINPUT64), .B1(new_n206), .B2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(KEYINPUT64), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n235), .A2(G1), .A3(G13), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n238), .A2(new_n207), .ZN(new_n239));
  OAI21_X1  g0039(.A(G50), .B1(G58), .B2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  AOI211_X1 g0041(.A(new_n212), .B(new_n232), .C1(new_n239), .C2(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n224), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT2), .B(G226), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G250), .B(G257), .Z(new_n247));
  XNOR2_X1  g0047(.A(G264), .B(G270), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g0053(.A(new_n253), .B(KEYINPUT65), .Z(new_n254));
  XOR2_X1   g0054(.A(G87), .B(G97), .Z(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  NAND2_X1  g0058(.A1(new_n228), .A2(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G77), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n259), .B1(new_n261), .B2(new_n202), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n234), .A2(new_n236), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT11), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n233), .A2(G1), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n259), .ZN(new_n274));
  XOR2_X1   g0074(.A(new_n274), .B(KEYINPUT12), .Z(new_n275));
  AOI21_X1  g0075(.A(new_n268), .B1(new_n206), .B2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n275), .B1(new_n277), .B2(new_n228), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G97), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n224), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  OAI211_X1 g0088(.A(G226), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n292), .A2(KEYINPUT69), .A3(G226), .A4(new_n286), .ZN(new_n293));
  AOI221_X4 g0093(.A(new_n282), .B1(G1698), .B2(new_n285), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n237), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n280), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT66), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(G1), .A2(G13), .ZN(new_n303));
  NAND3_X1  g0103(.A1(KEYINPUT66), .A2(G33), .A3(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n305), .A2(new_n298), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n300), .B1(new_n306), .B2(G238), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n291), .A2(new_n293), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n285), .A2(G1698), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n281), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n296), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(KEYINPUT70), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n297), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT13), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n297), .A2(new_n315), .A3(new_n307), .A4(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n279), .B1(new_n317), .B2(G200), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n314), .A2(G190), .A3(new_n316), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(G179), .A3(new_n316), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT71), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n314), .A2(new_n323), .A3(G179), .A4(new_n316), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n291), .A2(new_n293), .B1(G1698), .B2(new_n285), .ZN(new_n327));
  AOI211_X1 g0127(.A(new_n280), .B(new_n296), .C1(new_n327), .C2(new_n281), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT70), .B1(new_n310), .B2(new_n311), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n315), .B1(new_n330), .B2(new_n307), .ZN(new_n331));
  INV_X1    g0131(.A(new_n316), .ZN(new_n332));
  OAI21_X1  g0132(.A(G169), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n317), .A2(new_n335), .A3(G169), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT72), .B1(new_n326), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n335), .B1(new_n317), .B2(G169), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  AOI211_X1 g0140(.A(KEYINPUT14), .B(new_n340), .C1(new_n314), .C2(new_n316), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(new_n325), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n320), .B1(new_n345), .B2(new_n279), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT8), .B(G58), .Z(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT68), .Z(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT15), .B(G87), .Z(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n264), .B2(new_n351), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n233), .A2(new_n207), .A3(G1), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n352), .A2(new_n268), .B1(new_n265), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n276), .A2(G77), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n300), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n306), .A2(G244), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n292), .A2(G1698), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n359), .A2(new_n229), .B1(new_n225), .B2(new_n292), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n286), .B2(new_n285), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n357), .B(new_n358), .C1(new_n361), .C2(new_n296), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n340), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(G179), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n356), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n346), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n353), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n202), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n276), .B2(new_n202), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT67), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n203), .A2(G20), .ZN(new_n372));
  INV_X1    g0172(.A(G150), .ZN(new_n373));
  INV_X1    g0173(.A(new_n347), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n372), .B1(new_n373), .B2(new_n261), .C1(new_n374), .C2(new_n264), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n268), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT9), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(G222), .A2(G1698), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n286), .A2(G223), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n292), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n311), .B(new_n382), .C1(G77), .C2(new_n292), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n306), .A2(G226), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n357), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G200), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n371), .A2(KEYINPUT9), .A3(new_n376), .ZN(new_n387));
  INV_X1    g0187(.A(G190), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n379), .A2(new_n386), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT10), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n385), .A2(new_n340), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n385), .A2(G179), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n377), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(G223), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT75), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n292), .A2(KEYINPUT75), .A3(G223), .A4(new_n286), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n292), .A2(G226), .A3(G1698), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n311), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n305), .A2(G232), .A3(new_n298), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n357), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT76), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n398), .A2(new_n399), .A3(new_n402), .A4(new_n401), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n406), .B1(new_n411), .B2(new_n311), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT76), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n414), .A2(G200), .B1(G190), .B2(new_n408), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n347), .A2(new_n353), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n277), .B2(new_n347), .ZN(new_n417));
  XNOR2_X1  g0217(.A(G58), .B(G68), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n287), .A2(new_n288), .A3(new_n420), .A4(G20), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n228), .B1(new_n421), .B2(KEYINPUT73), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n283), .A2(new_n207), .A3(new_n284), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n420), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT73), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n283), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n284), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n422), .A2(new_n427), .A3(KEYINPUT74), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT74), .B1(new_n422), .B2(new_n427), .ZN(new_n429));
  OAI211_X1 g0229(.A(KEYINPUT16), .B(new_n419), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n268), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n424), .A2(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G68), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n419), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT16), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n417), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n415), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT17), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n410), .A2(new_n340), .A3(new_n413), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n408), .A2(G179), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n437), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT18), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n395), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n362), .A2(new_n388), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n362), .A2(G200), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n354), .A2(new_n448), .A3(new_n355), .A4(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n366), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G41), .ZN(new_n455));
  INV_X1    g0255(.A(G41), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT5), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n455), .A2(new_n457), .A3(new_n206), .A4(G45), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n458), .A2(new_n305), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G257), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n456), .A2(KEYINPUT5), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n462));
  INV_X1    g0262(.A(new_n457), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(KEYINPUT80), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n463), .A2(KEYINPUT80), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT79), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n359), .B2(new_n214), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n292), .A2(G244), .A3(new_n286), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT4), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT4), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n292), .A2(new_n472), .A3(G244), .A4(new_n286), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n460), .B(new_n466), .C1(new_n474), .C2(new_n296), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G200), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n475), .A2(new_n388), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n262), .A2(G1), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n268), .A2(new_n353), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G97), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n367), .A2(G97), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT78), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n217), .A2(new_n225), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G97), .A2(G107), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g0289(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n490));
  NAND2_X1  g0290(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(G107), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n486), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n485), .B(KEYINPUT78), .C1(new_n488), .C2(new_n487), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G20), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n432), .A2(G107), .B1(G77), .B2(new_n260), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n483), .B(new_n484), .C1(new_n498), .C2(new_n268), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n475), .A2(KEYINPUT81), .A3(G200), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n478), .A2(new_n479), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n268), .ZN(new_n502));
  INV_X1    g0302(.A(new_n484), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n482), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n475), .A2(new_n340), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n471), .A2(new_n473), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n311), .B1(new_n506), .B2(new_n469), .ZN(new_n507));
  INV_X1    g0307(.A(G179), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(new_n460), .A4(new_n466), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n501), .A2(KEYINPUT82), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT79), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n467), .B(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n207), .B1(new_n217), .B2(G33), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G20), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n515), .A2(KEYINPUT20), .A3(new_n268), .A4(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT20), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n513), .A2(new_n514), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n268), .A2(new_n517), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n481), .A2(G116), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n273), .A2(new_n517), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G200), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n292), .A2(G257), .A3(new_n286), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n287), .A2(new_n288), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G303), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n531), .C1(new_n359), .C2(new_n226), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n311), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n459), .A2(G270), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n466), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT85), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n532), .A2(new_n311), .B1(new_n465), .B2(new_n464), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT85), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(new_n534), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n528), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n535), .A2(KEYINPUT85), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n537), .B2(new_n534), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n527), .B(new_n540), .C1(G190), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n367), .A2(new_n350), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n292), .A2(new_n207), .A3(G68), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT84), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n263), .A2(new_n548), .A3(G97), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n488), .A2(new_n213), .B1(new_n281), .B2(new_n207), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n548), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n292), .A2(new_n552), .A3(new_n207), .A4(G68), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n545), .B1(new_n554), .B2(new_n268), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n481), .A2(new_n350), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G45), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n305), .B(G250), .C1(G1), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n462), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT83), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n292), .B1(G238), .B2(G1698), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n286), .A2(G244), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(new_n262), .B2(new_n516), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n311), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT83), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(new_n566), .A3(new_n462), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n561), .A2(new_n565), .A3(new_n508), .A4(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n561), .A2(new_n565), .A3(new_n567), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n557), .B(new_n568), .C1(new_n569), .C2(G169), .ZN(new_n570));
  NOR4_X1   g0370(.A1(new_n268), .A2(new_n213), .A3(new_n353), .A4(new_n480), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n545), .B(new_n571), .C1(new_n554), .C2(new_n268), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n561), .A2(new_n565), .A3(G190), .A4(new_n567), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n569), .C2(new_n528), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n292), .A2(G250), .A3(new_n286), .ZN(new_n575));
  INV_X1    g0375(.A(G294), .ZN(new_n576));
  OAI221_X1 g0376(.A(new_n575), .B1(new_n262), .B2(new_n576), .C1(new_n359), .C2(new_n218), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n311), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n459), .A2(G264), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n466), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G200), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT86), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n207), .B2(G107), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n263), .A2(G116), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n584), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n292), .A2(new_n207), .A3(G87), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n588), .B(KEYINPUT24), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n268), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n481), .A2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n272), .A2(G20), .A3(new_n225), .ZN(new_n598));
  XOR2_X1   g0398(.A(new_n598), .B(KEYINPUT25), .Z(new_n599));
  NAND4_X1  g0399(.A1(new_n581), .A2(new_n596), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n580), .A2(new_n388), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n570), .B(new_n574), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n544), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n580), .A2(G169), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n578), .A2(G179), .A3(new_n466), .A4(new_n579), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n527), .A2(G179), .A3(new_n534), .A4(new_n537), .ZN(new_n609));
  OAI211_X1 g0409(.A(G169), .B(new_n527), .C1(new_n541), .C2(new_n542), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n340), .B1(new_n536), .B2(new_n539), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n527), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n608), .B(new_n609), .C1(new_n611), .C2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT82), .B1(new_n501), .B2(new_n510), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n453), .A2(new_n511), .A3(new_n603), .A4(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n394), .ZN(new_n619));
  INV_X1    g0419(.A(new_n279), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n338), .B2(new_n344), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n320), .A2(new_n365), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n439), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n445), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n619), .B1(new_n624), .B2(new_n391), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT88), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n510), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n570), .A2(new_n574), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n504), .A2(new_n509), .A3(KEYINPUT88), .A4(new_n505), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n570), .A2(new_n574), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT26), .B1(new_n632), .B2(new_n510), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n631), .A2(new_n570), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n501), .A2(new_n510), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n602), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n613), .A2(new_n612), .A3(new_n527), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n608), .A2(KEYINPUT87), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT87), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n604), .A2(new_n607), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n639), .A2(new_n640), .A3(new_n609), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n625), .B1(new_n452), .B2(new_n645), .ZN(G369));
  NAND2_X1  g0446(.A1(new_n272), .A2(new_n207), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n647), .A2(KEYINPUT89), .A3(KEYINPUT27), .ZN(new_n648));
  INV_X1    g0448(.A(G213), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n647), .B2(KEYINPUT27), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT89), .B1(new_n647), .B2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n640), .B2(new_n642), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n639), .A2(new_n609), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n654), .ZN(new_n658));
  INV_X1    g0458(.A(new_n608), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n600), .A2(new_n601), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n655), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n656), .A2(new_n544), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n527), .B2(new_n654), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n657), .A2(new_n527), .A3(new_n654), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT90), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n604), .A2(new_n654), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n661), .A2(new_n669), .B1(new_n659), .B2(new_n654), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n662), .B1(new_n668), .B2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n210), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G1), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n488), .A2(new_n213), .A3(new_n516), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n675), .A2(new_n676), .B1(new_n240), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n654), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n617), .A2(new_n511), .A3(new_n603), .A4(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n606), .A2(new_n535), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n507), .A2(new_n460), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n569), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  AOI21_X1  g0487(.A(G179), .B1(new_n536), .B2(new_n539), .ZN(new_n688));
  INV_X1    g0488(.A(new_n569), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n688), .A2(new_n475), .A3(new_n689), .A4(new_n580), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n686), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n681), .A2(KEYINPUT31), .B1(new_n654), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n679), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n632), .A2(new_n510), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n628), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n570), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n699), .B1(KEYINPUT26), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n636), .A2(new_n615), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n654), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n654), .B1(new_n634), .B2(new_n644), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(KEYINPUT29), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n696), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n678), .B1(new_n708), .B2(G1), .ZN(G364));
  NOR2_X1   g0509(.A1(new_n233), .A2(G20), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G45), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n674), .A2(G1), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT91), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n668), .B(new_n714), .C1(G330), .C2(new_n666), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT100), .Z(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n664), .B2(new_n665), .ZN(new_n720));
  NAND3_X1  g0520(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT96), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n388), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(G190), .ZN(new_n724));
  XNOR2_X1  g0524(.A(KEYINPUT33), .B(G317), .ZN(new_n725));
  AOI22_X1  g0525(.A1(G326), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G322), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n207), .B2(new_n508), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n388), .A2(G200), .ZN(new_n730));
  NAND3_X1  g0530(.A1(KEYINPUT95), .A2(G20), .A3(G179), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n726), .B(new_n530), .C1(new_n727), .C2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n207), .A2(G179), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G190), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n733), .B1(G329), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(G190), .A3(G200), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT98), .Z(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G303), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n729), .A2(new_n735), .A3(new_n731), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n734), .A2(new_n388), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n744), .A2(G311), .B1(new_n746), .B2(G283), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n730), .A2(new_n508), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G294), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n738), .A2(new_n742), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n745), .A2(new_n225), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(G97), .B2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(new_n723), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n753), .B1(new_n213), .B2(new_n739), .C1(new_n754), .C2(new_n202), .ZN(new_n755));
  INV_X1    g0555(.A(new_n732), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n530), .B(new_n755), .C1(G58), .C2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT97), .B(G159), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n737), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(KEYINPUT32), .B1(new_n744), .B2(G77), .ZN(new_n760));
  INV_X1    g0560(.A(new_n724), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n757), .B(new_n760), .C1(new_n228), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n759), .A2(KEYINPUT32), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n751), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT99), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n238), .B1(G20), .B2(new_n340), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n672), .A2(new_n292), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G45), .B2(new_n240), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT93), .Z(new_n770));
  INV_X1    g0570(.A(new_n253), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n558), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n672), .A2(new_n530), .ZN(new_n773));
  XNOR2_X1  g0573(.A(G355), .B(KEYINPUT92), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n772), .B(new_n775), .C1(G116), .C2(new_n210), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT94), .Z(new_n777));
  NOR2_X1   g0577(.A1(new_n766), .A2(new_n718), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n720), .A2(new_n713), .A3(new_n767), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n715), .A2(new_n780), .ZN(G396));
  NAND2_X1  g0581(.A1(new_n356), .A2(new_n654), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n450), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n365), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n356), .A2(new_n363), .A3(new_n364), .A4(new_n680), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n705), .B(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n695), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n714), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n761), .A2(new_n791), .B1(new_n516), .B2(new_n743), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n756), .A2(G294), .B1(new_n749), .B2(G97), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT102), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(G107), .C2(new_n741), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n746), .A2(G87), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n723), .A2(G303), .B1(G311), .B2(new_n737), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n795), .A2(new_n530), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G137), .A2(new_n723), .B1(new_n724), .B2(G150), .ZN(new_n799));
  INV_X1    g0599(.A(G143), .ZN(new_n800));
  INV_X1    g0600(.A(new_n758), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n732), .C1(new_n801), .C2(new_n743), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT34), .Z(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G50), .B2(new_n741), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n746), .A2(G68), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n292), .B1(new_n736), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT103), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n807), .A2(new_n808), .B1(new_n749), .B2(G58), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n804), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n798), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n766), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n766), .A2(new_n716), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n714), .B1(new_n265), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(KEYINPUT101), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n786), .A2(new_n716), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n815), .A2(KEYINPUT101), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n813), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n790), .A2(new_n819), .ZN(G384));
  XNOR2_X1  g0620(.A(new_n694), .B(KEYINPUT113), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n693), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n366), .A2(new_n451), .A3(G330), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n786), .B1(new_n693), .B2(new_n822), .ZN(new_n825));
  INV_X1    g0625(.A(new_n430), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n419), .B1(new_n428), .B2(new_n429), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n431), .B1(new_n827), .B2(new_n435), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n826), .B1(new_n828), .B2(KEYINPUT105), .ZN(new_n829));
  INV_X1    g0629(.A(new_n419), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT74), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n832));
  OAI21_X1  g0632(.A(G68), .B1(new_n426), .B2(new_n425), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n422), .A2(new_n427), .A3(KEYINPUT74), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n268), .B1(new_n836), .B2(KEYINPUT16), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT105), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n417), .B1(new_n829), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT106), .B1(new_n840), .B2(new_n652), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n409), .B(new_n406), .C1(new_n311), .C2(new_n411), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT76), .B1(new_n404), .B2(new_n407), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(new_n528), .B1(new_n388), .B2(new_n412), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n430), .A2(new_n436), .ZN(new_n846));
  INV_X1    g0646(.A(new_n417), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(KEYINPUT105), .B(new_n268), .C1(new_n836), .C2(KEYINPUT16), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n430), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n827), .A2(new_n435), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT105), .B1(new_n852), .B2(new_n268), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n847), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n441), .B1(new_n844), .B2(new_n340), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT106), .ZN(new_n857));
  INV_X1    g0657(.A(new_n652), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n841), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT108), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n848), .B2(new_n858), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n437), .A2(KEYINPUT108), .A3(new_n652), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT107), .B1(new_n443), .B2(new_n437), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT107), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n855), .A2(new_n848), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n869), .A3(new_n438), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT109), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n444), .A2(new_n868), .B1(new_n415), .B2(new_n437), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n848), .A2(new_n863), .A3(new_n858), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT108), .B1(new_n437), .B2(new_n652), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT37), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT109), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n872), .A2(new_n875), .A3(new_n876), .A4(new_n867), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n861), .A2(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n439), .A2(new_n445), .B1(new_n841), .B2(new_n859), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT111), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n444), .B1(new_n849), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n873), .A2(new_n874), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n885), .B(new_n886), .C1(new_n884), .C2(new_n849), .ZN(new_n887));
  AOI22_X1  g0687(.A1(KEYINPUT37), .A2(new_n887), .B1(new_n871), .B2(new_n877), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n439), .B2(new_n445), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n883), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  AND4_X1   g0691(.A1(new_n343), .A2(new_n325), .A3(new_n334), .A4(new_n336), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n343), .B1(new_n342), .B2(new_n325), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n279), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n320), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n279), .A2(new_n654), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n621), .A2(new_n654), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n825), .A2(new_n891), .A3(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n346), .A2(new_n896), .B1(new_n621), .B2(new_n654), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n787), .B1(new_n692), .B2(new_n821), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n860), .A2(KEYINPUT37), .B1(new_n871), .B2(new_n877), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n883), .B1(new_n904), .B2(new_n880), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT40), .B1(new_n882), .B2(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(KEYINPUT40), .A2(new_n900), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n824), .B1(new_n907), .B2(new_n679), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n903), .B2(new_n891), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n906), .A2(new_n825), .A3(new_n899), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n823), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n908), .B1(new_n452), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n785), .B(KEYINPUT104), .Z(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n705), .B2(new_n787), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n897), .B2(new_n898), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n904), .A2(new_n883), .A3(new_n880), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n879), .B2(new_n881), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n445), .B2(new_n858), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT39), .B1(new_n918), .B2(new_n917), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT110), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n882), .A2(new_n890), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n882), .B2(new_n905), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT110), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n894), .A2(new_n654), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n920), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n913), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n625), .B1(new_n706), .B2(new_n452), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT112), .Z(new_n933));
  XNOR2_X1  g0733(.A(new_n931), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n206), .B2(new_n710), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n516), .B1(new_n495), .B2(KEYINPUT35), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(new_n239), .C1(KEYINPUT35), .C2(new_n495), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  OAI21_X1  g0738(.A(G77), .B1(new_n223), .B2(new_n228), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n939), .A2(new_n240), .B1(G50), .B2(new_n228), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(G1), .A3(new_n233), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n935), .A2(new_n938), .A3(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n658), .A2(new_n661), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n635), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT42), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n501), .B(new_n510), .C1(new_n499), .C2(new_n680), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n510), .B1(new_n946), .B2(new_n608), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n680), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n572), .A2(new_n680), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n629), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n570), .A2(new_n950), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n953), .ZN(new_n955));
  XOR2_X1   g0755(.A(KEYINPUT114), .B(KEYINPUT43), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n957), .B2(new_n949), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n668), .A2(new_n670), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n946), .B1(new_n510), .B2(new_n680), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n959), .B(new_n962), .Z(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT115), .B(KEYINPUT41), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n673), .B(new_n964), .Z(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n662), .A2(new_n961), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT45), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n662), .A2(new_n961), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT116), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT117), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(KEYINPUT116), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n960), .A4(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n670), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n943), .B1(new_n976), .B2(new_n658), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n668), .B(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n707), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n972), .A2(new_n960), .A3(new_n974), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n960), .A2(new_n971), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(KEYINPUT117), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n975), .B(new_n979), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n966), .B1(new_n983), .B2(new_n708), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n711), .A2(G1), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n963), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n714), .B1(new_n955), .B2(new_n719), .ZN(new_n987));
  INV_X1    g0787(.A(new_n768), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n778), .B1(new_n210), .B2(new_n351), .C1(new_n988), .C2(new_n249), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n761), .A2(new_n801), .B1(new_n202), .B2(new_n743), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT118), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n990), .A2(new_n991), .B1(G68), .B2(new_n749), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n265), .B2(new_n745), .C1(new_n800), .C2(new_n754), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n292), .B1(new_n732), .B2(new_n373), .ZN(new_n995));
  INV_X1    g0795(.A(G137), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n739), .A2(new_n223), .B1(new_n736), .B2(new_n996), .ZN(new_n997));
  NOR4_X1   g0797(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n723), .A2(G311), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT46), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n740), .A2(new_n1000), .A3(new_n516), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G294), .B2(new_n724), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n749), .A2(G107), .B1(new_n737), .B2(G317), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1000), .B1(new_n739), .B2(new_n516), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1002), .A2(new_n530), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(G303), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n791), .A2(new_n743), .B1(new_n732), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n745), .A2(new_n217), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n998), .B1(new_n999), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT47), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n766), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n987), .B(new_n989), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n986), .A2(new_n1013), .ZN(G387));
  NAND2_X1  g0814(.A1(new_n670), .A2(new_n719), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n246), .A2(new_n558), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1016), .A2(new_n768), .B1(new_n676), .B2(new_n773), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n347), .A2(new_n202), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n558), .B1(new_n228), .B2(new_n265), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1019), .A2(new_n676), .A3(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1017), .A2(new_n1021), .B1(G107), .B2(new_n210), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n714), .B1(new_n1022), .B2(new_n778), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n749), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n351), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G159), .B2(new_n723), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n228), .B2(new_n743), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n347), .B2(new_n724), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n739), .A2(new_n265), .B1(new_n736), .B2(new_n373), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1029), .A2(new_n1008), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n756), .A2(G50), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n292), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G311), .A2(new_n724), .B1(new_n723), .B2(G322), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1006), .B2(new_n743), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G317), .B2(new_n756), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT48), .Z(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n791), .B2(new_n1024), .C1(new_n576), .C2(new_n739), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT49), .Z(new_n1038));
  AOI21_X1  g0838(.A(new_n292), .B1(new_n737), .B2(G326), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n516), .B2(new_n745), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1032), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT119), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1015), .B(new_n1023), .C1(new_n1042), .C2(new_n1012), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n985), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n978), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n673), .B1(new_n1045), .B2(new_n708), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1043), .B1(new_n1044), .B2(new_n978), .C1(new_n1046), .C2(new_n979), .ZN(G393));
  XNOR2_X1  g0847(.A(new_n960), .B(new_n971), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n707), .B2(new_n978), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n983), .A2(new_n673), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n796), .A2(new_n292), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1024), .A2(new_n265), .B1(new_n800), .B2(new_n736), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n761), .A2(new_n202), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n756), .A2(G159), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n754), .B2(new_n373), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT51), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1052), .B(new_n1053), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .C1(new_n228), .C2(new_n739), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1051), .B(new_n1058), .C1(new_n347), .C2(new_n744), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n530), .B1(new_n736), .B2(new_n727), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n723), .A2(G317), .B1(new_n756), .B2(G311), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  NOR2_X1   g0862(.A1(new_n739), .A2(new_n791), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n752), .B(new_n1063), .C1(G116), .C2(new_n749), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1062), .B(new_n1064), .C1(new_n576), .C2(new_n743), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1060), .B(new_n1065), .C1(G303), .C2(new_n724), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n766), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n778), .B1(new_n217), .B2(new_n210), .C1(new_n988), .C2(new_n257), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n946), .B(new_n718), .C1(new_n510), .C2(new_n680), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1067), .A2(new_n713), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1048), .B2(new_n1044), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT120), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1050), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(G390));
  XNOR2_X1  g0874(.A(new_n925), .B(KEYINPUT110), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT121), .B1(new_n916), .B2(new_n929), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n929), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n901), .C2(new_n915), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1075), .A2(new_n924), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n695), .A2(new_n899), .A3(new_n787), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n914), .B1(new_n703), .B2(new_n787), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n891), .B(new_n1078), .C1(new_n901), .C2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1080), .A2(KEYINPUT122), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT122), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1079), .A2(new_n1076), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1083), .B1(new_n928), .B2(new_n1086), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n901), .A2(new_n679), .A3(new_n902), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1081), .B(new_n1083), .C1(new_n928), .C2(new_n1086), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1084), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n824), .B(new_n625), .C1(new_n452), .C2(new_n706), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n915), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n899), .B1(new_n695), .B2(new_n787), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n901), .B1(new_n679), .B2(new_n902), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1093), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1092), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1084), .B(new_n1099), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n673), .A3(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n985), .B(new_n1084), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1075), .A2(new_n716), .A3(new_n924), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n814), .A2(new_n374), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n292), .B1(new_n756), .B2(G116), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1107), .B(new_n805), .C1(new_n217), .C2(new_n743), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n741), .A2(G87), .B1(G283), .B2(new_n723), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1109), .B1(new_n265), .B2(new_n1024), .C1(new_n225), .C2(new_n761), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1108), .B(new_n1110), .C1(G294), .C2(new_n737), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n749), .A2(G159), .B1(new_n737), .B2(G125), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT53), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n739), .A2(new_n373), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .C1(new_n743), .C2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n724), .A2(G137), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n530), .B1(new_n746), .B2(G50), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n754), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1117), .B(new_n1121), .C1(G132), .C2(new_n756), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n766), .B1(new_n1111), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1105), .A2(new_n713), .A3(new_n1106), .A4(new_n1123), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1104), .A2(new_n1124), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1103), .A2(KEYINPUT123), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT123), .B1(new_n1103), .B2(new_n1125), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1126), .A2(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(new_n1093), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1102), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n377), .A2(new_n858), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT124), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n395), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n391), .A2(KEYINPUT124), .A3(new_n394), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n907), .B2(new_n679), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1141), .B(G330), .C1(new_n910), .C2(new_n911), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1143), .A2(new_n930), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n930), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1130), .A2(KEYINPUT57), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT125), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1150), .A2(new_n1151), .B1(new_n1102), .B2(new_n1129), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1148), .B(new_n673), .C1(new_n1152), .C2(KEYINPUT57), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1141), .A2(new_n717), .ZN(new_n1154));
  INV_X1    g0954(.A(G124), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n262), .B1(new_n736), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n723), .A2(G125), .B1(new_n744), .B2(G137), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1120), .B2(new_n732), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n761), .A2(new_n806), .B1(new_n739), .B2(new_n1116), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n373), .B2(new_n1024), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G41), .B(new_n1156), .C1(new_n1161), .C2(KEYINPUT59), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(KEYINPUT59), .B2(new_n1161), .C1(new_n801), .C2(new_n745), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n202), .B1(new_n287), .B2(G41), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n724), .A2(G97), .B1(G58), .B2(new_n746), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n225), .B2(new_n732), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n1024), .A2(new_n228), .B1(new_n351), .B2(new_n743), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n736), .A2(new_n791), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n456), .B1(new_n739), .B2(new_n265), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n530), .C1(new_n516), .C2(new_n754), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT58), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1163), .A2(new_n1164), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n766), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n814), .A2(new_n202), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NOR4_X1   g0977(.A1(new_n1154), .A2(new_n714), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n985), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1153), .A2(new_n1180), .ZN(G375));
  NAND3_X1  g0981(.A1(new_n1096), .A2(new_n1093), .A3(new_n1098), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1100), .A2(new_n965), .A3(new_n1182), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n516), .A2(new_n761), .B1(new_n754), .B2(new_n576), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1025), .B(new_n1184), .C1(G107), .C2(new_n744), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n741), .A2(G97), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n530), .B1(new_n745), .B2(new_n265), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT126), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1187), .A2(KEYINPUT126), .B1(new_n756), .B2(G283), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G303), .B2(new_n737), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n741), .A2(G159), .B1(G132), .B2(new_n723), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n996), .B2(new_n732), .C1(new_n761), .C2(new_n1116), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1024), .A2(new_n202), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n292), .B1(new_n745), .B2(new_n223), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT127), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n743), .A2(new_n373), .B1(new_n1120), .B2(new_n736), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1193), .A2(new_n1194), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n766), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n713), .B(new_n1199), .C1(new_n899), .C2(new_n717), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n228), .B2(new_n814), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n985), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1183), .A2(new_n1203), .ZN(G381));
  NAND2_X1  g1004(.A1(new_n1103), .A2(new_n1125), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(G375), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G381), .A2(G384), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1073), .A2(new_n986), .A3(new_n1013), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .A4(new_n1210), .ZN(G407));
  AOI21_X1  g1011(.A(new_n649), .B1(new_n1206), .B2(new_n653), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(G407), .ZN(G409));
  NOR2_X1   g1013(.A1(new_n649), .A2(G343), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1153), .B(new_n1180), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1152), .A2(new_n965), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1178), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1147), .A2(new_n985), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1205), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1214), .B1(new_n1215), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1182), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1182), .A2(new_n1223), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n673), .A3(new_n1100), .A4(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(G384), .A3(new_n1203), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G384), .B1(new_n1226), .B2(new_n1203), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1214), .A2(G2897), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1230), .B(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT63), .B1(new_n1222), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1222), .A2(new_n1230), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G387), .A2(G390), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1208), .ZN(new_n1237));
  AND2_X1   g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(new_n1210), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1236), .B(new_n1208), .C1(new_n1210), .C2(new_n1238), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1230), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1214), .B(new_n1243), .C1(new_n1215), .C2(new_n1221), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1242), .B1(new_n1244), .B2(KEYINPUT63), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1235), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1222), .A2(new_n1248), .A3(new_n1230), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1222), .B2(new_n1232), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(new_n1222), .B2(new_n1230), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1242), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1247), .B1(new_n1252), .B2(new_n1253), .ZN(G405));
  NAND2_X1  g1054(.A1(G375), .A2(new_n1220), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1255), .A2(new_n1215), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1242), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1242), .A2(new_n1256), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1243), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1259), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1257), .A3(new_n1230), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(G402));
endmodule


