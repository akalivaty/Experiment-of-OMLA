//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT65), .B(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT66), .B(G244), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT67), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n215), .A2(KEYINPUT67), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n203), .A2(G50), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT64), .B(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n209), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT0), .Z(new_n230));
  NOR4_X1   g0030(.A1(new_n222), .A2(new_n223), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT68), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(G1698), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n254), .B1(new_n213), .B2(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT71), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n263), .A2(new_n264), .A3(new_n226), .ZN(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT71), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G226), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n206), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n276), .A2(G274), .A3(new_n271), .A4(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n270), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT74), .B(G200), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n226), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n225), .A2(G33), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n285), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n295), .A2(new_n207), .A3(G1), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n285), .ZN(new_n297));
  INV_X1    g0097(.A(G50), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n206), .B2(G20), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n297), .A2(new_n299), .B1(new_n298), .B2(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n283), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n280), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT10), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n270), .A2(new_n279), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G190), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(new_n283), .A4(new_n302), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT72), .B1(new_n307), .B2(G169), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT72), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n301), .C1(new_n316), .C2(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n253), .A2(G232), .ZN(new_n318));
  INV_X1    g0118(.A(G107), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n318), .B1(new_n319), .B2(new_n259), .C1(new_n212), .C2(new_n261), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n269), .ZN(new_n321));
  INV_X1    g0121(.A(new_n214), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n273), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n323), .A2(new_n278), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(G190), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n295), .A2(G1), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G20), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n327), .A2(KEYINPUT73), .A3(G77), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT73), .B1(new_n327), .B2(G77), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n213), .B1(new_n206), .B2(G20), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n328), .A2(new_n329), .B1(new_n297), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT15), .B(G87), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n286), .A2(new_n332), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n213), .A2(new_n225), .B1(new_n287), .B2(new_n292), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n285), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n321), .A2(new_n324), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n325), .B(new_n336), .C1(new_n338), .C2(new_n281), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n313), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n336), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AND4_X1   g0143(.A1(new_n311), .A2(new_n317), .A3(new_n339), .A4(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT75), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT64), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G20), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n346), .A2(new_n348), .A3(G33), .A4(G77), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n291), .A2(G50), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT65), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G68), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n349), .B(new_n350), .C1(new_n207), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT11), .B1(new_n355), .B2(new_n285), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n345), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n358), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT75), .A3(new_n356), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT12), .B1(new_n296), .B2(new_n202), .ZN(new_n362));
  AND4_X1   g0162(.A1(KEYINPUT12), .A2(new_n211), .A3(G20), .A4(new_n326), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n364));
  AOI211_X1 g0164(.A(new_n362), .B(new_n363), .C1(new_n297), .C2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G226), .A2(G1698), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n234), .B2(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n259), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G97), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n269), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT13), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n273), .A2(G238), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n278), .A4(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n368), .A2(new_n259), .B1(G33), .B2(G97), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n271), .A2(new_n264), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n266), .A2(KEYINPUT71), .A3(new_n267), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n374), .B(new_n278), .C1(new_n376), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT13), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n375), .A2(new_n381), .A3(G190), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n375), .B2(new_n381), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n366), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n375), .A2(new_n381), .A3(KEYINPUT77), .A4(G179), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n375), .A2(new_n381), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(new_n313), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n341), .A2(KEYINPUT76), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT14), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT14), .ZN(new_n392));
  INV_X1    g0192(.A(new_n390), .ZN(new_n393));
  AOI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(new_n375), .C2(new_n381), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n386), .B(new_n389), .C1(new_n391), .C2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n385), .B1(new_n395), .B2(new_n366), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n344), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n287), .B1(new_n206), .B2(G20), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n297), .B1(new_n296), .B2(new_n287), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n203), .B1(new_n211), .B2(new_n201), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(G20), .B1(G159), .B2(new_n291), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n252), .A2(new_n225), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n257), .A2(new_n207), .A3(new_n258), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT7), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n405), .A3(G68), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n285), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n346), .A2(new_n348), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(new_n259), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n252), .A2(new_n402), .A3(new_n207), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n354), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT16), .B1(new_n401), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n399), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n271), .A2(G232), .A3(new_n272), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  INV_X1    g0216(.A(G226), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(G1698), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n259), .B1(G33), .B2(G87), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n278), .B(new_n415), .C1(new_n419), .C2(new_n379), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G169), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n313), .B2(new_n420), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT18), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n278), .A2(new_n415), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n417), .A2(G1698), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G223), .B2(G1698), .ZN(new_n427));
  INV_X1    g0227(.A(G87), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n427), .A2(new_n252), .B1(new_n256), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n269), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT78), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n425), .A2(new_n430), .A3(new_n431), .A4(new_n304), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT78), .B1(new_n420), .B2(G190), .ZN(new_n433));
  AOI21_X1  g0233(.A(G200), .B1(new_n425), .B2(new_n430), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n399), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n407), .A2(new_n285), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT16), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n410), .A2(new_n354), .A3(new_n411), .ZN(new_n440));
  INV_X1    g0240(.A(new_n203), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n354), .B2(G58), .ZN(new_n442));
  INV_X1    g0242(.A(G159), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n442), .A2(new_n207), .B1(new_n443), .B2(new_n292), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n439), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n437), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n436), .A2(new_n446), .A3(KEYINPUT17), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n414), .A2(new_n422), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n414), .B2(new_n435), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n424), .A2(new_n447), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT25), .B1(new_n296), .B2(new_n319), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n319), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n256), .A2(G1), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n296), .A2(new_n285), .A3(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n454), .A2(new_n455), .B1(new_n457), .B2(G107), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n263), .A2(new_n226), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G1), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n463), .A2(G264), .B1(new_n465), .B2(new_n462), .ZN(new_n466));
  OAI211_X1 g0266(.A(G257), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n467));
  INV_X1    g0267(.A(G1698), .ZN(new_n468));
  OAI211_X1 g0268(.A(G250), .B(new_n468), .C1(new_n250), .C2(new_n251), .ZN(new_n469));
  INV_X1    g0269(.A(G294), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n467), .B(new_n469), .C1(new_n256), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n269), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT86), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n466), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n466), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n304), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n466), .A2(new_n472), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT87), .B1(new_n477), .B2(G200), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n466), .A2(new_n472), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT87), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(new_n383), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT85), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n259), .A2(new_n225), .A3(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT22), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n259), .A2(new_n225), .A3(new_n486), .A4(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT23), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n319), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G116), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(new_n491), .B2(new_n489), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT23), .A2(G107), .ZN(new_n493));
  AOI211_X1 g0293(.A(new_n490), .B(new_n492), .C1(new_n409), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT24), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n488), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n483), .B1(new_n499), .B2(new_n285), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n488), .A2(new_n497), .A3(new_n494), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n497), .B1(new_n488), .B2(new_n494), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n483), .B(new_n285), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n458), .B(new_n482), .C1(new_n500), .C2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n474), .A2(new_n475), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G169), .B1(G179), .B2(new_n477), .ZN(new_n507));
  INV_X1    g0307(.A(new_n458), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n285), .B1(new_n501), .B2(new_n502), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT85), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n510), .B2(new_n503), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n505), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n259), .A2(G257), .A3(new_n468), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n252), .A2(G303), .ZN(new_n514));
  INV_X1    g0314(.A(G264), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n261), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n269), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n463), .A2(G270), .B1(new_n465), .B2(new_n462), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n341), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n327), .A2(G116), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n457), .B2(G116), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  INV_X1    g0322(.A(G97), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n225), .B(new_n522), .C1(G33), .C2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G116), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n284), .A2(new_n226), .B1(G20), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(KEYINPUT20), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT20), .B1(new_n524), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT21), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n517), .A2(new_n518), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  INV_X1    g0335(.A(new_n520), .ZN(new_n536));
  OR3_X1    g0336(.A1(new_n296), .A2(new_n285), .A3(new_n456), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(new_n525), .ZN(new_n538));
  INV_X1    g0338(.A(new_n529), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(new_n527), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n517), .A2(G190), .A3(new_n518), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n535), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n534), .A2(new_n313), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n530), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n519), .A2(KEYINPUT21), .A3(new_n530), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n533), .A2(new_n542), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n457), .A2(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n296), .A2(new_n523), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n410), .A2(G107), .A3(new_n411), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT80), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(G97), .B2(new_n319), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n523), .A2(KEYINPUT80), .A3(G107), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n319), .A2(G97), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n554));
  NAND2_X1  g0354(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  OAI22_X1  g0356(.A1(new_n552), .A2(new_n553), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT79), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(new_n523), .B2(G107), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT80), .B1(new_n523), .B2(G107), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n551), .A2(new_n319), .A3(G97), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n555), .A4(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n563), .A3(new_n409), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n291), .A2(G77), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n550), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n549), .B1(new_n566), .B2(new_n285), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G244), .B(new_n468), .C1(new_n250), .C2(new_n251), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT4), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n468), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n522), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n269), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n465), .A2(new_n462), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n463), .A2(G257), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n341), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n575), .A2(new_n313), .A3(new_n576), .A4(new_n577), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n568), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(G200), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n575), .A2(G190), .A3(new_n576), .A4(new_n577), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n567), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n546), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n332), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n327), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n537), .A2(new_n428), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n346), .A2(new_n348), .A3(G33), .A4(G97), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(KEYINPUT82), .A3(new_n591), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n259), .A2(new_n225), .A3(G68), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n428), .A2(new_n523), .A3(new_n319), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n370), .A2(new_n591), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n409), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n588), .B(new_n589), .C1(new_n600), .C2(new_n285), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n212), .A2(new_n468), .ZN(new_n602));
  INV_X1    g0402(.A(G244), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G1698), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n602), .B(new_n604), .C1(new_n250), .C2(new_n251), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n491), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n269), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT81), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n459), .B2(new_n464), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n271), .A2(KEYINPUT81), .A3(G274), .A4(new_n461), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n271), .B(G250), .C1(G1), .C2(new_n460), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n607), .A2(G190), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n614));
  INV_X1    g0414(.A(G250), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n459), .A2(new_n615), .A3(new_n461), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n269), .B2(new_n606), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT83), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(G190), .A4(new_n611), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n611), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n282), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n601), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n617), .A2(new_n313), .A3(new_n611), .ZN(new_n624));
  AOI21_X1  g0424(.A(G169), .B1(new_n617), .B2(new_n611), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n600), .A2(new_n285), .ZN(new_n627));
  INV_X1    g0427(.A(new_n588), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n457), .A2(new_n587), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT84), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n623), .A2(new_n631), .A3(KEYINPUT84), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n586), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NOR4_X1   g0436(.A1(new_n397), .A2(new_n452), .A3(new_n512), .A4(new_n636), .ZN(G372));
  NAND2_X1  g0437(.A1(new_n424), .A2(new_n449), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n395), .A2(new_n366), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n385), .B2(new_n343), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n447), .A2(new_n451), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT88), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n311), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n306), .A2(KEYINPUT88), .A3(new_n310), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n317), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT89), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n397), .A2(new_n452), .ZN(new_n649));
  INV_X1    g0449(.A(new_n631), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n601), .A2(new_n622), .A3(new_n613), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n581), .A2(new_n584), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n511), .B2(new_n482), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n533), .A2(new_n544), .A3(new_n545), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n511), .B2(new_n507), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n650), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n581), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n634), .A2(KEYINPUT26), .A3(new_n635), .A4(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n651), .A2(new_n631), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n581), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n649), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n648), .A2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(KEYINPUT90), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n225), .A2(new_n326), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n511), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n666), .B1(new_n512), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n458), .B1(new_n500), .B2(new_n504), .ZN(new_n676));
  INV_X1    g0476(.A(new_n507), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n672), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT90), .A4(new_n505), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n511), .A2(new_n507), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n672), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n681), .A2(KEYINPUT91), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT91), .B1(new_n681), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n673), .A2(new_n540), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n546), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n533), .A2(new_n544), .A3(new_n545), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n688), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n686), .A2(new_n687), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT92), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n690), .A2(new_n673), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT93), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n684), .B2(new_n685), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n682), .A2(new_n673), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n700), .A3(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n228), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n206), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n597), .A2(G116), .ZN(new_n706));
  INV_X1    g0506(.A(new_n224), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n705), .A2(new_n706), .B1(new_n707), .B2(new_n704), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT28), .Z(new_n709));
  NAND3_X1  g0509(.A1(new_n634), .A2(new_n635), .A3(new_n657), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT95), .A3(new_n659), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n631), .A4(new_n651), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT95), .B1(new_n710), .B2(new_n659), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n656), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .A3(new_n673), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n672), .B1(new_n656), .B2(new_n662), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n636), .ZN(new_n720));
  INV_X1    g0520(.A(new_n512), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(new_n673), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n621), .A2(new_n479), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n575), .A2(new_n577), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n543), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n543), .A2(new_n723), .A3(new_n724), .A4(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g0528(.A(G179), .B1(new_n617), .B2(new_n611), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n578), .A2(new_n479), .A3(new_n534), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n731), .B2(new_n672), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(KEYINPUT94), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT94), .ZN(new_n736));
  INV_X1    g0536(.A(new_n734), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(new_n737), .B2(new_n732), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n722), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n719), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n709), .B1(new_n742), .B2(G1), .ZN(G364));
  AOI21_X1  g0543(.A(new_n226), .B1(G20), .B2(new_n341), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n225), .A2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(new_n313), .A3(new_n383), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT33), .B(G317), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT100), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n225), .A2(new_n313), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G190), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G200), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n748), .A2(new_n750), .B1(new_n753), .B2(G322), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT101), .Z(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n259), .B1(new_n758), .B2(G329), .ZN(new_n759));
  INV_X1    g0559(.A(G311), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n751), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n752), .A2(new_n383), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(G326), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n281), .A2(G179), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n207), .A2(new_n304), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT99), .Z(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G303), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n746), .A2(new_n766), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT96), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n409), .B1(new_n304), .B2(new_n757), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT98), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G283), .A2(new_n772), .B1(new_n778), .B2(G294), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n755), .A2(new_n765), .A3(new_n770), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n772), .A2(G107), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n781), .B(new_n259), .C1(new_n428), .C2(new_n768), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  INV_X1    g0583(.A(new_n758), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n443), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT32), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n764), .ZN(new_n788));
  INV_X1    g0588(.A(new_n753), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n787), .B1(new_n298), .B2(new_n788), .C1(new_n201), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n778), .A2(G97), .ZN(new_n791));
  INV_X1    g0591(.A(new_n762), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n748), .A2(G68), .B1(G77), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n791), .B(new_n793), .C1(new_n786), .C2(new_n785), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n780), .B1(new_n783), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n745), .B1(new_n796), .B2(KEYINPUT102), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(KEYINPUT102), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n693), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n409), .A2(new_n295), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G45), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n705), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n245), .A2(G45), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n703), .A2(new_n259), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G45), .C2(new_n224), .ZN(new_n808));
  INV_X1    g0608(.A(G355), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n228), .A2(new_n259), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(G116), .B2(new_n228), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n801), .A2(new_n744), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n798), .A2(new_n802), .A3(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT103), .Z(new_n815));
  OAI21_X1  g0615(.A(new_n805), .B1(new_n693), .B2(new_n687), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n687), .B2(new_n693), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  INV_X1    g0619(.A(new_n805), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n673), .A2(new_n336), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n339), .A2(new_n821), .B1(new_n340), .B2(new_n342), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n340), .A2(new_n342), .A3(new_n673), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n717), .B(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n820), .B1(new_n826), .B2(new_n740), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n740), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n744), .A2(new_n799), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n820), .B1(G77), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G303), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n470), .A2(new_n789), .B1(new_n788), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n748), .ZN(new_n834));
  INV_X1    g0634(.A(G283), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n252), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n784), .A2(new_n760), .B1(new_n525), .B2(new_n762), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n772), .A2(G87), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n769), .A2(G107), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n838), .A2(new_n791), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n772), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n202), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G50), .B2(new_n769), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n259), .B1(new_n784), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n778), .B2(G58), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT34), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n748), .A2(G150), .B1(G159), .B2(new_n792), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n764), .A2(G137), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n753), .A2(G143), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n844), .B(new_n847), .C1(new_n848), .C2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n852), .A2(new_n848), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n841), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n831), .B1(new_n855), .B2(new_n744), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n800), .B2(new_n825), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n828), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G384));
  NOR2_X1   g0659(.A1(new_n803), .A2(new_n206), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT40), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n366), .A2(new_n672), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n862), .B(new_n385), .C1(new_n395), .C2(new_n366), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n395), .A2(new_n862), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n825), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n737), .A2(new_n732), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(new_n722), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n670), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n414), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n445), .A2(new_n285), .A3(new_n407), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n420), .A2(new_n383), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n425), .A2(new_n304), .A3(new_n430), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT78), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(new_n399), .A3(new_n432), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n423), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n423), .A2(new_n870), .A3(new_n875), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(KEYINPUT105), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n870), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n452), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT105), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n876), .A2(new_n883), .A3(KEYINPUT37), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT16), .B1(new_n401), .B2(new_n406), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n399), .B1(new_n408), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n869), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n452), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(new_n422), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n893), .A2(new_n890), .A3(new_n875), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n879), .B1(new_n894), .B2(new_n878), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n887), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n861), .B1(new_n868), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n892), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n892), .B2(new_n895), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n861), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n325), .A2(new_n336), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n281), .B1(new_n321), .B2(new_n324), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n821), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n343), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n823), .ZN(new_n906));
  INV_X1    g0706(.A(new_n862), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n396), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n908), .B2(new_n864), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n636), .A2(new_n512), .A3(new_n672), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n733), .A2(new_n734), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n898), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n722), .A2(new_n867), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n649), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n916), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(G330), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT106), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n716), .A2(new_n649), .A3(new_n718), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n648), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n639), .A2(new_n672), .ZN(new_n923));
  INV_X1    g0723(.A(new_n900), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n899), .B1(new_n886), .B2(new_n885), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n923), .B(new_n925), .C1(new_n926), .C2(KEYINPUT39), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n863), .A2(new_n865), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n896), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n672), .B(new_n906), .C1(new_n656), .C2(new_n662), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n824), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n638), .A2(new_n670), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n927), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n922), .B(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n860), .B1(new_n920), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n920), .B2(new_n935), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n225), .A2(new_n525), .A3(new_n226), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n557), .A2(new_n563), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT35), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n939), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT36), .Z(new_n943));
  AOI211_X1 g0743(.A(new_n213), .B(new_n224), .C1(new_n354), .C2(G58), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT104), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n944), .A2(new_n945), .B1(new_n298), .B2(G68), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(G1), .A3(new_n295), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n937), .A2(new_n943), .A3(new_n948), .ZN(G367));
  INV_X1    g0749(.A(new_n768), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT46), .B1(new_n950), .B2(G116), .ZN(new_n951));
  INV_X1    g0751(.A(new_n769), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n952), .A2(new_n953), .A3(new_n525), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n951), .B(new_n954), .C1(G294), .C2(new_n748), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT110), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT110), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n832), .A2(new_n789), .B1(new_n788), .B2(new_n760), .ZN(new_n958));
  INV_X1    g0758(.A(new_n771), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G97), .A2(new_n959), .B1(new_n792), .B2(G283), .ZN(new_n960));
  INV_X1    g0760(.A(G317), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n252), .C1(new_n961), .C2(new_n784), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n958), .B(new_n962), .C1(G107), .C2(new_n778), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n956), .A2(new_n957), .A3(new_n963), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n298), .A2(new_n762), .B1(new_n768), .B2(new_n201), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT111), .B(G137), .Z(new_n966));
  OAI22_X1  g0766(.A1(new_n784), .A2(new_n966), .B1(new_n213), .B2(new_n771), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n965), .B(new_n967), .C1(G68), .C2(new_n778), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n259), .B1(new_n834), .B2(new_n443), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G143), .B2(new_n764), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n968), .B(new_n970), .C1(new_n290), .C2(new_n789), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT47), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n744), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n601), .A2(new_n673), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n660), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n650), .A2(new_n975), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n801), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n807), .A2(new_n240), .ZN(new_n979));
  INV_X1    g0779(.A(new_n812), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n703), .B2(new_n587), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n805), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n974), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n657), .A2(new_n672), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n581), .B(new_n584), .C1(new_n567), .C2(new_n673), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n700), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n581), .B1(new_n678), .B2(new_n985), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n988), .A2(KEYINPUT42), .B1(new_n673), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT108), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT108), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n976), .A2(new_n977), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT107), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n993), .A2(new_n995), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1000), .B1(KEYINPUT43), .B2(new_n996), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n993), .B2(new_n995), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1002), .A2(new_n1005), .B1(new_n696), .B2(new_n987), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1005), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n696), .A2(new_n987), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n1008), .A3(new_n1001), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n804), .A2(G1), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n700), .A2(new_n701), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n987), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n701), .A4(new_n986), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT44), .B1(new_n1013), .B2(new_n987), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1013), .A2(KEYINPUT44), .A3(new_n987), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n694), .B(KEYINPUT92), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n696), .B(new_n1016), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n686), .A2(new_n698), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n700), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n693), .A2(new_n687), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(KEYINPUT109), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1025), .B(KEYINPUT109), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n1023), .B2(new_n700), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1021), .A2(new_n1022), .A3(new_n742), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n742), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n704), .B(KEYINPUT41), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1011), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n983), .B1(new_n1010), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT112), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(G387));
  NAND2_X1  g0838(.A1(new_n1030), .A2(new_n742), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n741), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n704), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n686), .A2(new_n801), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n810), .A2(new_n706), .B1(G107), .B2(new_n228), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n237), .A2(new_n460), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n706), .ZN(new_n1045));
  AOI211_X1 g0845(.A(G45), .B(new_n1045), .C1(G68), .C2(G77), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n287), .A2(G50), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT50), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n703), .B(new_n259), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1043), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n820), .B1(new_n1050), .B2(new_n980), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n950), .A2(G77), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n259), .B(new_n1052), .C1(new_n789), .C2(new_n298), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G159), .B2(new_n764), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n772), .A2(G97), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n778), .A2(new_n587), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n784), .A2(new_n290), .B1(new_n202), .B2(new_n762), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n287), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n748), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n748), .A2(G311), .B1(G303), .B2(new_n792), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n764), .A2(G322), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n961), .C2(new_n789), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n778), .A2(G283), .B1(G294), .B2(new_n950), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT49), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n259), .B1(new_n758), .B2(G326), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n525), .C2(new_n771), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1060), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1051), .B1(new_n1074), .B2(new_n744), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1030), .A2(new_n1011), .B1(new_n1042), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1041), .A2(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(KEYINPUT114), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1021), .A2(new_n1022), .A3(new_n1078), .ZN(new_n1079));
  OR3_X1    g0879(.A1(new_n1019), .A2(new_n1078), .A3(new_n1020), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT115), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT115), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n1011), .A3(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1031), .A2(new_n704), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1079), .A2(new_n1080), .A3(new_n1039), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n987), .A2(new_n801), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n812), .B1(new_n523), .B2(new_n228), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n807), .B2(new_n248), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G311), .A2(new_n753), .B1(new_n764), .B2(G317), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n834), .A2(new_n832), .B1(new_n835), .B2(new_n768), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G322), .B2(new_n758), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n259), .B1(new_n792), .B2(G294), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n778), .A2(G116), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1093), .A2(new_n781), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n834), .A2(new_n298), .B1(new_n211), .B2(new_n768), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G143), .B2(new_n758), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n252), .B1(new_n792), .B2(new_n1058), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n777), .A2(new_n213), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n839), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G150), .A2(new_n764), .B1(new_n753), .B2(G159), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT51), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1091), .A2(new_n1096), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n805), .B(new_n1089), .C1(new_n1105), .C2(new_n744), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1085), .A2(new_n1086), .B1(new_n1087), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1084), .A2(new_n1107), .ZN(G390));
  AOI22_X1  g0908(.A1(G128), .A2(new_n764), .B1(new_n753), .B2(G132), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n950), .A2(G150), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(KEYINPUT53), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(KEYINPUT53), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1112), .B1(new_n762), .B2(new_n1113), .C1(new_n834), .C2(new_n966), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1111), .B(new_n1114), .C1(G159), .C2(new_n778), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n259), .B1(new_n771), .B2(new_n298), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G125), .B2(new_n758), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT117), .Z(new_n1118));
  AOI211_X1 g0918(.A(new_n1100), .B(new_n843), .C1(G87), .C2(new_n769), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n525), .A2(new_n789), .B1(new_n788), .B2(new_n835), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n252), .B1(new_n834), .B2(new_n319), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n784), .A2(new_n470), .B1(new_n523), .B2(new_n762), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1115), .A2(new_n1118), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n820), .B1(new_n1058), .B2(new_n830), .C1(new_n1124), .C2(new_n745), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT118), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n925), .B1(new_n926), .B2(KEYINPUT39), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n799), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n658), .A2(new_n661), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n690), .B1(new_n676), .B2(new_n677), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n581), .A2(new_n584), .A3(new_n651), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n505), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n631), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n673), .B(new_n825), .C1(new_n1129), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n928), .B1(new_n1134), .B2(new_n823), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT39), .B1(new_n887), .B2(new_n896), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1135), .A2(new_n923), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n715), .A2(new_n673), .A3(new_n905), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n928), .B1(new_n1139), .B2(new_n823), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n926), .A2(new_n923), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1138), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT116), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n687), .B1(new_n722), .B2(new_n867), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n909), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1143), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n739), .A2(G330), .A3(new_n825), .A4(new_n929), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1138), .B(new_n1149), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1144), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1148), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1128), .B1(new_n1153), .B2(new_n1011), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1145), .A2(new_n825), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1149), .B1(new_n1155), .B2(new_n929), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1139), .A2(new_n823), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n739), .A2(G330), .A3(new_n825), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1158), .A2(new_n928), .B1(new_n1145), .B2(new_n909), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n824), .B1(new_n717), .B2(new_n825), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1156), .A2(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n649), .A2(new_n1145), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n648), .A2(new_n921), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n704), .B1(new_n1153), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT95), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n623), .A2(KEYINPUT84), .A3(new_n631), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT84), .B1(new_n623), .B2(new_n631), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1169), .A2(new_n1170), .A3(new_n581), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1168), .B1(new_n1171), .B2(KEYINPUT26), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(new_n712), .A3(new_n711), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n672), .B(new_n822), .C1(new_n1173), .C2(new_n656), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n929), .B1(new_n1174), .B2(new_n824), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1160), .A2(new_n928), .B1(new_n639), .B2(new_n672), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1175), .A2(new_n1141), .B1(new_n1127), .B2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(KEYINPUT116), .B(new_n1150), .C1(new_n1177), .C2(new_n1146), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1143), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1165), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1154), .B1(new_n1167), .B2(new_n1180), .ZN(G378));
  INV_X1    g0981(.A(G41), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1052), .A2(new_n1182), .A3(new_n252), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1183), .A2(KEYINPUT119), .B1(new_n778), .B2(G68), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(KEYINPUT119), .B2(new_n1183), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G283), .A2(new_n758), .B1(new_n792), .B2(new_n587), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n959), .A2(G58), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n523), .C2(new_n834), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n319), .A2(new_n789), .B1(new_n788), .B2(new_n525), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1185), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n252), .A2(new_n1182), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G50), .B1(new_n256), .B2(new_n1182), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1190), .A2(KEYINPUT58), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n834), .A2(new_n845), .B1(new_n768), .B2(new_n1113), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G137), .B2(new_n792), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G125), .A2(new_n764), .B1(new_n753), .B2(G128), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n290), .C2(new_n777), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n256), .B(new_n1182), .C1(new_n771), .C2(new_n443), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G124), .B2(new_n758), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1193), .B1(KEYINPUT58), .B2(new_n1190), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n744), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n805), .B1(new_n298), .B2(new_n829), .ZN(new_n1205));
  XOR2_X1   g1005(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1206));
  INV_X1    g1006(.A(KEYINPUT120), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n306), .A2(KEYINPUT88), .A3(new_n310), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT88), .B1(new_n306), .B2(new_n310), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1207), .B1(new_n1210), .B2(new_n317), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n1207), .A2(new_n644), .A3(new_n317), .A4(new_n645), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1206), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n869), .A2(new_n301), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n317), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT120), .B1(new_n646), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1210), .A2(new_n1207), .A3(new_n317), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1206), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1213), .A2(new_n1215), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1215), .B1(new_n1213), .B2(new_n1220), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1204), .B(new_n1205), .C1(new_n1223), .C2(new_n800), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(G330), .B1(new_n898), .B2(new_n913), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1135), .A2(new_n930), .B1(new_n638), .B2(new_n670), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n927), .A3(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT40), .B1(new_n926), .B2(new_n912), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n868), .A2(new_n861), .A3(new_n930), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n687), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n934), .A2(new_n1231), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1228), .A2(new_n1232), .A3(new_n1223), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1223), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1225), .B1(new_n1235), .B2(new_n1011), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1164), .B1(new_n1152), .B2(new_n1165), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1237), .B2(new_n1235), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n704), .B1(new_n1238), .B2(KEYINPUT122), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1235), .B1(new_n1180), .B2(new_n1163), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(KEYINPUT122), .A3(new_n1241), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1233), .A2(new_n1234), .A3(new_n1241), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT121), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(KEYINPUT121), .C1(new_n1180), .C2(new_n1163), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1242), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1236), .B1(new_n1239), .B2(new_n1247), .ZN(G375));
  NAND2_X1  g1048(.A1(new_n1187), .A2(new_n259), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT125), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n952), .A2(new_n443), .B1(new_n298), .B2(new_n777), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G128), .A2(new_n758), .B1(new_n792), .B2(G150), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n834), .B2(new_n1113), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n845), .A2(new_n788), .B1(new_n789), .B2(new_n966), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n748), .A2(G116), .B1(G107), .B2(new_n792), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n470), .B2(new_n788), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT124), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n952), .A2(new_n523), .B1(new_n842), .B2(new_n213), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n259), .B1(new_n758), .B2(G303), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1056), .B(new_n1260), .C1(new_n835), .C2(new_n789), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1250), .A2(new_n1255), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n820), .B1(G68), .B2(new_n830), .C1(new_n1263), .C2(new_n745), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n928), .B2(new_n799), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1011), .B(KEYINPUT123), .Z(new_n1266));
  AOI21_X1  g1066(.A(new_n1265), .B1(new_n1161), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1165), .A2(new_n1034), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1268), .B2(new_n1269), .ZN(G381));
  INV_X1    g1070(.A(G378), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1236), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1243), .B1(new_n1180), .B2(new_n1163), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT121), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1238), .A2(KEYINPUT122), .B1(new_n1275), .B2(new_n1245), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n704), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT122), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1272), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n858), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(G390), .A2(G381), .A3(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1037), .A2(new_n1271), .A3(new_n1281), .A4(new_n1284), .ZN(G407));
  NAND2_X1  g1085(.A1(new_n671), .A2(G213), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1281), .A2(new_n1271), .A3(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G407), .A2(G213), .A3(new_n1288), .ZN(G409));
  INV_X1    g1089(.A(new_n1036), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT112), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n818), .B1(new_n1041), .B2(new_n1076), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1282), .B2(new_n1292), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1084), .A2(new_n1107), .A3(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1282), .A2(new_n1292), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1084), .B2(new_n1107), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1290), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1282), .A2(new_n1292), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G390), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1084), .A2(new_n1107), .A3(new_n1293), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1300), .A3(new_n1036), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G378), .B(new_n1236), .C1(new_n1239), .C2(new_n1247), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1237), .A2(new_n1034), .A3(new_n1235), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1225), .B1(new_n1235), .B2(new_n1266), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G378), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1165), .A2(KEYINPUT60), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n1269), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1165), .A2(KEYINPUT60), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1312), .B(KEYINPUT126), .C1(new_n1164), .C2(new_n1161), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1277), .B1(new_n1269), .B2(KEYINPUT60), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1311), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(G384), .A3(new_n1267), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G384), .B1(new_n1315), .B2(new_n1267), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1308), .A2(new_n1286), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT62), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1287), .B1(new_n1303), .B2(new_n1307), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(new_n1323), .A3(new_n1319), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1287), .A2(G2897), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1318), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(new_n1316), .A3(new_n1326), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1306), .B1(new_n1281), .B2(G378), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1331), .B1(new_n1332), .B2(new_n1287), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT61), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT127), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1302), .B1(new_n1325), .B2(new_n1335), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1337));
  AND4_X1   g1137(.A1(KEYINPUT63), .A2(new_n1308), .A3(new_n1286), .A4(new_n1319), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT63), .B1(new_n1322), .B2(new_n1319), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1337), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT127), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1334), .B1(new_n1322), .B2(new_n1342), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1340), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1336), .A2(new_n1345), .ZN(G405));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1271), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1303), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1348), .A2(new_n1319), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1319), .ZN(new_n1350));
  OR3_X1    g1150(.A1(new_n1349), .A2(new_n1350), .A3(new_n1302), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1302), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(G402));
endmodule


