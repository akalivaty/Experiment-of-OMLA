//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(G64gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G92gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G211gat), .B(G218gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n207), .A3(new_n211), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  AND2_X1   g028(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n230));
  NOR2_X1   g029(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n228), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(KEYINPUT23), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n237), .A2(KEYINPUT23), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n219), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT64), .B(G169gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(G176gat), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n239), .B1(new_n246), .B2(KEYINPUT23), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(new_n227), .A3(new_n220), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n241), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n222), .A2(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n234), .B1(new_n254), .B2(new_n229), .ZN(new_n255));
  INV_X1    g054(.A(new_n235), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(KEYINPUT68), .A3(new_n242), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(new_n252), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n237), .ZN(new_n260));
  OR3_X1    g059(.A1(new_n260), .A2(KEYINPUT70), .A3(KEYINPUT26), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(KEYINPUT26), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n260), .A2(KEYINPUT26), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT70), .B1(G169gat), .B2(G176gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n261), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT27), .B(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n266), .A2(new_n226), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n226), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(new_n267), .A3(KEYINPUT28), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n265), .A2(new_n270), .A3(new_n229), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n259), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G226gat), .A2(G233gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT79), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n277), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n259), .A2(KEYINPUT78), .A3(new_n273), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT78), .B1(new_n259), .B2(new_n273), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(KEYINPUT79), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n218), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n275), .B(new_n277), .C1(new_n280), .C2(new_n281), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n274), .A2(new_n277), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n218), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n206), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT78), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n257), .A2(KEYINPUT68), .A3(new_n242), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT68), .B1(new_n257), .B2(new_n242), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT25), .B1(new_n247), .B2(new_n250), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n273), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n259), .A2(KEYINPUT78), .A3(new_n273), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n277), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT79), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n259), .B2(new_n273), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(new_n279), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n284), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n217), .ZN(new_n305));
  INV_X1    g104(.A(new_n206), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n289), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n291), .A2(KEYINPUT30), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT40), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT39), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G120gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT72), .B(G120gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(new_n311), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n315));
  XOR2_X1   g114(.A(G127gat), .B(G134gat), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT73), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G113gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n322), .A2(KEYINPUT71), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n315), .B1(new_n322), .B2(KEYINPUT71), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n316), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n314), .A2(new_n317), .A3(new_n326), .A4(new_n315), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G155gat), .B(G162gat), .Z(new_n329));
  AND2_X1   g128(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G148gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT80), .B1(new_n334), .B2(G141gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336));
  INV_X1    g135(.A(G141gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(G148gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n335), .B(new_n338), .C1(new_n337), .C2(G148gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n334), .A2(G141gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n337), .A2(G148gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n331), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n333), .A2(new_n339), .B1(new_n342), .B2(new_n329), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n319), .A2(new_n325), .A3(new_n343), .A4(new_n327), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT83), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n346), .B(KEYINPUT4), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n328), .B(new_n352), .C1(new_n344), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  AOI211_X1 g154(.A(new_n310), .B(new_n350), .C1(new_n355), .C2(new_n349), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n310), .A3(new_n349), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G85gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n309), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n350), .B1(new_n355), .B2(new_n349), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT39), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n365), .A2(KEYINPUT40), .A3(new_n361), .A4(new_n357), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n347), .B2(new_n349), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n346), .A2(new_n349), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n355), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n354), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n361), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n363), .A2(new_n366), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n305), .A2(new_n377), .A3(new_n289), .A4(new_n306), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n308), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n380), .B(G22gat), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n353), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n343), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(new_n217), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT29), .B1(new_n215), .B2(new_n216), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n344), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n386), .A2(new_n387), .A3(new_n352), .A4(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(new_n352), .C1(new_n217), .C2(new_n384), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT85), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT31), .B(G50gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n353), .B1(new_n389), .B2(new_n397), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n343), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n388), .B1(new_n400), .B2(new_n385), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n394), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n396), .B1(new_n394), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n382), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n394), .A2(new_n401), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n395), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n381), .A3(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n379), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT37), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n305), .A2(new_n413), .A3(new_n289), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT87), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n305), .A2(new_n416), .A3(new_n413), .A4(new_n289), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n298), .B2(new_n299), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n287), .B1(new_n419), .B2(new_n277), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT86), .B1(new_n420), .B2(new_n218), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n283), .A2(new_n218), .A3(new_n284), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n286), .A2(new_n288), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n217), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT38), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n418), .A2(new_n427), .A3(new_n206), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n370), .A2(new_n372), .A3(new_n361), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n375), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n373), .A2(KEYINPUT6), .A3(new_n374), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n307), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT38), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n306), .B1(new_n415), .B2(new_n417), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT37), .B1(new_n285), .B2(new_n290), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n412), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT76), .ZN(new_n441));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(G71gat), .ZN(new_n443));
  INV_X1    g242(.A(G99gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(KEYINPUT74), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT33), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n328), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n259), .A2(new_n449), .A3(new_n273), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n259), .B2(new_n273), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G227gat), .ZN(new_n453));
  INV_X1    g252(.A(G233gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT32), .B(new_n448), .C1(new_n452), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n274), .A2(new_n328), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n259), .A2(new_n449), .A3(new_n273), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n460), .A2(new_n455), .B1(new_n461), .B2(KEYINPUT33), .ZN(new_n462));
  INV_X1    g261(.A(new_n445), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT34), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n460), .B2(new_n455), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n452), .A2(KEYINPUT34), .A3(new_n456), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n441), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n470));
  OAI22_X1  g269(.A1(new_n452), .A2(new_n456), .B1(KEYINPUT32), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n445), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n466), .A2(new_n467), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT76), .A4(new_n457), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n472), .B2(new_n457), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT75), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n464), .A2(new_n468), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT75), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n478), .A3(KEYINPUT36), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(new_n479), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n308), .A2(new_n378), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n431), .A2(new_n432), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n481), .A2(new_n484), .B1(new_n487), .B2(new_n409), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n475), .A2(new_n410), .A3(new_n480), .A4(new_n478), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT35), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n475), .A2(new_n410), .A3(new_n479), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT35), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n486), .A4(new_n485), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n440), .A2(new_n488), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n495), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(KEYINPUT16), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(G1gat), .B1(new_n495), .B2(KEYINPUT91), .ZN(new_n499));
  OAI21_X1  g298(.A(G8gat), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n497), .A2(KEYINPUT16), .ZN(new_n501));
  INV_X1    g300(.A(new_n499), .ZN(new_n502));
  INV_X1    g301(.A(G8gat), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n496), .ZN(new_n504));
  NOR2_X1   g303(.A1(G29gat), .A2(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT14), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n509));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n506), .A2(new_n508), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G50gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G43gat), .ZN(new_n513));
  INV_X1    g312(.A(G43gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G50gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT15), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n511), .A2(new_n516), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n506), .A2(new_n508), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n512), .B2(G43gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n513), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n520), .A2(new_n524), .A3(new_n525), .A4(new_n510), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT17), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n511), .A2(new_n516), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n516), .ZN(new_n529));
  AND4_X1   g328(.A1(KEYINPUT17), .A2(new_n528), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n500), .B(new_n504), .C1(new_n527), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n519), .A2(new_n526), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n500), .A2(new_n504), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n500), .A3(new_n504), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n540), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT92), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n532), .B(KEYINPUT13), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n532), .A4(new_n536), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n539), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT11), .B(G169gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XOR2_X1   g349(.A(G113gat), .B(G141gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT12), .A3(new_n553), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n547), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n559), .A2(new_n539), .A3(new_n545), .A4(new_n546), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n494), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567));
  INV_X1    g366(.A(G57gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n567), .B(G64gat), .C1(new_n568), .C2(KEYINPUT94), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT93), .B1(new_n203), .B2(G57gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n203), .A2(G57gat), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n569), .B(new_n570), .C1(KEYINPUT94), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  INV_X1    g372(.A(G71gat), .ZN(new_n574));
  INV_X1    g373(.A(G78gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n572), .A2(KEYINPUT95), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n572), .A2(new_n578), .A3(new_n576), .ZN(new_n579));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n566), .A2(new_n580), .A3(new_n573), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n566), .A2(new_n577), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n584), .A2(KEYINPUT96), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(KEYINPUT96), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT97), .B(G211gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n587), .ZN(new_n589));
  INV_X1    g388(.A(new_n586), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n584), .A2(KEYINPUT96), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n566), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n579), .A2(new_n581), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n535), .B1(KEYINPUT21), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n225), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n582), .A2(new_n583), .ZN(new_n598));
  OAI21_X1  g397(.A(G183gat), .B1(new_n598), .B2(new_n535), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(new_n597), .B2(new_n599), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n588), .B(new_n592), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n592), .A2(new_n588), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n597), .A2(new_n599), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n604), .A2(new_n609), .A3(new_n613), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G134gat), .B(G162gat), .Z(new_n618));
  NAND2_X1  g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT102), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G106gat), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT98), .B1(new_n444), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(G99gat), .A3(G106gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(KEYINPUT8), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G85gat), .A2(G92gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT7), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT99), .B(G85gat), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n629), .B(new_n631), .C1(G92gat), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G99gat), .B(G106gat), .Z(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n205), .ZN(new_n637));
  INV_X1    g436(.A(new_n634), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n629), .A4(new_n631), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n527), .B2(new_n530), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n642));
  OAI22_X1  g441(.A1(new_n533), .A2(new_n640), .B1(new_n620), .B2(new_n619), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI221_X1 g444(.A(KEYINPUT101), .B1(new_n620), .B2(new_n619), .C1(new_n533), .C2(new_n640), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n642), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n642), .A2(new_n647), .A3(new_n652), .A4(new_n648), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n624), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n622), .A2(KEYINPUT102), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n651), .A2(new_n656), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n617), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT104), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G120gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n635), .A2(new_n639), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n595), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n582), .A2(new_n640), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n665), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n663), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT106), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(new_n677), .B2(new_n664), .ZN(new_n678));
  INV_X1    g477(.A(new_n663), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR4_X1   g479(.A1(new_n672), .A2(KEYINPUT105), .A3(new_n673), .A4(new_n663), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n659), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n565), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n486), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G1gat), .ZN(G1324gat));
  INV_X1    g489(.A(new_n485), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT16), .B(G8gat), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT107), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(G8gat), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697));
  OAI211_X1 g496(.A(KEYINPUT107), .B(new_n697), .C1(new_n692), .C2(new_n693), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(G1325gat));
  NAND2_X1  g498(.A1(new_n484), .A2(new_n481), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n687), .A2(G15gat), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n482), .ZN(new_n703));
  AOI21_X1  g502(.A(G15gat), .B1(new_n687), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n686), .A2(new_n410), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  NOR3_X1   g507(.A1(new_n684), .A2(new_n617), .A3(new_n658), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n565), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(G29gat), .A3(new_n486), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n490), .A2(new_n493), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n418), .A2(new_n206), .A3(new_n438), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT38), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n433), .B1(new_n437), .B2(new_n427), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n411), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n487), .A2(new_n409), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n700), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n716), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n657), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n654), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(KEYINPUT44), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT44), .B1(new_n723), .B2(new_n725), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n604), .A2(new_n609), .A3(new_n613), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n613), .B1(new_n604), .B2(new_n609), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n615), .A2(KEYINPUT109), .A3(new_n616), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(new_n564), .A3(new_n684), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n729), .A2(new_n688), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G29gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n715), .A2(new_n738), .ZN(G1328gat));
  NOR3_X1   g538(.A1(new_n712), .A2(G36gat), .A3(new_n485), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n729), .A2(new_n691), .A3(new_n736), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G36gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(G1329gat));
  NAND2_X1  g545(.A1(new_n723), .A2(new_n725), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n749), .A2(new_n701), .A3(new_n726), .A4(new_n736), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G43gat), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT47), .B1(new_n751), .B2(KEYINPUT110), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n565), .A2(new_n710), .A3(new_n711), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n514), .A3(new_n703), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n751), .B(new_n754), .C1(KEYINPUT110), .C2(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1330gat));
  NAND4_X1  g557(.A1(new_n749), .A2(new_n409), .A3(new_n726), .A4(new_n736), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G50gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n753), .A2(new_n512), .A3(new_n409), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1331gat));
  NOR2_X1   g563(.A1(new_n683), .A2(new_n563), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n617), .A3(new_n658), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT111), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT112), .B1(new_n494), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  INV_X1    g568(.A(new_n767), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n723), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n486), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n568), .ZN(G1332gat));
  NOR2_X1   g573(.A1(new_n772), .A2(new_n485), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT49), .B(G64gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n775), .B2(new_n778), .ZN(G1333gat));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n768), .A2(new_n703), .A3(new_n771), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n574), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n771), .A3(G71gat), .A4(new_n701), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n780), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(KEYINPUT50), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(G1334gat));
  NOR2_X1   g591(.A1(new_n772), .A2(new_n410), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(new_n575), .ZN(G1335gat));
  INV_X1    g593(.A(new_n617), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n765), .A2(new_n795), .ZN(new_n796));
  NOR4_X1   g595(.A1(new_n727), .A2(new_n728), .A3(new_n636), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n617), .A2(new_n563), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT51), .B1(new_n747), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n723), .A2(new_n801), .A3(new_n725), .A4(new_n798), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n800), .A2(new_n688), .A3(new_n684), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n797), .A2(new_n688), .B1(new_n803), .B2(new_n636), .ZN(G1336gat));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805));
  INV_X1    g604(.A(new_n796), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n729), .A2(new_n805), .A3(new_n691), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n749), .A2(new_n691), .A3(new_n726), .A4(new_n806), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n807), .A2(G92gat), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n485), .A2(G92gat), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n800), .A2(new_n684), .A3(new_n802), .A4(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(G92gat), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n812), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n810), .A2(new_n814), .B1(new_n816), .B2(new_n813), .ZN(G1337gat));
  NOR4_X1   g616(.A1(new_n727), .A2(new_n728), .A3(new_n700), .A4(new_n796), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n800), .A2(new_n444), .A3(new_n684), .A4(new_n802), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n818), .A2(new_n444), .B1(new_n819), .B2(new_n482), .ZN(G1338gat));
  NOR2_X1   g619(.A1(new_n410), .A2(G106gat), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n800), .A2(new_n684), .A3(new_n802), .A4(new_n821), .ZN(new_n822));
  NOR4_X1   g621(.A1(new_n727), .A2(new_n728), .A3(new_n410), .A4(new_n796), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n625), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g624(.A1(new_n733), .A2(new_n734), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n544), .B1(new_n541), .B2(new_n542), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n532), .B1(new_n531), .B2(new_n536), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n552), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n562), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n675), .B2(new_n682), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n677), .A2(new_n664), .ZN(new_n832));
  INV_X1    g631(.A(new_n673), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n833), .A3(new_n679), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT105), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n678), .A2(new_n676), .A3(new_n679), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n670), .A2(new_n665), .A3(new_n671), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT54), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n672), .ZN(new_n841));
  XOR2_X1   g640(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n677), .A2(new_n664), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n663), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n838), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n679), .B1(new_n672), .B2(new_n842), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n846), .B(KEYINPUT55), .C1(new_n672), .C2(new_n840), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n837), .A2(new_n563), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n725), .B1(new_n831), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n837), .A2(new_n830), .A3(new_n845), .A4(new_n847), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n658), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n826), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n617), .A2(new_n683), .A3(new_n658), .A4(new_n564), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(KEYINPUT116), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n485), .A2(new_n688), .ZN(new_n859));
  NOR4_X1   g658(.A1(new_n858), .A2(new_n409), .A3(new_n482), .A4(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n564), .ZN(new_n862));
  INV_X1    g661(.A(new_n489), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n856), .A2(new_n688), .A3(new_n863), .A4(new_n857), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT117), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n485), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n563), .A2(new_n311), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT119), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n862), .B1(new_n868), .B2(new_n870), .ZN(G1340gat));
  OAI21_X1  g670(.A(G120gat), .B1(new_n861), .B2(new_n683), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n683), .A2(new_n313), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n868), .B2(new_n873), .ZN(G1341gat));
  INV_X1    g673(.A(G127gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n861), .A2(new_n875), .A3(new_n826), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n865), .A2(new_n485), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n617), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(new_n875), .ZN(G1342gat));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n658), .A2(G134gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n877), .A2(new_n881), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT56), .ZN(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n861), .B2(new_n658), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n877), .A2(new_n887), .A3(new_n880), .A4(new_n881), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n883), .A2(new_n885), .A3(new_n886), .A4(new_n888), .ZN(G1343gat));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n852), .A2(KEYINPUT116), .A3(new_n853), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT116), .B1(new_n852), .B2(new_n853), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n891), .A2(new_n892), .A3(new_n410), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n890), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT121), .B(new_n895), .C1(new_n858), .C2(new_n410), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n831), .A2(new_n848), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n658), .ZN(new_n898));
  INV_X1    g697(.A(new_n851), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n617), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n853), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT57), .B(new_n409), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n894), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n701), .A2(new_n859), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n563), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G141gat), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n893), .A2(new_n904), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n337), .A3(new_n563), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT58), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1344gat));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n903), .A2(new_n904), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n914), .B(G148gat), .C1(new_n915), .C2(new_n683), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n898), .A2(new_n899), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT123), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n853), .B1(new_n918), .B2(new_n617), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n895), .A3(new_n409), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT57), .B1(new_n858), .B2(new_n410), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n920), .A2(new_n684), .A3(new_n904), .A4(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(G148gat), .ZN(new_n923));
  XOR2_X1   g722(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n924));
  OAI21_X1  g723(.A(new_n916), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n334), .A3(new_n684), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1345gat));
  AOI21_X1  g726(.A(G155gat), .B1(new_n907), .B2(new_n617), .ZN(new_n928));
  INV_X1    g727(.A(new_n915), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n735), .A2(G155gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G1346gat));
  NOR2_X1   g730(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n330), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n907), .A2(new_n725), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT124), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n915), .A2(new_n658), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n933), .B2(new_n936), .ZN(G1347gat));
  INV_X1    g736(.A(new_n858), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n485), .A2(new_n688), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n491), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n564), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n858), .A2(new_n489), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n939), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n564), .A2(new_n245), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1348gat));
  INV_X1    g744(.A(G176gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n940), .A2(new_n946), .A3(new_n683), .ZN(new_n947));
  INV_X1    g746(.A(new_n943), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n684), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n949), .B2(new_n946), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n940), .B2(new_n826), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n617), .A2(new_n266), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n943), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n948), .A2(new_n226), .A3(new_n725), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n940), .A2(new_n658), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(G1351gat));
  AND2_X1   g760(.A1(new_n700), .A2(new_n939), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n893), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT125), .ZN(new_n964));
  INV_X1    g763(.A(G197gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n965), .A3(new_n563), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n920), .A2(new_n921), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n967), .A2(new_n962), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(new_n563), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n969), .B2(new_n965), .ZN(G1352gat));
  XNOR2_X1  g769(.A(KEYINPUT126), .B(G204gat), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n963), .A2(new_n684), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g772(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n974));
  NOR2_X1   g773(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n967), .A2(new_n684), .A3(new_n962), .ZN(new_n977));
  OAI221_X1 g776(.A(new_n976), .B1(new_n974), .B2(new_n973), .C1(new_n977), .C2(new_n972), .ZN(G1353gat));
  NAND3_X1  g777(.A1(new_n964), .A2(new_n209), .A3(new_n617), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n967), .A2(new_n617), .A3(new_n962), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  AOI21_X1  g782(.A(G218gat), .B1(new_n964), .B2(new_n725), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n658), .A2(new_n210), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n984), .B1(new_n968), .B2(new_n985), .ZN(G1355gat));
endmodule


