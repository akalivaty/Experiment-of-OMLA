//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT80), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G141gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n207), .B(new_n209), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218));
  INV_X1    g017(.A(G113gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G120gat), .ZN(new_n220));
  INV_X1    g019(.A(G120gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G113gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G134gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G127gat), .ZN(new_n225));
  INV_X1    g024(.A(G127gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n225), .A2(new_n227), .A3(new_n218), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT69), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n219), .B2(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n219), .A2(G120gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n221), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n212), .A2(G141gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n210), .A2(G148gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n239), .A2(new_n215), .A3(new_n207), .A4(new_n209), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n217), .A2(new_n229), .A3(new_n236), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n223), .A2(new_n228), .B1(new_n230), .B2(new_n235), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n245), .A2(KEYINPUT82), .A3(new_n217), .A4(new_n240), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT81), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n217), .A2(new_n240), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n229), .A2(new_n236), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n217), .A2(new_n254), .A3(new_n240), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n251), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(KEYINPUT4), .A3(new_n245), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n247), .A2(new_n250), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n251), .A2(new_n253), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n246), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n261), .A2(new_n262), .A3(new_n249), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n261), .B2(new_n249), .ZN(new_n264));
  OAI211_X1 g063(.A(KEYINPUT5), .B(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n256), .A2(new_n250), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n244), .B1(new_n243), .B2(new_n246), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n241), .A2(new_n244), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n206), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT6), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n265), .A2(new_n206), .A3(new_n271), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n274), .B(new_n275), .C1(new_n272), .C2(KEYINPUT85), .ZN(new_n276));
  INV_X1    g075(.A(new_n270), .ZN(new_n277));
  NOR4_X1   g076(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT5), .A4(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n249), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT83), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n261), .A2(new_n262), .A3(new_n249), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n278), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n284), .A2(new_n285), .A3(new_n206), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n273), .B1(new_n276), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G8gat), .B(G36gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(KEYINPUT79), .ZN(new_n291));
  AND2_X1   g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G211gat), .A2(G218gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT75), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G211gat), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n298));
  NAND2_X1  g097(.A1(G211gat), .A2(G218gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(KEYINPUT74), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G197gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G204gat), .ZN(new_n305));
  INV_X1    g104(.A(G204gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G197gat), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n292), .B2(KEYINPUT22), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n301), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT74), .B1(new_n299), .B2(new_n302), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n294), .B(new_n300), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n310), .A2(new_n303), .A3(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n294), .A4(new_n300), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT29), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  NOR3_X1   g126(.A1(KEYINPUT68), .A2(G169gat), .A3(G176gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329));
  AND3_X1   g128(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n333));
  INV_X1    g132(.A(G169gat), .ZN(new_n334));
  INV_X1    g133(.A(G176gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(KEYINPUT26), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n327), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT27), .B(G183gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT27), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n341), .ZN(new_n345));
  INV_X1    g144(.A(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n339), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G183gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT27), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n351), .A2(new_n339), .A3(G190gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n338), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT24), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n327), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n346), .ZN(new_n358));
  NAND3_X1  g157(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n334), .A2(KEYINPUT64), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT64), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G169gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT65), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n361), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n360), .A2(new_n366), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n330), .B2(new_n331), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n335), .A2(KEYINPUT23), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT25), .B1(new_n375), .B2(G169gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT66), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n327), .A2(new_n378), .A3(new_n356), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n327), .B2(new_n356), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n358), .B(new_n359), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n355), .A2(new_n373), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n326), .B1(new_n354), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n336), .A2(KEYINPUT26), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n328), .A2(new_n329), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n371), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n351), .A2(KEYINPUT67), .ZN(new_n387));
  AOI21_X1  g186(.A(G190gat), .B1(new_n344), .B2(new_n341), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT28), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n327), .B(new_n386), .C1(new_n389), .C2(new_n352), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n355), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n377), .A2(new_n381), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n393), .A3(KEYINPUT78), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n325), .B1(new_n383), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n393), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n322), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n321), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n323), .A3(new_n394), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n322), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n399), .A2(new_n320), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n291), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n398), .A2(new_n291), .A3(new_n403), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n290), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n398), .A2(new_n290), .A3(new_n403), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n398), .A2(new_n403), .A3(KEYINPUT30), .A4(new_n290), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n287), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n318), .B(new_n301), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n254), .B1(new_n416), .B2(new_n400), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n255), .A2(new_n401), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n417), .A2(new_n251), .B1(new_n320), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G228gat), .A2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n320), .A2(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n421), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n316), .A2(new_n424), .A3(new_n319), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n257), .B1(new_n425), .B2(new_n254), .ZN(new_n426));
  OAI22_X1  g225(.A1(new_n419), .A2(new_n421), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n415), .B1(new_n427), .B2(G22gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n423), .A2(new_n426), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n400), .B1(new_n311), .B2(new_n315), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n251), .B1(new_n434), .B2(KEYINPUT3), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n421), .B1(new_n422), .B2(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n433), .A2(G22gat), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n425), .A2(new_n254), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n251), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n420), .B1(new_n320), .B2(new_n418), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n435), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n420), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n438), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n428), .A2(new_n432), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(G22gat), .B1(new_n433), .B2(new_n436), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(new_n438), .A3(new_n444), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n415), .A4(new_n431), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n446), .A2(KEYINPUT87), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT87), .B1(new_n446), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n414), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n390), .A2(new_n393), .A3(new_n245), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT70), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n396), .A2(new_n253), .ZN(new_n456));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT70), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n390), .A2(new_n393), .A3(new_n458), .A4(new_n245), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n455), .A2(new_n456), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT72), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(KEYINPUT34), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT32), .ZN(new_n467));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT33), .B1(new_n470), .B2(KEYINPUT71), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(KEYINPUT71), .B2(new_n470), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n459), .A3(new_n456), .ZN(new_n473));
  INV_X1    g272(.A(new_n457), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n467), .B(new_n472), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n470), .B1(new_n476), .B2(KEYINPUT32), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT33), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT73), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n466), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n466), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n484), .A2(new_n478), .A3(new_n470), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT73), .B(new_n483), .C1(new_n485), .C2(new_n475), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(KEYINPUT36), .A3(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n485), .A2(new_n483), .A3(new_n475), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n480), .A2(new_n466), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n487), .B1(new_n490), .B2(KEYINPUT36), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n243), .A2(new_n246), .A3(new_n250), .A4(new_n260), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT39), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT39), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n268), .A2(new_n498), .A3(new_n277), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n495), .B(new_n497), .C1(new_n499), .C2(new_n250), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n269), .A2(new_n256), .A3(new_n270), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n249), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n206), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n272), .B1(new_n492), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n500), .A2(KEYINPUT40), .A3(new_n206), .A4(new_n503), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n505), .B(new_n506), .C1(new_n407), .C2(new_n412), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n440), .A2(new_n441), .B1(new_n443), .B2(new_n420), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT86), .B1(new_n508), .B2(new_n438), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n509), .A2(new_n431), .B1(new_n447), .B2(new_n448), .ZN(new_n510));
  INV_X1    g309(.A(new_n449), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n265), .A2(new_n271), .ZN(new_n513));
  INV_X1    g312(.A(new_n206), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(new_n274), .A3(new_n275), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n398), .A2(new_n517), .A3(new_n403), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n320), .B1(new_n395), .B2(new_n397), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n399), .A2(new_n321), .A3(new_n402), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT37), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT38), .ZN(new_n522));
  INV_X1    g321(.A(new_n290), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n518), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n516), .A2(new_n273), .A3(new_n408), .A4(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n398), .A2(new_n291), .A3(new_n403), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT37), .B1(new_n526), .B2(new_n404), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n518), .A2(new_n523), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n507), .B(new_n512), .C1(new_n525), .C2(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n453), .A2(new_n491), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n273), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n512), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n480), .B(new_n466), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n523), .B1(new_n526), .B2(new_n404), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT35), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n410), .A4(new_n411), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n533), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n512), .A2(new_n482), .A3(new_n486), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT35), .B1(new_n414), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT89), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT89), .B(KEYINPUT35), .C1(new_n414), .C2(new_n539), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n531), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n547), .B2(new_n546), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT91), .B(G36gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G29gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n552), .A2(G29gat), .A3(G36gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n549), .B1(new_n557), .B2(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n559), .A2(KEYINPUT17), .ZN(new_n560));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT16), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(G1gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(G1gat), .B2(new_n561), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(G8gat), .Z(new_n565));
  AND2_X1   g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(KEYINPUT17), .ZN(new_n567));
  INV_X1    g366(.A(new_n559), .ZN(new_n568));
  INV_X1    g367(.A(new_n565), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n566), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(KEYINPUT18), .A3(new_n571), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n565), .B(new_n559), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n571), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G197gat), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT11), .B(G169gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT12), .Z(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n574), .A2(new_n586), .A3(new_n575), .A4(new_n578), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n544), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n224), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G162gat), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT7), .ZN(new_n597));
  INV_X1    g396(.A(G99gat), .ZN(new_n598));
  INV_X1    g397(.A(G106gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT8), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n597), .B(new_n600), .C1(G85gat), .C2(G92gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(G99gat), .B(G106gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n560), .A2(new_n567), .A3(new_n604), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n568), .A2(new_n603), .B1(KEYINPUT41), .B2(new_n591), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n595), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n594), .B1(new_n607), .B2(KEYINPUT96), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT97), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT97), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n605), .A2(new_n606), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n595), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n611), .A2(new_n614), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT93), .ZN(new_n620));
  INV_X1    g419(.A(G71gat), .ZN(new_n621));
  INV_X1    g420(.A(G78gat), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT92), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n620), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G57gat), .B(G64gat), .Z(new_n625));
  INV_X1    g424(.A(new_n619), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(KEYINPUT9), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  OR3_X1    g428(.A1(new_n627), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(KEYINPUT94), .A3(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n635), .A2(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G127gat), .B(G155gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT20), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G183gat), .B(G211gat), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n569), .B1(new_n635), .B2(KEYINPUT21), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n646), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n646), .B2(new_n651), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n618), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n635), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n604), .A2(new_n631), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n635), .B2(new_n604), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n658), .B2(KEYINPUT10), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(G230gat), .A3(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT98), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n662), .ZN(new_n668));
  INV_X1    g467(.A(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n590), .A2(new_n655), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT99), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n287), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(G1gat), .Z(G1324gat));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n674), .A2(new_n413), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G8gat), .B1(new_n674), .B2(new_n413), .ZN(new_n681));
  NOR2_X1   g480(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n682));
  MUX2_X1   g481(.A(KEYINPUT100), .B(new_n682), .S(new_n679), .Z(new_n683));
  AOI22_X1  g482(.A1(new_n680), .A2(new_n681), .B1(new_n678), .B2(new_n683), .ZN(G1325gat));
  XNOR2_X1  g483(.A(new_n491), .B(KEYINPUT101), .ZN(new_n685));
  OAI21_X1  g484(.A(G15gat), .B1(new_n674), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n534), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n674), .B2(new_n687), .ZN(G1326gat));
  INV_X1    g487(.A(new_n452), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NAND3_X1  g491(.A1(new_n453), .A2(new_n491), .A3(new_n530), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n533), .A2(new_n537), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n490), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n512), .A2(new_n482), .A3(new_n486), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n535), .A2(new_n410), .A3(new_n411), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n285), .B1(new_n284), .B2(new_n206), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT6), .B1(new_n284), .B2(new_n206), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n272), .A2(KEYINPUT85), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n697), .B1(new_n273), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n536), .B1(new_n696), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n695), .B1(new_n703), .B2(KEYINPUT89), .ZN(new_n704));
  INV_X1    g503(.A(new_n543), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n693), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n616), .A2(new_n617), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n652), .A2(new_n653), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n588), .A3(new_n672), .ZN(new_n710));
  NOR4_X1   g509(.A1(new_n708), .A2(G29gat), .A3(new_n287), .A4(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT103), .Z(new_n712));
  XOR2_X1   g511(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n544), .B2(new_n618), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n706), .A2(KEYINPUT44), .A3(new_n707), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n710), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n721), .B2(new_n287), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n714), .A2(new_n715), .A3(new_n722), .ZN(G1328gat));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724));
  AOI211_X1 g523(.A(new_n550), .B(new_n618), .C1(new_n724), .C2(KEYINPUT46), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n652), .A2(new_n653), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n671), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n590), .A2(new_n725), .A3(new_n697), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n724), .A2(KEYINPUT46), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT105), .B1(new_n721), .B2(new_n413), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n550), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n721), .A2(KEYINPUT105), .A3(new_n413), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(G1329gat));
  INV_X1    g533(.A(new_n491), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n735), .A3(new_n720), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G43gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n534), .A2(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n708), .A2(new_n710), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(KEYINPUT47), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n685), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n717), .A2(new_n718), .A3(new_n743), .A4(new_n720), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G43gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n741), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT106), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n740), .B1(new_n744), .B2(G43gat), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT47), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n742), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n742), .B(KEYINPUT107), .C1(new_n748), .C2(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1330gat));
  OAI21_X1  g555(.A(G50gat), .B1(new_n721), .B2(new_n512), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n708), .A2(new_n710), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n689), .A2(G50gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(KEYINPUT48), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n719), .A2(new_n452), .A3(new_n720), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n762), .A2(G50gat), .B1(new_n758), .B2(new_n759), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g563(.A1(new_n706), .A2(new_n655), .A3(new_n589), .A4(new_n671), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n287), .B(KEYINPUT109), .Z(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g572(.A1(new_n413), .A2(KEYINPUT110), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n413), .A2(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  AND2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n778), .B2(new_n779), .ZN(G1333gat));
  NOR2_X1   g581(.A1(new_n685), .A2(new_n621), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n766), .A2(KEYINPUT111), .A3(new_n767), .A4(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n621), .B1(new_n768), .B2(new_n534), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT50), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1334gat));
  NOR2_X1   g593(.A1(new_n768), .A2(new_n689), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n622), .ZN(G1335gat));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n709), .A2(new_n589), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n708), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n708), .B2(new_n798), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(KEYINPUT112), .B(new_n797), .C1(new_n708), .C2(new_n798), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n672), .A2(G85gat), .A3(new_n287), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n798), .A2(new_n672), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n719), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G85gat), .B1(new_n807), .B2(new_n287), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1336gat));
  NAND3_X1  g608(.A1(new_n799), .A2(KEYINPUT113), .A3(new_n801), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n777), .A2(new_n672), .A3(G92gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n797), .C1(new_n708), .C2(new_n798), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G92gat), .B1(new_n807), .B2(new_n413), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT52), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n719), .A2(new_n776), .A3(new_n806), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n818), .B2(G92gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n811), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n819), .B2(new_n820), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n817), .B1(new_n822), .B2(new_n823), .ZN(G1337gat));
  XNOR2_X1  g623(.A(KEYINPUT115), .B(G99gat), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n672), .A2(new_n534), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n802), .A2(new_n803), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n807), .B2(new_n685), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1338gat));
  NOR3_X1   g628(.A1(new_n672), .A2(G106gat), .A3(new_n512), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n802), .A2(new_n803), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G106gat), .B1(new_n807), .B2(new_n512), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n810), .A2(new_n813), .A3(new_n830), .ZN(new_n835));
  OAI21_X1  g634(.A(G106gat), .B1(new_n807), .B2(new_n689), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT116), .B1(new_n837), .B2(KEYINPUT53), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n839), .B(new_n833), .C1(new_n835), .C2(new_n836), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n834), .B1(new_n838), .B2(new_n840), .ZN(G1339gat));
  NOR3_X1   g640(.A1(new_n654), .A2(new_n588), .A3(new_n671), .ZN(new_n842));
  XNOR2_X1  g641(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n669), .B1(new_n661), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n659), .A2(new_n660), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n661), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT118), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n846), .B2(new_n849), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n570), .A2(new_n571), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n576), .A2(new_n577), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n583), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n587), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n849), .A3(KEYINPUT55), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n667), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n857), .A2(new_n707), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n861), .B1(new_n667), .B2(new_n670), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n588), .A2(new_n667), .A3(new_n863), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n857), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n865), .B1(new_n868), .B2(new_n707), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n842), .B1(new_n869), .B2(new_n709), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n770), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n696), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n776), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n219), .A3(new_n588), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n709), .ZN(new_n875));
  INV_X1    g674(.A(new_n842), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n776), .A2(new_n287), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n452), .A2(new_n534), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n880), .A2(new_n589), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT119), .B1(new_n881), .B2(G113gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(G1340gat));
  OAI21_X1  g683(.A(G120gat), .B1(new_n880), .B2(new_n672), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n672), .A2(G120gat), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n696), .A3(new_n777), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT120), .Z(G1341gat));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n226), .A3(new_n726), .ZN(new_n890));
  OAI21_X1  g689(.A(G127gat), .B1(new_n880), .B2(new_n709), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1342gat));
  NOR2_X1   g691(.A1(new_n618), .A2(new_n697), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n224), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n872), .A2(KEYINPUT56), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n880), .B2(new_n618), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT56), .B1(new_n872), .B2(new_n894), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1343gat));
  NAND3_X1  g697(.A1(new_n588), .A2(new_n667), .A3(new_n863), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n854), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n618), .B1(new_n900), .B2(new_n866), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n726), .B1(new_n901), .B2(new_n865), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n452), .B1(new_n902), .B2(new_n842), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT57), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  INV_X1    g704(.A(new_n512), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n899), .B1(new_n853), .B2(new_n856), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n618), .B1(new_n907), .B2(new_n866), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n726), .B1(new_n908), .B2(new_n865), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n905), .B(new_n906), .C1(new_n909), .C2(new_n842), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n735), .A2(new_n776), .A3(new_n287), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G141gat), .B1(new_n912), .B2(new_n589), .ZN(new_n913));
  OR2_X1    g712(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n685), .A2(new_n906), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n870), .A2(new_n915), .A3(new_n770), .A4(new_n776), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n589), .A2(G141gat), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n916), .A2(new_n917), .B1(KEYINPUT121), .B2(KEYINPUT58), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n913), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n914), .B1(new_n913), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1344gat));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  AOI211_X1 g721(.A(new_n922), .B(G148gat), .C1(new_n916), .C2(new_n671), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n912), .B2(new_n672), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT57), .B1(new_n870), .B2(new_n512), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n905), .B(new_n452), .C1(new_n902), .C2(new_n842), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n911), .A2(KEYINPUT59), .A3(new_n671), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n923), .B1(new_n929), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g729(.A(G155gat), .B1(new_n912), .B2(new_n709), .ZN(new_n931));
  INV_X1    g730(.A(new_n916), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n709), .A2(G155gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n912), .B2(new_n618), .ZN(new_n935));
  INV_X1    g734(.A(G162gat), .ZN(new_n936));
  INV_X1    g735(.A(new_n915), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n871), .A2(new_n936), .A3(new_n893), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(G1347gat));
  NOR2_X1   g738(.A1(new_n771), .A2(new_n413), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n877), .A2(new_n879), .A3(new_n940), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n941), .A2(new_n589), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n942), .A2(new_n943), .A3(G169gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n942), .B2(G169gat), .ZN(new_n945));
  INV_X1    g744(.A(new_n287), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n870), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n777), .A2(new_n539), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n287), .B(new_n949), .C1(new_n909), .C2(new_n842), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n588), .A2(new_n363), .A3(new_n365), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n944), .A2(new_n945), .B1(new_n953), .B2(new_n954), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n941), .B2(new_n672), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n671), .A2(new_n335), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n953), .B2(new_n957), .ZN(G1349gat));
  OAI21_X1  g757(.A(G183gat), .B1(new_n941), .B2(new_n709), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n726), .A2(new_n340), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n951), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g761(.A1(new_n950), .A2(new_n952), .A3(new_n346), .A4(new_n707), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n877), .A2(new_n707), .A3(new_n879), .A4(new_n940), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n964), .A2(new_n965), .A3(G190gat), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n964), .B2(G190gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n963), .B(KEYINPUT124), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1351gat));
  NAND2_X1  g771(.A1(new_n937), .A2(new_n776), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n870), .A2(new_n946), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(G197gat), .B1(new_n974), .B2(new_n588), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n940), .A2(new_n685), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n925), .A2(new_n926), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n589), .A2(new_n304), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NAND4_X1  g778(.A1(new_n925), .A2(new_n671), .A3(new_n926), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G204gat), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n672), .A2(G204gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n974), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n974), .A2(new_n985), .A3(new_n982), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n981), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(KEYINPUT125), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n981), .A2(new_n989), .A3(new_n984), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n295), .A3(new_n726), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n925), .A2(new_n726), .A3(new_n926), .A4(new_n976), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(G211gat), .ZN(new_n994));
  NOR2_X1   g793(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n994), .A2(new_n995), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(G1354gat));
  NAND3_X1  g799(.A1(new_n925), .A2(new_n926), .A3(new_n976), .ZN(new_n1001));
  OAI21_X1  g800(.A(G218gat), .B1(new_n1001), .B2(new_n618), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n974), .A2(new_n296), .A3(new_n707), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(KEYINPUT127), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1002), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1005), .A2(new_n1007), .ZN(G1355gat));
endmodule


