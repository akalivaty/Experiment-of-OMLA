//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(G146), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  OAI211_X1 g007(.A(G128), .B(new_n190), .C1(new_n191), .C2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n195), .B(new_n196), .C1(KEYINPUT1), .C2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(G125), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT0), .A4(G128), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n199), .B1(G125), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G224), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G953), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n204), .B(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G110), .B(G122), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT73), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT73), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G101), .ZN(new_n220));
  AOI21_X1  g034(.A(G101), .B1(new_n210), .B2(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  INV_X1    g038(.A(G119), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT64), .B1(new_n225), .B2(G116), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(G119), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT2), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT2), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n230), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n230), .B2(new_n232), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n224), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n227), .B1(new_n228), .B2(G119), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n225), .A2(KEYINPUT64), .A3(G116), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n232), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n237), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n230), .A2(new_n232), .A3(new_n237), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT65), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n219), .A2(new_n248), .A3(G101), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n223), .A2(new_n240), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n233), .B1(new_n231), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n243), .B2(new_n251), .ZN(new_n253));
  AOI21_X1  g067(.A(G104), .B1(new_n213), .B2(new_n215), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n210), .A2(G107), .ZN(new_n255));
  OAI21_X1  g069(.A(G101), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n253), .A2(new_n246), .A3(new_n222), .A4(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n209), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT77), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT77), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n262), .A3(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n240), .A2(new_n247), .ZN(new_n265));
  INV_X1    g079(.A(G101), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(G104), .B2(new_n212), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT73), .B(G107), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(new_n211), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(new_n270), .B2(new_n217), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n249), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n209), .B(new_n257), .C1(new_n265), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n250), .A2(KEYINPUT75), .A3(new_n209), .A4(new_n257), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n258), .A2(new_n259), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n278), .A2(KEYINPUT76), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT76), .B1(new_n278), .B2(new_n279), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n208), .B(new_n264), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n204), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(new_n209), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n256), .A2(new_n222), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(new_n238), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n243), .A2(new_n251), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n252), .B(KEYINPUT79), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n253), .A2(new_n246), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n287), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n286), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n284), .B(new_n294), .C1(new_n208), .C2(new_n283), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n295), .B2(new_n278), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n282), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n282), .A2(new_n296), .A3(new_n298), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n188), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G217), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(G234), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n225), .A2(G128), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n225), .A2(G128), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(KEYINPUT23), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT24), .B(G110), .Z(new_n311));
  XNOR2_X1  g125(.A(G119), .B(G128), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n310), .A2(G110), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT16), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n316), .A2(KEYINPUT16), .A3(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G146), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(G146), .B1(new_n318), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n313), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n310), .A2(G110), .B1(new_n311), .B2(new_n312), .ZN(new_n324));
  XNOR2_X1  g138(.A(G125), .B(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n192), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n320), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(new_n327), .A3(new_n332), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n304), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT70), .B1(KEYINPUT71), .B2(KEYINPUT25), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n306), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT70), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n334), .A2(new_n340), .A3(new_n304), .A4(new_n335), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n341), .A2(KEYINPUT71), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n339), .B1(new_n342), .B2(KEYINPUT25), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n334), .A2(new_n335), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n305), .A2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT72), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n338), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n305), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT25), .B1(new_n341), .B2(KEYINPUT71), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT72), .B(new_n346), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n203), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT11), .ZN(new_n355));
  INV_X1    g169(.A(G134), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(G137), .ZN(new_n357));
  INV_X1    g171(.A(G137), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT11), .A3(G134), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(G137), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G131), .ZN(new_n362));
  INV_X1    g176(.A(G131), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n357), .A2(new_n359), .A3(new_n363), .A4(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n354), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n194), .A2(new_n198), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n356), .A2(G137), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n358), .A2(G134), .ZN(new_n369));
  OAI21_X1  g183(.A(G131), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n238), .A2(new_n239), .A3(new_n224), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT65), .B1(new_n245), .B2(new_n246), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n366), .B(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n203), .B1(new_n362), .B2(new_n364), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n367), .A2(new_n371), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n240), .B(new_n247), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n380));
  INV_X1    g194(.A(G237), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n330), .A3(G210), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G101), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n385), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n375), .B2(new_n378), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT67), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n375), .B2(new_n390), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n380), .B(new_n389), .C1(new_n391), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT68), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n375), .A2(new_n378), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n376), .A2(new_n377), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT28), .B1(new_n398), .B2(new_n265), .ZN(new_n399));
  OAI22_X1  g213(.A1(new_n397), .A2(new_n390), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n400), .A2(KEYINPUT68), .A3(new_n389), .A4(new_n380), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n373), .A2(new_n374), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n372), .A2(new_n366), .A3(KEYINPUT30), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n376), .B2(new_n377), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n375), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT29), .B1(new_n407), .B2(new_n388), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n396), .A2(new_n401), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n391), .A2(new_n410), .ZN(new_n411));
  AOI211_X1 g225(.A(KEYINPUT69), .B(new_n390), .C1(new_n375), .C2(new_n378), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n411), .A2(new_n412), .A3(new_n399), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n389), .A2(KEYINPUT29), .ZN(new_n414));
  AOI21_X1  g228(.A(G902), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G472), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n380), .B1(new_n391), .B2(new_n393), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT66), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT31), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n386), .A2(new_n387), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n398), .B2(new_n265), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n406), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n419), .A2(KEYINPUT31), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n422), .B(new_n406), .C1(new_n419), .C2(KEYINPUT31), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n418), .A2(new_n388), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G472), .A2(G902), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT32), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT32), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n389), .B1(new_n400), .B2(new_n380), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n425), .A2(new_n426), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n431), .B(new_n428), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n353), .B1(new_n417), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n330), .A2(G227), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n256), .A2(new_n198), .A3(new_n194), .A4(new_n222), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT74), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT10), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT10), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(KEYINPUT74), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n223), .A2(new_n354), .A3(new_n249), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n365), .ZN(new_n449));
  INV_X1    g263(.A(new_n365), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(new_n450), .A3(new_n446), .A4(new_n447), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n441), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n441), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n287), .A2(new_n367), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n442), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT12), .B1(new_n455), .B2(new_n365), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  AOI211_X1 g271(.A(new_n457), .B(new_n450), .C1(new_n454), .C2(new_n442), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n437), .B(new_n304), .C1(new_n452), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n451), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n440), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n449), .A2(new_n451), .A3(new_n441), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(G469), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n437), .A2(new_n304), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT9), .B(G234), .ZN(new_n469));
  OAI21_X1  g283(.A(G221), .B1(new_n469), .B2(G902), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n469), .A2(new_n303), .A3(G953), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n213), .A2(new_n215), .ZN(new_n473));
  INV_X1    g287(.A(G122), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G116), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n228), .A2(G122), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G116), .B(G122), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n269), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n197), .B2(G143), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n189), .A2(KEYINPUT81), .A3(G128), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n197), .A2(G143), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n356), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT13), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT82), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT82), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n483), .A2(new_n484), .A3(new_n491), .A4(KEYINPUT13), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n485), .A2(new_n489), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n490), .A2(new_n492), .A3(new_n486), .A4(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n488), .B1(new_n494), .B2(G134), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n485), .A2(new_n356), .A3(new_n486), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n356), .B1(new_n485), .B2(new_n486), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT83), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n480), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(new_n474), .B2(G116), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n475), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n476), .A2(KEYINPUT14), .ZN(new_n503));
  OAI21_X1  g317(.A(G107), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n269), .A2(new_n479), .A3(KEYINPUT83), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n472), .B1(new_n495), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT85), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n510), .B(new_n472), .C1(new_n495), .C2(new_n507), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n495), .A2(new_n507), .ZN(new_n513));
  INV_X1    g327(.A(new_n472), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR4_X1   g329(.A1(new_n495), .A2(new_n507), .A3(KEYINPUT84), .A4(new_n472), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n509), .B(new_n511), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n304), .ZN(new_n518));
  INV_X1    g332(.A(G478), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n517), .A2(new_n304), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G237), .A2(G953), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(G143), .A3(G214), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(G143), .B1(new_n529), .B2(G214), .ZN(new_n532));
  OAI21_X1  g346(.A(G131), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n381), .A2(new_n330), .A3(G214), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n189), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n363), .A3(new_n530), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT80), .B(KEYINPUT19), .Z(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n325), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n315), .A2(new_n317), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT80), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n540), .B1(new_n541), .B2(KEYINPUT19), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n542), .A3(new_n192), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(new_n320), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(KEYINPUT18), .B(G131), .C1(new_n531), .C2(new_n532), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(G146), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n326), .ZN(new_n547));
  NAND2_X1  g361(.A1(KEYINPUT18), .A2(G131), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n535), .A2(new_n530), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G113), .B(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n210), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n321), .A2(new_n322), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n533), .A2(new_n557), .A3(new_n536), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n363), .B1(new_n535), .B2(new_n530), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT17), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n553), .A3(new_n550), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(G475), .A2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT20), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT20), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(new_n562), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n553), .B1(new_n561), .B2(new_n550), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n304), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n566), .A2(new_n568), .B1(G475), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(G234), .A2(G237), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(G902), .A3(G953), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT87), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT21), .B(G898), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n573), .A2(G952), .A3(new_n330), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n471), .A2(new_n528), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n302), .A2(new_n436), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  NOR2_X1   g398(.A1(new_n347), .A2(new_n352), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT88), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(G472), .C1(new_n427), .C2(G902), .ZN(new_n587));
  INV_X1    g401(.A(G472), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n391), .A2(new_n393), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n392), .B(new_n390), .C1(new_n375), .C2(new_n378), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n388), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n425), .A2(new_n426), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n588), .B1(new_n593), .B2(new_n304), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT88), .B1(new_n593), .B2(new_n428), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n585), .B(new_n587), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n471), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT89), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n517), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n513), .A2(new_n514), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(KEYINPUT33), .A3(new_n508), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n519), .A2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n518), .A2(new_n519), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n572), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n282), .A2(new_n296), .A3(new_n298), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n298), .B1(new_n282), .B2(new_n296), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n187), .B(new_n606), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n598), .A2(new_n580), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND2_X1  g427(.A1(new_n571), .A2(G475), .ZN(new_n614));
  INV_X1    g428(.A(new_n568), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n567), .B1(new_n563), .B2(new_n564), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT90), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT90), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n566), .A2(new_n618), .A3(new_n568), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n580), .B(KEYINPUT91), .Z(new_n621));
  AND4_X1   g435(.A1(new_n528), .A2(new_n614), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n622), .B(new_n187), .C1(new_n608), .C2(new_n607), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(KEYINPUT92), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT92), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n302), .B2(new_n622), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n598), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT93), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NOR2_X1   g444(.A1(new_n333), .A2(KEYINPUT36), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n328), .B(new_n631), .Z(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n345), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n343), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n587), .B(new_n635), .C1(new_n594), .C2(new_n595), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT94), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n427), .B2(G902), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n586), .B1(new_n427), .B2(new_n429), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n587), .A4(new_n635), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n637), .A2(new_n302), .A3(new_n582), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  NAND2_X1  g459(.A1(new_n300), .A2(new_n301), .ZN(new_n646));
  INV_X1    g460(.A(new_n528), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n620), .A2(new_n614), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n578), .B1(new_n575), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(new_n651), .A3(new_n187), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n416), .A2(G472), .B1(new_n430), .B2(new_n434), .ZN(new_n654));
  INV_X1    g468(.A(new_n635), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n471), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  OAI21_X1  g472(.A(new_n304), .B1(new_n379), .B2(new_n389), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n388), .B1(new_n406), .B2(new_n375), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n435), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n572), .B1(new_n525), .B2(new_n527), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n187), .A2(new_n662), .A3(new_n655), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n300), .A2(new_n301), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n665), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n646), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT96), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT96), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n664), .A2(new_n671), .A3(new_n666), .A4(new_n668), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n468), .A2(new_n470), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n650), .B(KEYINPUT39), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT40), .Z(new_n676));
  NAND3_X1  g490(.A1(new_n670), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT97), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n670), .A2(new_n672), .A3(KEYINPUT97), .A4(new_n676), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  OAI21_X1  g496(.A(new_n187), .B1(new_n607), .B2(new_n608), .ZN(new_n683));
  INV_X1    g497(.A(new_n650), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n606), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT98), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT98), .ZN(new_n687));
  AOI211_X1 g501(.A(new_n650), .B(new_n572), .C1(new_n604), .C2(new_n605), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n302), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n686), .A2(new_n689), .A3(new_n656), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n646), .A2(new_n187), .A3(new_n580), .A4(new_n606), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n417), .A2(new_n435), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n452), .A2(new_n460), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n470), .A3(new_n461), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n694), .A2(new_n585), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n692), .B1(new_n693), .B2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n654), .A2(new_n353), .A3(new_n697), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n610), .A2(new_n701), .A3(KEYINPUT99), .A4(new_n580), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND2_X1  g519(.A1(new_n623), .A2(KEYINPUT92), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n302), .A2(new_n625), .A3(new_n622), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n699), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n228), .ZN(G18));
  AOI21_X1  g523(.A(new_n655), .B1(new_n417), .B2(new_n435), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n528), .A2(new_n581), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n302), .A2(new_n710), .A3(new_n711), .A4(new_n698), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND2_X1  g527(.A1(new_n343), .A2(new_n346), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT69), .B1(new_n397), .B2(new_n390), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n399), .B1(new_n391), .B2(new_n410), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n389), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT100), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n433), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n638), .B(new_n715), .C1(new_n722), .C2(new_n429), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n621), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n697), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n302), .A2(new_n724), .A3(new_n663), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NOR3_X1   g542(.A1(new_n683), .A2(new_n685), .A3(new_n697), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n718), .A2(new_n719), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n388), .A3(new_n721), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n592), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n594), .B1(new_n732), .B2(new_n428), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT101), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n635), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n638), .B(new_n635), .C1(new_n722), .C2(new_n429), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT101), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT102), .B(G125), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G27));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n300), .A2(new_n688), .A3(new_n187), .A4(new_n301), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n465), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n463), .A2(KEYINPUT103), .A3(G469), .A4(new_n464), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n461), .A3(new_n467), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n470), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n588), .B1(new_n409), .B2(new_n415), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n751), .B2(new_n435), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n430), .A2(new_n434), .A3(KEYINPUT104), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n714), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n742), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n607), .A2(new_n608), .A3(new_n188), .ZN(new_n756));
  INV_X1    g570(.A(new_n748), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n436), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT105), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(new_n688), .A3(new_n757), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n431), .B1(new_n593), .B2(new_n428), .ZN(new_n762));
  AOI211_X1 g576(.A(KEYINPUT32), .B(new_n429), .C1(new_n591), .C2(new_n592), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n751), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n417), .A3(new_n753), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n715), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT42), .B1(new_n761), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT105), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n654), .A2(new_n748), .A3(new_n353), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n756), .A3(new_n758), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n760), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT106), .B(G131), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G33));
  NAND4_X1  g588(.A1(new_n756), .A2(new_n436), .A3(new_n651), .A4(new_n757), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n769), .A2(KEYINPUT107), .A3(new_n651), .A4(new_n756), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  NAND3_X1  g594(.A1(new_n300), .A2(new_n187), .A3(new_n301), .ZN(new_n781));
  INV_X1    g595(.A(new_n602), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n517), .B2(new_n599), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n783), .A2(new_n603), .B1(new_n518), .B2(new_n519), .ZN(new_n784));
  INV_X1    g598(.A(new_n572), .ZN(new_n785));
  OR3_X1    g599(.A1(new_n784), .A2(KEYINPUT43), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT43), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n640), .A2(new_n587), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n635), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n781), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n463), .A2(new_n464), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n437), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n467), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n461), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT108), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n797), .A2(new_n467), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT46), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(KEYINPUT108), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n470), .A3(new_n674), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n793), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n358), .ZN(G39));
  NOR3_X1   g621(.A1(new_n743), .A2(new_n694), .A3(new_n585), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n470), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT47), .B1(new_n804), .B2(new_n470), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT109), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  NAND2_X1  g630(.A1(new_n696), .A2(new_n461), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(KEYINPUT49), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(KEYINPUT49), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n818), .A2(new_n819), .A3(new_n785), .A4(new_n784), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n668), .A2(new_n666), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n715), .A2(new_n187), .A3(new_n470), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n662), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n647), .A2(new_n785), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n597), .A2(new_n302), .A3(new_n621), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n643), .A3(new_n712), .A4(new_n727), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n708), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n673), .A2(new_n585), .A3(new_n640), .A4(new_n587), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n609), .A2(new_n829), .A3(new_n725), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n762), .A2(new_n763), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n585), .B1(new_n831), .B2(new_n750), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n673), .A2(new_n711), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n832), .A2(new_n683), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT110), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n597), .A2(new_n621), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n836), .B(new_n583), .C1(new_n837), .C2(new_n609), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n828), .A2(new_n839), .A3(new_n703), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n648), .A2(new_n528), .A3(new_n650), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n756), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n756), .A2(KEYINPUT111), .A3(new_n841), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n656), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n749), .A2(new_n738), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n779), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n840), .A2(new_n772), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n663), .B(new_n187), .C1(new_n607), .C2(new_n608), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n635), .B(new_n650), .C1(new_n435), .C2(new_n661), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n757), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n690), .A2(new_n657), .A3(new_n739), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n738), .A2(new_n729), .B1(new_n653), .B2(new_n656), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n690), .A4(new_n853), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT53), .B1(new_n849), .B2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n755), .A2(KEYINPUT105), .A3(new_n759), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n768), .B1(new_n767), .B2(new_n770), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n701), .B1(new_n624), .B2(new_n626), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n643), .A2(new_n712), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n825), .B(new_n187), .C1(new_n608), .C2(new_n607), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n829), .A2(new_n725), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n723), .A2(new_n725), .A3(new_n697), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n867), .A2(new_n868), .B1(new_n851), .B2(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n703), .A2(new_n864), .A3(new_n865), .A4(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n779), .A2(new_n846), .A3(new_n847), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n863), .A2(new_n871), .A3(new_n839), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n855), .A2(new_n858), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n856), .A2(new_n857), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(KEYINPUT53), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT54), .B1(new_n860), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n788), .A2(KEYINPUT112), .A3(new_n578), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n786), .A2(new_n578), .A3(new_n787), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT112), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n723), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n697), .A2(new_n187), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n821), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT113), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT113), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n821), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n883), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT50), .Z(new_n890));
  NOR2_X1   g704(.A1(new_n781), .A2(new_n697), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n662), .A2(new_n353), .A3(new_n579), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n893), .A2(new_n572), .A3(new_n784), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n879), .A2(new_n882), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n738), .A3(new_n891), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT114), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(KEYINPUT114), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n890), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT115), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n890), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n809), .A2(new_n810), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n470), .B2(new_n817), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n756), .A3(new_n883), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n901), .A2(KEYINPUT51), .A3(new_n903), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n895), .A2(new_n754), .A3(new_n891), .ZN(new_n908));
  XNOR2_X1  g722(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(G952), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n911), .B(G953), .C1(new_n893), .C2(new_n606), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT48), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(KEYINPUT116), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n895), .A2(new_n754), .A3(new_n891), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n883), .A2(new_n302), .A3(new_n698), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n910), .A2(new_n912), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT117), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n906), .A2(new_n890), .A3(new_n899), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n873), .B2(new_n874), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n828), .A2(new_n839), .A3(new_n703), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n767), .A2(KEYINPUT53), .A3(new_n770), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n875), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n859), .A2(new_n925), .A3(new_n872), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n923), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  AND4_X1   g743(.A1(new_n878), .A2(new_n907), .A3(new_n921), .A4(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(G952), .A2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n824), .B1(new_n930), .B2(new_n931), .ZN(G75));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n923), .A2(new_n928), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(G902), .ZN(new_n935));
  INV_X1    g749(.A(G210), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n264), .B1(new_n280), .B2(new_n281), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n207), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n282), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT55), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n330), .A2(G952), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n937), .A2(new_n941), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(G51));
  XNOR2_X1  g761(.A(new_n695), .B(KEYINPUT118), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n934), .A2(KEYINPUT54), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(new_n929), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n466), .B(KEYINPUT57), .Z(new_n951));
  OAI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n935), .A2(new_n797), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n943), .B1(new_n952), .B2(new_n953), .ZN(G54));
  NAND4_X1  g768(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n955));
  INV_X1    g769(.A(new_n563), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n955), .A2(KEYINPUT119), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n944), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT119), .B1(new_n955), .B2(new_n956), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G60));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT59), .Z(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n878), .B2(new_n929), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n944), .B1(new_n963), .B2(new_n783), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n949), .A2(new_n929), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n962), .B(new_n782), .C1(new_n517), .C2(new_n599), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT120), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT120), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n965), .A2(new_n969), .A3(new_n966), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n964), .B1(new_n968), .B2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT121), .Z(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT60), .Z(new_n974));
  AND4_X1   g788(.A1(new_n859), .A2(new_n925), .A3(new_n872), .A4(new_n927), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n860), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n344), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n943), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n979), .A2(new_n934), .A3(new_n633), .A4(new_n974), .ZN(new_n980));
  INV_X1    g794(.A(new_n974), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n923), .B2(new_n928), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n982), .B2(new_n633), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n978), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n978), .B(KEYINPUT61), .C1(new_n980), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(G66));
  NAND2_X1  g802(.A1(new_n840), .A2(new_n330), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT123), .Z(new_n990));
  OAI21_X1  g804(.A(G953), .B1(new_n576), .B2(new_n205), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n938), .B1(G898), .B2(new_n330), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(G69));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n856), .A2(new_n690), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n754), .A2(new_n851), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n805), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n779), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n998), .A2(new_n806), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n815), .A2(new_n1000), .A3(new_n863), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n330), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n403), .A2(new_n405), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n539), .A2(new_n542), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n649), .A2(G953), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT125), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n436), .B1(new_n606), .B2(new_n825), .ZN(new_n1010));
  OR3_X1    g824(.A1(new_n1010), .A2(new_n675), .A3(new_n781), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(new_n793), .B2(new_n805), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n813), .B2(new_n814), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT62), .B1(new_n681), .B2(new_n996), .ZN(new_n1014));
  AND4_X1   g828(.A1(KEYINPUT62), .A2(new_n679), .A3(new_n680), .A4(new_n996), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1005), .A2(G953), .ZN(new_n1017));
  AOI22_X1  g831(.A1(new_n1002), .A2(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n330), .B1(G227), .B2(G900), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT124), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n995), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1020), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1008), .B1(new_n1001), .B2(new_n330), .ZN(new_n1024));
  OAI211_X1 g838(.A(KEYINPUT126), .B(new_n1022), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(G72));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  OAI21_X1  g843(.A(new_n1029), .B1(new_n1001), .B2(new_n840), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n407), .A2(new_n389), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n943), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1013), .B(new_n925), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n1029), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n660), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1029), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n1031), .A2(new_n660), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1038), .B1(new_n860), .B2(new_n877), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1039), .A2(KEYINPUT127), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1039), .A2(KEYINPUT127), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(G57));
endmodule


