//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116, new_n1117, new_n1118;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  INV_X1    g038(.A(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G2104), .ZN(new_n465));
  OAI22_X1  g040(.A1(new_n462), .A2(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n460), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  INV_X1    g045(.A(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G136), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n460), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  INV_X1    g053(.A(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n480), .A2(new_n482), .A3(G126), .A4(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n480), .A2(new_n482), .A3(G138), .A4(new_n461), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n460), .A2(new_n490), .A3(G138), .A4(new_n461), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(G164));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n499), .B2(KEYINPUT66), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .A3(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n493), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G50), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n504), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n497), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n500), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  NAND2_X1  g087(.A1(new_n494), .A2(new_n496), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n502), .B2(new_n504), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G89), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n505), .A2(G51), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n497), .A2(G63), .A3(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n515), .A2(new_n516), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(KEYINPUT67), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(KEYINPUT67), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(G168));
  NAND2_X1  g098(.A1(G77), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G64), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n514), .A2(G90), .B1(new_n505), .B2(G52), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n526), .A2(KEYINPUT68), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  NAND2_X1  g108(.A1(G68), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G56), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n513), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT69), .Z(new_n538));
  AOI22_X1  g113(.A1(new_n514), .A2(G81), .B1(new_n505), .B2(G43), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT70), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n505), .A2(G53), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n550));
  INV_X1    g125(.A(G65), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n494), .B2(new_n496), .ZN(new_n553));
  NOR3_X1   g128(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n514), .A2(G91), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n549), .A2(new_n557), .A3(new_n558), .ZN(G299));
  AND2_X1   g134(.A1(new_n521), .A2(new_n522), .ZN(G286));
  NAND2_X1  g135(.A1(new_n514), .A2(G87), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n505), .A2(G49), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  NAND2_X1  g139(.A1(new_n505), .A2(G48), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT72), .Z(new_n566));
  AOI22_X1  g141(.A1(new_n497), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n499), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n570), .B2(new_n508), .ZN(G305));
  AOI22_X1  g146(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n499), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(G47), .B2(new_n505), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n514), .A2(G85), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(G301), .A2(G868), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT73), .Z(new_n579));
  NAND3_X1  g154(.A1(new_n497), .A2(new_n507), .A3(G92), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n505), .A2(G54), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  NOR3_X1   g159(.A1(new_n550), .A2(new_n584), .A3(new_n553), .ZN(new_n585));
  AND2_X1   g160(.A1(G79), .A2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n582), .B(new_n583), .C1(new_n587), .C2(new_n499), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n579), .B1(G868), .B2(new_n589), .ZN(G284));
  OAI21_X1  g165(.A(new_n579), .B1(G868), .B2(new_n589), .ZN(G321));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(G299), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G168), .B2(new_n592), .ZN(G280));
  XOR2_X1   g169(.A(G280), .B(KEYINPUT74), .Z(G297));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n538), .A2(new_n539), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n592), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n588), .A2(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n592), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n471), .A2(G135), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n473), .A2(G123), .ZN(new_n604));
  OAI21_X1  g179(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n461), .A2(G111), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(G2096), .Z(new_n608));
  NAND3_X1  g183(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(G2100), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(G156));
  XOR2_X1   g188(.A(KEYINPUT76), .B(G2438), .Z(new_n614));
  XNOR2_X1  g189(.A(G2427), .B(G2430), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT15), .B(G2435), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT14), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2451), .B(G2454), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n621), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n627), .A2(G14), .ZN(G401));
  XOR2_X1   g203(.A(G2084), .B(G2090), .Z(new_n629));
  XNOR2_X1  g204(.A(G2072), .B(G2078), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT17), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2067), .B(G2678), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n630), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT78), .ZN(new_n635));
  INV_X1    g210(.A(new_n629), .ZN(new_n636));
  NOR3_X1   g211(.A1(new_n631), .A2(new_n636), .A3(new_n632), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT79), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n629), .A2(new_n632), .A3(new_n630), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT77), .B(KEYINPUT18), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n635), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT80), .Z(new_n643));
  XNOR2_X1  g218(.A(G2096), .B(G2100), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G227));
  XOR2_X1   g221(.A(G1971), .B(G1976), .Z(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1956), .B(G2474), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1961), .B(G1966), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n649), .A2(KEYINPUT83), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  NOR3_X1   g232(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G1986), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT84), .B(G1981), .Z(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G229));
  MUX2_X1   g243(.A(G6), .B(G305), .S(G16), .Z(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT32), .B(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(G16), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G22), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(G166), .B2(new_n672), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1971), .ZN(new_n675));
  NOR2_X1   g250(.A1(G16), .A2(G23), .ZN(new_n676));
  INV_X1    g251(.A(G288), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(G16), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT33), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n671), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT34), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n672), .A2(G24), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n576), .B2(new_n672), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n683), .B(new_n684), .S(KEYINPUT87), .Z(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n473), .A2(G119), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT85), .Z(new_n689));
  INV_X1    g264(.A(G131), .ZN(new_n690));
  OAI21_X1  g265(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n461), .A2(G107), .ZN(new_n692));
  OAI22_X1  g267(.A1(new_n462), .A2(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT86), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT35), .B(G1991), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n682), .A2(new_n687), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(KEYINPUT88), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(G29), .A2(G32), .ZN(new_n704));
  AOI22_X1  g279(.A1(G141), .A2(new_n471), .B1(new_n473), .B2(G129), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT26), .Z(new_n707));
  INV_X1    g282(.A(G105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n707), .C1(new_n708), .C2(new_n465), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT95), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n607), .A2(new_n710), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT96), .ZN(new_n716));
  INV_X1    g291(.A(G11), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT31), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n714), .A2(new_n716), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G16), .A2(G21), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G168), .B2(G16), .ZN(new_n722));
  INV_X1    g297(.A(G1966), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(G171), .A2(G16), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G1961), .C1(G5), .C2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT97), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n711), .A2(new_n713), .ZN(new_n728));
  OR2_X1    g303(.A1(G29), .A2(G33), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n471), .A2(G139), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT25), .Z(new_n732));
  AOI22_X1  g307(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n730), .B(new_n732), .C1(new_n461), .C2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n729), .B1(new_n734), .B2(new_n710), .ZN(new_n735));
  INV_X1    g310(.A(G2072), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT93), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n724), .A2(new_n727), .A3(new_n728), .A4(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n725), .B1(G5), .B2(G16), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n720), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n735), .A2(new_n736), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  OR2_X1    g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n745), .A2(new_n710), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n710), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G2084), .Z(new_n749));
  NOR2_X1   g324(.A1(G27), .A2(G29), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G164), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2078), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT30), .B(G28), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n710), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n742), .A2(new_n744), .A3(new_n749), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT98), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n700), .A2(KEYINPUT88), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n699), .A2(new_n702), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n672), .A2(KEYINPUT23), .A3(G20), .ZN(new_n760));
  AOI21_X1  g335(.A(KEYINPUT23), .B1(new_n672), .B2(G20), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n760), .B(new_n761), .C1(G299), .C2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n710), .A2(G26), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT92), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n471), .A2(G140), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n473), .A2(G128), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(G104), .A2(G2105), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n772), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n473), .A2(KEYINPUT90), .A3(G128), .ZN(new_n774));
  AND4_X1   g349(.A1(new_n768), .A2(new_n771), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT91), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(KEYINPUT91), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n767), .B1(new_n778), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G2067), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n764), .B(new_n781), .C1(new_n755), .C2(new_n756), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n703), .A2(new_n757), .A3(new_n759), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n672), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n540), .B2(new_n672), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT89), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1341), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n672), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n589), .B2(new_n672), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n710), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n710), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT29), .B(G2090), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT99), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n783), .A2(new_n787), .A3(new_n792), .A4(new_n798), .ZN(G311));
  INV_X1    g374(.A(new_n783), .ZN(new_n800));
  INV_X1    g375(.A(new_n787), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n800), .A2(new_n801), .A3(new_n791), .A4(new_n797), .ZN(G150));
  AOI22_X1  g377(.A1(new_n497), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(new_n499), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n514), .A2(G93), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT100), .B(G55), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n505), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT102), .B(G860), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT37), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n589), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT39), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n808), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n808), .A2(new_n815), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n540), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n598), .A2(new_n815), .A3(new_n808), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n814), .B(new_n820), .Z(new_n821));
  OAI21_X1  g396(.A(new_n811), .B1(new_n821), .B2(new_n809), .ZN(G145));
  XNOR2_X1  g397(.A(new_n778), .B(G164), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n709), .B(new_n734), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n694), .B(new_n610), .ZN(new_n826));
  OR2_X1    g401(.A1(G106), .A2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n827), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n828));
  INV_X1    g403(.A(G142), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n462), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G130), .B2(new_n473), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n826), .B(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT103), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n825), .A2(new_n832), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n825), .A2(KEYINPUT103), .A3(new_n832), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n607), .B(G160), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G162), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(G37), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n833), .A2(new_n835), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g420(.A1(new_n808), .A2(new_n592), .ZN(new_n846));
  XNOR2_X1  g421(.A(G303), .B(G288), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G305), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G290), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT42), .Z(new_n850));
  OR2_X1    g425(.A1(new_n585), .A2(new_n586), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G651), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n852), .A2(new_n853), .A3(new_n583), .A4(new_n582), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n588), .A2(KEYINPUT104), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n855), .A3(G299), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n588), .A2(G299), .A3(KEYINPUT104), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT41), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n856), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(KEYINPUT105), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n863), .A3(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n820), .B(new_n600), .ZN(new_n866));
  MUX2_X1   g441(.A(new_n858), .B(new_n865), .S(new_n866), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n850), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n846), .B1(new_n868), .B2(new_n592), .ZN(G295));
  OAI21_X1  g444(.A(new_n846), .B1(new_n868), .B2(new_n592), .ZN(G331));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n871));
  NAND2_X1  g446(.A1(G286), .A2(G301), .ZN(new_n872));
  NAND2_X1  g447(.A1(G168), .A2(G171), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n820), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n872), .A2(new_n818), .A3(new_n819), .A4(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n862), .A2(new_n877), .A3(new_n864), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT106), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n877), .A2(new_n858), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n862), .A2(new_n877), .A3(new_n882), .A4(new_n864), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n879), .A2(new_n849), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  INV_X1    g460(.A(new_n849), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n876), .A2(new_n875), .B1(new_n859), .B2(new_n861), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n891), .A2(new_n886), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n884), .A2(new_n885), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT43), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n890), .B1(new_n894), .B2(KEYINPUT107), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n890), .A2(KEYINPUT107), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n871), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT108), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n884), .A2(new_n885), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n891), .A2(new_n886), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(KEYINPUT44), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT109), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n906), .B(new_n871), .C1(new_n895), .C2(new_n896), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n898), .A2(new_n905), .A3(new_n907), .ZN(G397));
  NOR2_X1   g483(.A1(G164), .A2(G1384), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(KEYINPUT110), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(KEYINPUT110), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G160), .A2(G40), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n778), .A2(G2067), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n776), .A2(new_n780), .A3(new_n777), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G1996), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n709), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n694), .B(new_n697), .Z(new_n925));
  AOI21_X1  g500(.A(new_n916), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n916), .A2(G1986), .A3(G290), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT48), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n915), .B1(new_n919), .B2(new_n709), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n916), .B2(G1996), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n915), .A2(KEYINPUT46), .A3(new_n921), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT127), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n935), .B(KEYINPUT47), .Z(new_n936));
  OR2_X1    g511(.A1(new_n694), .A2(new_n697), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n918), .B1(new_n923), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g513(.A(new_n929), .B(new_n936), .C1(new_n915), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT126), .ZN(new_n940));
  INV_X1    g515(.A(G8), .ZN(new_n941));
  NAND2_X1  g516(.A1(G303), .A2(G8), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT55), .ZN(new_n944));
  XNOR2_X1  g519(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n489), .A2(new_n491), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n483), .A2(new_n486), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n952));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G40), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n466), .A2(new_n469), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n948), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n957), .A2(G2090), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT113), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n911), .B1(G164), .B2(G1384), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n951), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n956), .ZN(new_n962));
  INV_X1    g537(.A(G1971), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT112), .Z(new_n965));
  AOI211_X1 g540(.A(new_n941), .B(new_n947), .C1(new_n959), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n909), .A2(new_n956), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(G8), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n968), .B(KEYINPUT115), .Z(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(G1976), .B2(new_n677), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n970), .B(new_n971), .C1(G1976), .C2(new_n677), .ZN(new_n973));
  INV_X1    g548(.A(new_n969), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT116), .B(G86), .Z(new_n975));
  OAI21_X1  g550(.A(new_n569), .B1(new_n508), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G1981), .ZN(new_n977));
  INV_X1    g552(.A(G1981), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n569), .B(new_n978), .C1(new_n570), .C2(new_n508), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(KEYINPUT117), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT49), .B1(new_n980), .B2(KEYINPUT118), .ZN(new_n981));
  NAND2_X1  g556(.A1(KEYINPUT118), .A2(KEYINPUT49), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n977), .A2(new_n979), .B1(KEYINPUT117), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n974), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n972), .A2(new_n973), .A3(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n958), .A2(new_n964), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(new_n941), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n966), .B(new_n985), .C1(new_n947), .C2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n962), .A2(new_n723), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT119), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n957), .A2(G2084), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n962), .A2(new_n992), .A3(new_n723), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT122), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n990), .A2(new_n991), .A3(KEYINPUT122), .A4(new_n993), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(G168), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G8), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT51), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n1001));
  AOI211_X1 g576(.A(KEYINPUT51), .B(new_n941), .C1(new_n1001), .C2(G168), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT123), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n996), .A2(new_n997), .ZN(new_n1006));
  NOR2_X1   g581(.A1(G168), .A2(new_n941), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1007), .ZN(new_n1009));
  AOI211_X1 g584(.A(KEYINPUT123), .B(new_n1009), .C1(new_n996), .C2(new_n997), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n957), .A2(new_n740), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n962), .A2(G2078), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT124), .Z(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1018));
  AOI21_X1  g593(.A(G301), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n962), .A2(new_n992), .A3(new_n723), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n992), .B1(new_n962), .B2(new_n723), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT122), .B1(new_n1022), .B2(new_n991), .ZN(new_n1023));
  INV_X1    g598(.A(new_n997), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1007), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT123), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1006), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1002), .B1(new_n999), .B2(KEYINPUT51), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT62), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1012), .A2(new_n1019), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1033));
  AND4_X1   g608(.A1(G40), .A2(G160), .A3(new_n953), .A4(new_n951), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT58), .B(G1341), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n962), .A2(G1996), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n540), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(KEYINPUT59), .A3(new_n540), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n790), .A2(new_n957), .B1(new_n1034), .B2(new_n780), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(new_n589), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n957), .A2(new_n790), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(G2067), .B2(new_n967), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n589), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1041), .A2(new_n588), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT56), .B(G2072), .Z(new_n1051));
  OR2_X1    g626(.A1(new_n962), .A2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n957), .A2(KEYINPUT120), .A3(new_n763), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT120), .B1(new_n957), .B2(new_n763), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n1056));
  XNOR2_X1  g631(.A(G299), .B(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT61), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1057), .B(new_n1052), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1050), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1047), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT121), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1069), .B(new_n1061), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1064), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1072));
  XNOR2_X1  g647(.A(G301), .B(KEYINPUT54), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G2078), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  OAI21_X1  g651(.A(G40), .B1(new_n466), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1076), .B2(new_n466), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n1015), .B(new_n469), .C1(new_n909), .C2(KEYINPUT45), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n913), .A2(new_n1075), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1073), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1018), .A3(new_n1081), .A4(new_n1013), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1033), .A2(new_n1071), .A3(new_n1074), .A4(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1001), .A2(new_n941), .A3(G286), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT63), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n988), .B1(new_n1032), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n985), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n966), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n981), .A2(new_n983), .ZN(new_n1091));
  OR2_X1    g666(.A1(G288), .A2(G1976), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n979), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n974), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n959), .A2(new_n965), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n946), .B1(new_n1095), .B2(G8), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1084), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n985), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1090), .B(new_n1094), .C1(new_n1098), .C2(new_n1085), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1088), .A2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n916), .A2(new_n686), .A3(new_n576), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n927), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT111), .Z(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(new_n926), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n940), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1012), .A2(new_n1019), .A3(new_n1031), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1099), .B1(new_n1109), .B2(new_n988), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1106), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1110), .A2(KEYINPUT126), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n939), .B1(new_n1107), .B2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g688(.A1(new_n890), .A2(KEYINPUT107), .ZN(new_n1115));
  AND2_X1   g689(.A1(new_n894), .A2(KEYINPUT107), .ZN(new_n1116));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1116), .B2(new_n890), .ZN(new_n1117));
  AOI211_X1 g691(.A(G401), .B(G229), .C1(new_n841), .C2(new_n843), .ZN(new_n1118));
  AND4_X1   g692(.A1(G319), .A2(new_n1117), .A3(new_n645), .A4(new_n1118), .ZN(G308));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(G319), .A4(new_n645), .ZN(G225));
endmodule


