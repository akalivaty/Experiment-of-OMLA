

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586;

  XOR2_X1 U321 ( .A(n425), .B(n424), .Z(n462) );
  XNOR2_X1 U322 ( .A(n447), .B(KEYINPUT122), .ZN(n569) );
  XNOR2_X1 U323 ( .A(n339), .B(KEYINPUT46), .ZN(n359) );
  XNOR2_X1 U324 ( .A(n417), .B(G22GAT), .ZN(n419) );
  XNOR2_X1 U325 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U326 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U327 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n369) );
  XNOR2_X1 U328 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U329 ( .A(n370), .B(n369), .ZN(n549) );
  NOR2_X1 U330 ( .A1(n517), .A2(n481), .ZN(n473) );
  INV_X1 U331 ( .A(G190GAT), .ZN(n448) );
  XNOR2_X1 U332 ( .A(n473), .B(n472), .ZN(n501) );
  XNOR2_X1 U333 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U334 ( .A(n474), .B(KEYINPUT40), .ZN(n475) );
  XNOR2_X1 U335 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XNOR2_X1 U336 ( .A(n476), .B(n475), .ZN(G1330GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n290) );
  NAND2_X1 U338 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U339 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U340 ( .A(n291), .B(KEYINPUT10), .Z(n296) );
  XOR2_X1 U341 ( .A(G43GAT), .B(G50GAT), .Z(n293) );
  XNOR2_X1 U342 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n330) );
  XNOR2_X1 U344 ( .A(G29GAT), .B(G134GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n294), .B(KEYINPUT77), .ZN(n389) );
  XNOR2_X1 U346 ( .A(n330), .B(n389), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U348 ( .A(G92GAT), .B(G106GAT), .Z(n298) );
  XNOR2_X1 U349 ( .A(G162GAT), .B(G218GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U351 ( .A(n300), .B(n299), .Z(n302) );
  XOR2_X1 U352 ( .A(G36GAT), .B(G190GAT), .Z(n371) );
  XOR2_X1 U353 ( .A(G99GAT), .B(G85GAT), .Z(n313) );
  XNOR2_X1 U354 ( .A(n371), .B(n313), .ZN(n301) );
  XOR2_X1 U355 ( .A(n302), .B(n301), .Z(n545) );
  INV_X1 U356 ( .A(n545), .ZN(n559) );
  XOR2_X1 U357 ( .A(KEYINPUT74), .B(G64GAT), .Z(n304) );
  XNOR2_X1 U358 ( .A(G176GAT), .B(G92GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U360 ( .A(G204GAT), .B(n305), .Z(n375) );
  XOR2_X1 U361 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n307) );
  XNOR2_X1 U362 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n375), .B(n308), .ZN(n319) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(G78GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n309), .B(KEYINPUT73), .ZN(n416) );
  XOR2_X1 U367 ( .A(n416), .B(KEYINPUT31), .Z(n311) );
  NAND2_X1 U368 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n317) );
  XNOR2_X1 U370 ( .A(G120GAT), .B(G148GAT), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n312), .B(G57GAT), .ZN(n398) );
  XNOR2_X1 U372 ( .A(n398), .B(n313), .ZN(n315) );
  XOR2_X1 U373 ( .A(G71GAT), .B(KEYINPUT13), .Z(n340) );
  INV_X1 U374 ( .A(n340), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n364) );
  XNOR2_X1 U376 ( .A(KEYINPUT41), .B(n364), .ZN(n504) );
  XOR2_X1 U377 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n321) );
  XNOR2_X1 U378 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n338) );
  XOR2_X1 U380 ( .A(G113GAT), .B(G36GAT), .Z(n323) );
  XNOR2_X1 U381 ( .A(G169GAT), .B(G29GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U383 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n325) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(G197GAT), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U386 ( .A(n327), .B(n326), .Z(n336) );
  XOR2_X1 U387 ( .A(G1GAT), .B(G8GAT), .Z(n329) );
  XNOR2_X1 U388 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n334) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G22GAT), .Z(n350) );
  XOR2_X1 U391 ( .A(n330), .B(n350), .Z(n332) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n532) );
  NAND2_X1 U397 ( .A1(n504), .A2(n532), .ZN(n339) );
  XOR2_X1 U398 ( .A(n340), .B(KEYINPUT12), .Z(n342) );
  NAND2_X1 U399 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U401 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n344) );
  XNOR2_X1 U402 ( .A(KEYINPUT81), .B(KEYINPUT79), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U404 ( .A(n346), .B(n345), .Z(n352) );
  XOR2_X1 U405 ( .A(KEYINPUT82), .B(KEYINPUT15), .Z(n348) );
  XNOR2_X1 U406 ( .A(G57GAT), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U410 ( .A(G8GAT), .B(KEYINPUT78), .Z(n372) );
  XOR2_X1 U411 ( .A(G1GAT), .B(G127GAT), .Z(n395) );
  XOR2_X1 U412 ( .A(n372), .B(n395), .Z(n354) );
  XNOR2_X1 U413 ( .A(G155GAT), .B(G211GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U415 ( .A(n356), .B(n355), .Z(n358) );
  XNOR2_X1 U416 ( .A(G183GAT), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n581) );
  NAND2_X1 U418 ( .A1(n359), .A2(n581), .ZN(n360) );
  NOR2_X1 U419 ( .A1(n559), .A2(n360), .ZN(n362) );
  XNOR2_X1 U420 ( .A(KEYINPUT115), .B(KEYINPUT47), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n545), .B(KEYINPUT36), .ZN(n584) );
  NOR2_X1 U423 ( .A1(n581), .A2(n584), .ZN(n363) );
  XNOR2_X1 U424 ( .A(KEYINPUT45), .B(n363), .ZN(n365) );
  NAND2_X1 U425 ( .A1(n365), .A2(n364), .ZN(n366) );
  NOR2_X1 U426 ( .A1(n532), .A2(n366), .ZN(n367) );
  NOR2_X1 U427 ( .A1(n368), .A2(n367), .ZN(n370) );
  XOR2_X1 U428 ( .A(n372), .B(n371), .Z(n374) );
  NAND2_X1 U429 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U431 ( .A(n376), .B(n375), .Z(n386) );
  XNOR2_X1 U432 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n377), .B(KEYINPUT89), .ZN(n378) );
  XOR2_X1 U434 ( .A(n378), .B(KEYINPUT17), .Z(n380) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(G183GAT), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n441) );
  XOR2_X1 U437 ( .A(KEYINPUT21), .B(G218GAT), .Z(n382) );
  XNOR2_X1 U438 ( .A(KEYINPUT91), .B(G211GAT), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U440 ( .A(G197GAT), .B(n383), .Z(n424) );
  INV_X1 U441 ( .A(n424), .ZN(n384) );
  XOR2_X1 U442 ( .A(n441), .B(n384), .Z(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n523) );
  XNOR2_X1 U444 ( .A(n523), .B(KEYINPUT120), .ZN(n387) );
  NOR2_X1 U445 ( .A1(n549), .A2(n387), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n388), .B(KEYINPUT54), .ZN(n410) );
  XOR2_X1 U447 ( .A(n389), .B(KEYINPUT4), .Z(n391) );
  NAND2_X1 U448 ( .A1(G225GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n409) );
  XOR2_X1 U450 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n393) );
  XNOR2_X1 U451 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n394), .B(KEYINPUT94), .Z(n397) );
  XNOR2_X1 U454 ( .A(n395), .B(G85GAT), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n399) );
  XOR2_X1 U456 ( .A(n399), .B(n398), .Z(n407) );
  XOR2_X1 U457 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n401) );
  XNOR2_X1 U458 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n434) );
  XNOR2_X1 U460 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n402), .B(KEYINPUT3), .ZN(n403) );
  XOR2_X1 U462 ( .A(n403), .B(KEYINPUT92), .Z(n405) );
  XNOR2_X1 U463 ( .A(G141GAT), .B(G162GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n418) );
  XNOR2_X1 U465 ( .A(n434), .B(n418), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n460) );
  XOR2_X1 U468 ( .A(KEYINPUT95), .B(n460), .Z(n550) );
  INV_X1 U469 ( .A(n550), .ZN(n520) );
  NAND2_X1 U470 ( .A1(n410), .A2(n520), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n411), .B(KEYINPUT65), .ZN(n573) );
  XOR2_X1 U472 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n413) );
  XNOR2_X1 U473 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U475 ( .A(G50GAT), .B(G148GAT), .Z(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n421) );
  XOR2_X1 U477 ( .A(KEYINPUT24), .B(n416), .Z(n417) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n423) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n425) );
  NAND2_X1 U481 ( .A1(n573), .A2(n462), .ZN(n427) );
  XOR2_X1 U482 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n446) );
  XOR2_X1 U484 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n429) );
  XNOR2_X1 U485 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U487 ( .A(KEYINPUT88), .B(G99GAT), .Z(n431) );
  XNOR2_X1 U488 ( .A(G15GAT), .B(G190GAT), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n445) );
  XOR2_X1 U491 ( .A(n434), .B(G134GAT), .Z(n436) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U494 ( .A(G71GAT), .B(G120GAT), .Z(n438) );
  XNOR2_X1 U495 ( .A(G176GAT), .B(G127GAT), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U497 ( .A(n440), .B(n439), .Z(n443) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X2 U500 ( .A(n445), .B(n444), .Z(n525) );
  INV_X1 U501 ( .A(n525), .ZN(n535) );
  NAND2_X1 U502 ( .A1(n446), .A2(n535), .ZN(n447) );
  NOR2_X1 U503 ( .A1(n569), .A2(n545), .ZN(n451) );
  XNOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT126), .ZN(n449) );
  NOR2_X1 U505 ( .A1(n523), .A2(n525), .ZN(n452) );
  XNOR2_X1 U506 ( .A(KEYINPUT97), .B(n452), .ZN(n453) );
  NAND2_X1 U507 ( .A1(n453), .A2(n462), .ZN(n456) );
  XOR2_X1 U508 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n454) );
  XNOR2_X1 U509 ( .A(KEYINPUT25), .B(n454), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(n459) );
  XOR2_X1 U511 ( .A(n523), .B(KEYINPUT27), .Z(n464) );
  NOR2_X1 U512 ( .A1(n462), .A2(n535), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n457), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U514 ( .A1(n464), .A2(n572), .ZN(n548) );
  XOR2_X1 U515 ( .A(KEYINPUT96), .B(n548), .Z(n458) );
  NOR2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n467) );
  XOR2_X1 U518 ( .A(n462), .B(KEYINPUT66), .Z(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT28), .B(n463), .Z(n528) );
  AND2_X1 U520 ( .A1(n550), .A2(n464), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n528), .A2(n465), .ZN(n533) );
  NOR2_X1 U522 ( .A1(n533), .A2(n535), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U524 ( .A(KEYINPUT100), .B(n468), .ZN(n479) );
  NOR2_X1 U525 ( .A1(n584), .A2(n479), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n469), .A2(n581), .ZN(n471) );
  INV_X1 U527 ( .A(KEYINPUT37), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(n517) );
  NAND2_X1 U529 ( .A1(n364), .A2(n532), .ZN(n481) );
  INV_X1 U530 ( .A(KEYINPUT38), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n501), .A2(n525), .ZN(n476) );
  INV_X1 U532 ( .A(G43GAT), .ZN(n474) );
  INV_X1 U533 ( .A(G1GAT), .ZN(n487) );
  INV_X1 U534 ( .A(KEYINPUT102), .ZN(n484) );
  NOR2_X1 U535 ( .A1(n559), .A2(n581), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  NOR2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n480) );
  XOR2_X1 U538 ( .A(n480), .B(KEYINPUT101), .Z(n505) );
  INV_X1 U539 ( .A(n481), .ZN(n482) );
  AND2_X1 U540 ( .A1(n505), .A2(n482), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n494) );
  NOR2_X1 U542 ( .A1(n520), .A2(n494), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(n485), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  XNOR2_X1 U545 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n489) );
  NOR2_X1 U546 ( .A1(n523), .A2(n494), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  NOR2_X1 U548 ( .A1(n525), .A2(n494), .ZN(n493) );
  XOR2_X1 U549 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n491) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  INV_X1 U553 ( .A(KEYINPUT106), .ZN(n496) );
  NOR2_X1 U554 ( .A1(n528), .A2(n494), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n497), .ZN(G1327GAT) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  NOR2_X1 U558 ( .A1(n520), .A2(n501), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n523), .A2(n501), .ZN(n500) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n528), .A2(n501), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  XNOR2_X1 U565 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n509) );
  XOR2_X1 U566 ( .A(KEYINPUT108), .B(n504), .Z(n564) );
  NOR2_X1 U567 ( .A1(n532), .A2(n564), .ZN(n518) );
  NAND2_X1 U568 ( .A1(n505), .A2(n518), .ZN(n514) );
  NOR2_X1 U569 ( .A1(n520), .A2(n514), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n523), .A2(n514), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NOR2_X1 U576 ( .A1(n525), .A2(n514), .ZN(n512) );
  XOR2_X1 U577 ( .A(KEYINPUT112), .B(n512), .Z(n513) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  NOR2_X1 U579 ( .A1(n528), .A2(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  INV_X1 U582 ( .A(n517), .ZN(n519) );
  NAND2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n527) );
  NOR2_X1 U584 ( .A1(n520), .A2(n527), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n527), .ZN(n524) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U589 ( .A1(n525), .A2(n527), .ZN(n526) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n530) );
  XNOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT114), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n531), .Z(G1339GAT) );
  INV_X1 U595 ( .A(n532), .ZN(n574) );
  NOR2_X1 U596 ( .A1(n533), .A2(n549), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n544) );
  NOR2_X1 U598 ( .A1(n574), .A2(n544), .ZN(n536) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(n536), .Z(n537) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  NOR2_X1 U601 ( .A1(n544), .A2(n564), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n539) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NOR2_X1 U606 ( .A1(n581), .A2(n544), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(n542), .Z(n543) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n557) );
  NOR2_X1 U614 ( .A1(n574), .A2(n557), .ZN(n553) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  INV_X1 U618 ( .A(n557), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n560), .A2(n504), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n581), .A2(n557), .ZN(n558) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n569), .A2(n574), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(n562), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(KEYINPUT123), .ZN(G1348GAT) );
  XNOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n568) );
  NOR2_X1 U630 ( .A1(n569), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  XNOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n571) );
  NOR2_X1 U635 ( .A1(n581), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1350GAT) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n583) );
  NOR2_X1 U638 ( .A1(n574), .A2(n583), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n364), .A2(n583), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

