//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n446, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT64), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT64), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G217));
  NOR3_X1   g029(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n455));
  NAND3_X1  g030(.A1(new_n437), .A2(new_n438), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AND2_X1   g036(.A1(new_n457), .A2(G2106), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(new_n463), .B1(G567), .B2(new_n459), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(G319));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(G137), .A3(new_n470), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n468), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(KEYINPUT68), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n484), .A3(G125), .ZN(new_n485));
  NAND2_X1  g060(.A1(G113), .A2(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n476), .B1(new_n487), .B2(G2105), .ZN(G160));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n474), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n482), .A2(KEYINPUT70), .A3(new_n483), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n470), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n470), .A2(G112), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n490), .A2(new_n491), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n470), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n497), .A2(new_n500), .A3(new_n470), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n496), .B1(new_n502), .B2(G136), .ZN(G162));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n504), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n480), .A2(new_n484), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g081(.A(G138), .B(new_n470), .C1(new_n478), .C2(new_n479), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(G126), .A2(G2105), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n510), .B1(new_n478), .B2(new_n479), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n470), .A2(G114), .ZN(new_n512));
  OAI21_X1  g087(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(KEYINPUT72), .B1(new_n509), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(G164));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT73), .Z(new_n522));
  OAI21_X1  g097(.A(G651), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(G543), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(G88), .B1(new_n531), .B2(G50), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n537), .B2(new_n530), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n525), .A2(new_n524), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT6), .B(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  INV_X1    g123(.A(G52), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n528), .A2(new_n548), .B1(new_n530), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  NAND3_X1  g126(.A1(new_n519), .A2(new_n540), .A3(G81), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n540), .A2(G43), .A3(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(G56), .B1(new_n525), .B2(new_n524), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n546), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g135(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND3_X1  g139(.A1(new_n540), .A2(G53), .A3(G543), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT75), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n567), .B(KEYINPUT9), .C1(KEYINPUT75), .C2(new_n565), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  OAI211_X1 g144(.A(KEYINPUT75), .B(new_n569), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n546), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n519), .A2(new_n540), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(G91), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n568), .A2(new_n570), .A3(new_n572), .A4(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  OR2_X1    g154(.A1(new_n519), .A2(G74), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G49), .B2(new_n531), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n573), .A2(G87), .A3(new_n575), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n546), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n573), .A2(G86), .A3(new_n575), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n573), .A2(new_n588), .A3(G86), .A4(new_n575), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n531), .A2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  XNOR2_X1  g167(.A(KEYINPUT79), .B(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n528), .A2(new_n593), .B1(new_n530), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n546), .B2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n602), .B(new_n603), .C1(new_n539), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n530), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n573), .A2(G92), .A3(new_n575), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n573), .A2(KEYINPUT10), .A3(G92), .A4(new_n575), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  AND4_X1   g191(.A1(new_n568), .A2(new_n570), .A3(new_n572), .A4(new_n576), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT82), .Z(G148));
  NAND2_X1  g197(.A1(new_n613), .A2(new_n620), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g201(.A1(new_n472), .A2(new_n480), .A3(new_n484), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2100), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n502), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n492), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n470), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n642), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(G14), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n649), .ZN(G401));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n636), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT83), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n669), .A2(new_n670), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n677), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(new_n672), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n678), .C1(new_n668), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT85), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n681), .B(new_n683), .Z(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT84), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n684), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  NAND2_X1  g265(.A1(new_n502), .A2(G131), .ZN(new_n691));
  OAI21_X1  g266(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n692));
  INV_X1    g267(.A(G107), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(G2105), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n492), .A2(G119), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(KEYINPUT86), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n492), .A2(new_n697), .A3(G119), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n694), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT87), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT88), .B(G16), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G24), .B(G290), .S(new_n706), .Z(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G6), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G305), .B2(G16), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  MUX2_X1   g290(.A(G23), .B(G288), .S(G16), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n706), .A2(G22), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n706), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n714), .A2(new_n715), .A3(new_n718), .A4(new_n722), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n704), .B(new_n709), .C1(KEYINPUT34), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(KEYINPUT34), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT89), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G33), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT25), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n480), .A2(new_n484), .A3(G127), .ZN(new_n735));
  INV_X1    g310(.A(G115), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n468), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n734), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n499), .A2(new_n501), .ZN(new_n739));
  INV_X1    g314(.A(G139), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n732), .B1(new_n741), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2072), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT90), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n731), .A2(G35), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT94), .Z(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n731), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n745), .B1(G2090), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n742), .A2(new_n743), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n731), .A2(G27), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(KEYINPUT93), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n753), .B(new_n754), .C1(G164), .C2(new_n731), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2078), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n710), .A2(G5), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G171), .B2(new_n710), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT92), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n502), .A2(G141), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT26), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n472), .A2(G105), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n765), .B(new_n766), .C1(new_n492), .C2(G129), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(new_n731), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n731), .B2(G32), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n757), .B(new_n762), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G28), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT30), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(KEYINPUT30), .ZN(new_n776));
  OR2_X1    g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  NAND2_X1  g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G1341), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n558), .A2(new_n705), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G19), .B2(new_n705), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n779), .B1(new_n780), .B2(new_n782), .C1(new_n635), .C2(new_n731), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G21), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G168), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT91), .B(G1966), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n782), .A2(new_n780), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n731), .B1(new_n789), .B2(G34), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n789), .B2(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G160), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n783), .A2(new_n788), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n755), .A2(G2078), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n770), .B2(new_n771), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n750), .A2(new_n773), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n731), .A2(G26), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT28), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n502), .A2(G140), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G116), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G2105), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n492), .B2(G128), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2067), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n710), .A2(G4), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n613), .B2(new_n710), .ZN(new_n811));
  INV_X1    g386(.A(G1348), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n705), .A2(G20), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT23), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n617), .B2(new_n710), .ZN(new_n816));
  INV_X1    g391(.A(G1956), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n809), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n749), .A2(G2090), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n799), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n730), .A2(new_n824), .ZN(G311));
  NAND2_X1  g400(.A1(new_n730), .A2(new_n824), .ZN(G150));
  NAND3_X1  g401(.A1(new_n519), .A2(new_n540), .A3(G93), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT96), .B(G55), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n540), .A2(new_n828), .A3(G543), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n827), .B(new_n829), .C1(new_n830), .C2(new_n546), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT99), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n613), .A2(G559), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT38), .Z(new_n836));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n827), .A2(new_n829), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n519), .A2(G67), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n546), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n555), .A2(new_n556), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n553), .B(new_n552), .C1(new_n843), .C2(new_n546), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n837), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n558), .A2(new_n831), .A3(KEYINPUT97), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n842), .A2(KEYINPUT98), .A3(new_n844), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n558), .B2(new_n831), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n836), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  INV_X1    g430(.A(G860), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n834), .B1(new_n855), .B2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n635), .B(G160), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(G162), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n509), .A2(new_n515), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT100), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n741), .B(new_n862), .Z(new_n863));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n700), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n691), .A2(new_n699), .A3(KEYINPUT102), .ZN(new_n866));
  INV_X1    g441(.A(new_n628), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n863), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n741), .B(new_n862), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n866), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n628), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  INV_X1    g451(.A(G142), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n739), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n502), .A2(KEYINPUT101), .A3(G142), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  INV_X1    g456(.A(G118), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(G2105), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n492), .B2(G130), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n763), .A2(new_n767), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(new_n807), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n807), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n880), .B(new_n884), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n880), .A2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n807), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n768), .A2(new_n802), .A3(new_n806), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n870), .A2(new_n875), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n873), .A2(new_n871), .A3(new_n874), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n895), .A2(new_n896), .B1(new_n892), .B2(new_n888), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n860), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n893), .B1(new_n870), .B2(new_n875), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n859), .B(G162), .Z(new_n901));
  NAND4_X1  g476(.A1(new_n895), .A2(new_n896), .A3(new_n892), .A4(new_n888), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g480(.A(G305), .B(G290), .ZN(new_n906));
  XOR2_X1   g481(.A(G288), .B(G303), .Z(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n852), .B(new_n623), .ZN(new_n912));
  INV_X1    g487(.A(new_n613), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n617), .A2(new_n613), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n913), .A2(G299), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n617), .A2(new_n613), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT41), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n914), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n918), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT103), .B1(new_n916), .B2(KEYINPUT41), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n917), .B1(new_n926), .B2(new_n912), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n911), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n926), .A2(new_n912), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n910), .B(new_n909), .C1(new_n929), .C2(new_n917), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n928), .B(new_n930), .C1(new_n910), .C2(new_n909), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G868), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n842), .A2(G868), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(G295));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n932), .B2(new_n934), .ZN(new_n937));
  AOI211_X1 g512(.A(KEYINPUT105), .B(new_n933), .C1(new_n931), .C2(G868), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n847), .A2(new_n851), .A3(G301), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G301), .B1(new_n847), .B2(new_n851), .ZN(new_n943));
  OAI21_X1  g518(.A(G286), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n852), .A2(G171), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(G168), .A3(new_n941), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n921), .A2(new_n923), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n950));
  INV_X1    g525(.A(new_n916), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n944), .A2(new_n946), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n954), .B2(new_n908), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n944), .A2(new_n946), .A3(new_n957), .A4(new_n951), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n947), .B1(new_n924), .B2(new_n925), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(KEYINPUT106), .B(new_n947), .C1(new_n924), .C2(new_n925), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n908), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n955), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT43), .B1(new_n964), .B2(new_n965), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n963), .ZN(new_n970));
  INV_X1    g545(.A(new_n959), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n908), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n973), .A3(new_n899), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n940), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n899), .A3(new_n966), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n976), .A2(KEYINPUT43), .B1(new_n955), .B2(new_n969), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n940), .B2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n885), .B(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G2067), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n807), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n861), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n470), .B1(new_n485), .B2(new_n486), .ZN(new_n986));
  INV_X1    g561(.A(G40), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n986), .A2(new_n987), .A3(new_n476), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n700), .A2(new_n703), .ZN(new_n992));
  INV_X1    g567(.A(new_n703), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n691), .A2(new_n699), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(G290), .B(new_n708), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n989), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(G303), .A2(G8), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT110), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(KEYINPUT110), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT111), .Z(new_n1004));
  AND3_X1   g579(.A1(new_n999), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n999), .B2(new_n1002), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(new_n984), .C1(new_n516), .C2(new_n517), .ZN(new_n1009));
  INV_X1    g584(.A(G2090), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n514), .B1(new_n506), .B2(new_n508), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(G1384), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1009), .A2(new_n1010), .A3(new_n988), .A4(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n988), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n984), .B1(new_n516), .B2(new_n517), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1014), .B1(new_n1019), .B2(G1971), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT112), .B(G8), .Z(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1007), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1012), .A2(new_n1017), .A3(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n487), .A2(G2105), .ZN(new_n1027));
  INV_X1    g602(.A(new_n476), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(G40), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT72), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n861), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1012), .A2(KEYINPUT72), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n1034), .B2(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n721), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1012), .A2(G1384), .A3(new_n1011), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(new_n1029), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n1010), .C1(new_n1034), .C2(new_n1008), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1025), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1023), .A2(new_n1024), .B1(new_n1040), .B2(new_n1007), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G288), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n509), .B2(new_n515), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1046), .B(new_n1021), .C1(new_n988), .C2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(G160), .A3(G40), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT113), .B1(new_n1049), .B2(new_n1022), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1044), .B(new_n1045), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n861), .A2(new_n984), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1022), .B1(new_n1029), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1046), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(KEYINPUT113), .A3(new_n1022), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1043), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1051), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  INV_X1    g635(.A(new_n591), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(G86), .B2(new_n529), .ZN(new_n1062));
  INV_X1    g637(.A(new_n585), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n587), .A2(new_n589), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1061), .A2(G1981), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT114), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n590), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1070));
  AOI211_X1 g645(.A(new_n1059), .B(new_n1064), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1064), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1070), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1069), .B1(new_n590), .B2(new_n1066), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n1077), .B2(new_n1059), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1058), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1018), .A2(new_n1017), .ZN(new_n1080));
  AOI21_X1  g655(.A(G1971), .B1(new_n1080), .B2(new_n1030), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1008), .A2(new_n984), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1013), .A2(new_n988), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1083), .A2(new_n1084), .A3(G2090), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1022), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1007), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT116), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n985), .A2(new_n1029), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT45), .B(new_n984), .C1(new_n516), .C2(new_n517), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1038), .B(new_n793), .C1(new_n1034), .C2(new_n1008), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1022), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(G286), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1041), .A2(new_n1079), .A3(new_n1089), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT63), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT52), .B1(new_n1073), .B2(new_n1043), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1064), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(KEYINPUT49), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1051), .B(new_n1103), .C1(new_n1106), .C2(new_n1071), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1040), .A2(new_n1007), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1078), .A2(new_n1072), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n988), .B1(new_n1052), .B2(new_n1011), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(KEYINPUT50), .B2(new_n1018), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1010), .A2(new_n1112), .B1(new_n1035), .B2(new_n721), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1087), .B1(new_n1113), .B2(new_n1025), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1058), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1110), .A2(new_n1114), .A3(new_n1115), .A4(KEYINPUT117), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1096), .A2(KEYINPUT63), .A3(G168), .A4(new_n1022), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1007), .B2(new_n1040), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1109), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1101), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1040), .A2(new_n1007), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1107), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G288), .A2(G1976), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1106), .B2(new_n1071), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1073), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(KEYINPUT115), .A3(new_n1125), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1122), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1086), .A2(new_n1024), .A3(new_n1087), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1121), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1024), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1132), .A2(new_n1107), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G168), .A2(new_n1021), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(KEYINPUT51), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1097), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1025), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT51), .B1(new_n1138), .B2(new_n1135), .ZN(new_n1139));
  AOI211_X1 g714(.A(G168), .B(new_n1021), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1137), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G2078), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1030), .B(new_n1144), .C1(new_n1034), .C2(KEYINPUT45), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(G2078), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1090), .A2(new_n1091), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1038), .B1(new_n1034), .B2(new_n1008), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n761), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(KEYINPUT62), .B(new_n1137), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1134), .A2(new_n1143), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1120), .A2(new_n1130), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n817), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT118), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1161), .B(new_n817), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n617), .B(KEYINPUT57), .ZN(new_n1164));
  XNOR2_X1  g739(.A(KEYINPUT56), .B(G2072), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1019), .A2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1164), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1158), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1160), .A2(new_n1162), .B1(new_n1019), .B2(new_n1165), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT119), .B1(new_n1174), .B2(new_n1164), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1164), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1173), .A2(KEYINPUT61), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT59), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1080), .A2(new_n979), .A3(new_n1030), .ZN(new_n1179));
  XOR2_X1   g754(.A(KEYINPUT58), .B(G1341), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n1049), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1178), .B1(new_n1182), .B2(new_n558), .ZN(new_n1183));
  AOI211_X1 g758(.A(KEYINPUT59), .B(new_n844), .C1(new_n1179), .C2(new_n1181), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1049), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n981), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n613), .B2(KEYINPUT121), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1186), .B(new_n1188), .C1(new_n1112), .C2(G1348), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n613), .A2(KEYINPUT121), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1183), .A2(new_n1184), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1150), .A2(new_n812), .B1(new_n981), .B2(new_n1185), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1193), .A2(KEYINPUT60), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g771(.A(KEYINPUT120), .B(new_n1158), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1171), .A2(new_n1177), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1173), .B(new_n1175), .C1(new_n913), .C2(new_n1193), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1176), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1090), .A2(new_n1015), .A3(new_n1148), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1147), .A2(G301), .A3(new_n1151), .A4(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(KEYINPUT54), .B1(new_n1153), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1204), .A2(KEYINPUT122), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n1206));
  AOI211_X1 g781(.A(new_n1206), .B(KEYINPUT54), .C1(new_n1153), .C2(new_n1203), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT51), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1096), .A2(G8), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1135), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1140), .ZN(new_n1213));
  AOI22_X1  g788(.A1(new_n1212), .A2(new_n1213), .B1(new_n1097), .B2(new_n1136), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1107), .A2(new_n1133), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1147), .A2(new_n1151), .A3(new_n1202), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(G171), .ZN(new_n1217));
  OAI211_X1 g792(.A(new_n1217), .B(KEYINPUT54), .C1(G171), .C2(new_n1152), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1214), .A2(new_n1215), .A3(new_n1218), .A4(new_n1041), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1208), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1201), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n998), .B1(new_n1157), .B2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n807), .A2(G2067), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n701), .A2(new_n993), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1223), .B1(new_n991), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n1226));
  OR2_X1    g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n989), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1228));
  AND2_X1   g803(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g804(.A1(G290), .A2(new_n989), .A3(G1986), .ZN(new_n1230));
  XOR2_X1   g805(.A(new_n1230), .B(KEYINPUT48), .Z(new_n1231));
  AND2_X1   g806(.A1(new_n996), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT46), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1233), .B1(new_n989), .B2(G1996), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n990), .A2(KEYINPUT46), .A3(new_n979), .ZN(new_n1235));
  AND2_X1   g810(.A1(new_n982), .A2(new_n768), .ZN(new_n1236));
  OAI211_X1 g811(.A(new_n1234), .B(new_n1235), .C1(new_n1236), .C2(new_n989), .ZN(new_n1237));
  XOR2_X1   g812(.A(KEYINPUT124), .B(KEYINPUT47), .Z(new_n1238));
  XNOR2_X1  g813(.A(new_n1237), .B(new_n1238), .ZN(new_n1239));
  NOR3_X1   g814(.A1(new_n1229), .A2(new_n1232), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1240), .ZN(new_n1241));
  OAI21_X1  g816(.A(KEYINPUT125), .B1(new_n1222), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1243));
  NAND3_X1  g818(.A1(new_n1120), .A2(new_n1130), .A3(new_n1156), .ZN(new_n1244));
  AOI21_X1  g819(.A(new_n1244), .B1(new_n1201), .B2(new_n1220), .ZN(new_n1245));
  OAI211_X1 g820(.A(new_n1243), .B(new_n1240), .C1(new_n1245), .C2(new_n998), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1242), .A2(new_n1246), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g822(.A(new_n899), .B1(new_n964), .B2(new_n965), .ZN(new_n1249));
  AOI211_X1 g823(.A(new_n908), .B(new_n959), .C1(new_n962), .C2(new_n963), .ZN(new_n1250));
  OAI21_X1  g824(.A(KEYINPUT43), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g825(.A1(new_n969), .A2(new_n955), .ZN(new_n1252));
  NAND2_X1  g826(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g827(.A1(G319), .A2(new_n665), .ZN(new_n1254));
  OR3_X1    g828(.A1(G401), .A2(new_n1254), .A3(KEYINPUT126), .ZN(new_n1255));
  OAI21_X1  g829(.A(KEYINPUT126), .B1(G401), .B2(new_n1254), .ZN(new_n1256));
  AND3_X1   g830(.A1(new_n689), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g831(.A1(new_n904), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g832(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g833(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1261));
  AOI211_X1 g835(.A(new_n1261), .B(new_n1258), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1262));
  NOR2_X1   g836(.A1(new_n1260), .A2(new_n1262), .ZN(G308));
  OAI21_X1  g837(.A(new_n1261), .B1(new_n977), .B2(new_n1258), .ZN(new_n1264));
  NAND3_X1  g838(.A1(new_n1253), .A2(KEYINPUT127), .A3(new_n1259), .ZN(new_n1265));
  NAND2_X1  g839(.A1(new_n1264), .A2(new_n1265), .ZN(G225));
endmodule


