//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1111, new_n1112,
    new_n1113;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  INV_X1    g033(.A(new_n451), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n474), .A2(new_n475), .A3(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(G2105), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n474), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G137), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n481), .A2(G136), .ZN(new_n485));
  INV_X1    g060(.A(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n486), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  AND2_X1   g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n479), .A2(new_n486), .A3(new_n474), .A4(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n474), .A2(new_n475), .A3(G138), .A4(new_n486), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n479), .A2(new_n474), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n486), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT69), .Z(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(new_n507), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  INV_X1    g091(.A(new_n514), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n511), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n509), .A2(G51), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n507), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n517), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n509), .A2(G52), .ZN(new_n533));
  INV_X1    g108(.A(new_n515), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n519), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(new_n509), .A2(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n519), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n509), .A2(G53), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT70), .B(KEYINPUT9), .Z(new_n552));
  OR3_X1    g127(.A1(new_n551), .A2(KEYINPUT71), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT71), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n515), .A2(G91), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n519), .C2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  XOR2_X1   g135(.A(new_n531), .B(KEYINPUT72), .Z(G286));
  NAND2_X1  g136(.A1(new_n515), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n509), .A2(G49), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  AOI22_X1  g140(.A1(new_n515), .A2(G86), .B1(new_n509), .B2(G48), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n519), .B2(new_n567), .ZN(G305));
  AND2_X1   g143(.A1(new_n517), .A2(G60), .ZN(new_n569));
  AND2_X1   g144(.A1(G72), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(KEYINPUT73), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(KEYINPUT73), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n515), .A2(G85), .B1(new_n509), .B2(G47), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n515), .A2(G92), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT10), .Z(new_n578));
  NOR2_X1   g153(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n579));
  INV_X1    g154(.A(G54), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n514), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n581), .A2(new_n582), .B1(G651), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n576), .B1(new_n587), .B2(G868), .ZN(G284));
  OAI21_X1  g163(.A(new_n576), .B1(new_n587), .B2(G868), .ZN(G321));
  MUX2_X1   g164(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g165(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g166(.A(KEYINPUT75), .B(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n587), .B1(G860), .B2(new_n592), .ZN(G148));
  NAND2_X1  g168(.A1(new_n587), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g172(.A1(new_n474), .A2(new_n475), .ZN(new_n598));
  NOR3_X1   g173(.A1(new_n467), .A2(G2105), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT12), .Z(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT13), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(G2100), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n481), .A2(G135), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n487), .A2(G123), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n486), .A2(G111), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(G2096), .Z(new_n608));
  NAND2_X1  g183(.A1(new_n602), .A2(new_n608), .ZN(G156));
  INV_X1    g184(.A(KEYINPUT14), .ZN(new_n610));
  XNOR2_X1  g185(.A(G2427), .B(G2438), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(G2430), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT15), .B(G2435), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(new_n612), .ZN(new_n615));
  XNOR2_X1  g190(.A(G2451), .B(G2454), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT16), .ZN(new_n617));
  XNOR2_X1  g192(.A(G1341), .B(G1348), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n615), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2443), .B(G2446), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n622), .A2(G14), .A3(new_n623), .ZN(G401));
  INV_X1    g199(.A(KEYINPUT18), .ZN(new_n625));
  XOR2_X1   g200(.A(G2084), .B(G2090), .Z(new_n626));
  XNOR2_X1  g201(.A(G2067), .B(G2678), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT17), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  XOR2_X1   g207(.A(G2072), .B(G2078), .Z(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n628), .B2(KEYINPUT18), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2096), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(G227));
  XOR2_X1   g211(.A(G1971), .B(G1976), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT19), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1956), .B(G2474), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1961), .B(G1966), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NOR3_X1   g217(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n641), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT20), .Z(new_n645));
  AOI211_X1 g220(.A(new_n643), .B(new_n645), .C1(new_n638), .C2(new_n642), .ZN(new_n646));
  XOR2_X1   g221(.A(G1981), .B(G1986), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT76), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1991), .B(G1996), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G229));
  INV_X1    g228(.A(G29), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(G33), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n481), .A2(G139), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n486), .A2(G103), .A3(G2104), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT25), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT83), .Z(new_n660));
  NAND2_X1  g235(.A1(G115), .A2(G2104), .ZN(new_n661));
  INV_X1    g236(.A(G127), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n598), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(G2105), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n655), .B1(new_n664), .B2(new_n654), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(G2072), .Z(new_n666));
  INV_X1    g241(.A(G16), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G20), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT23), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(G299), .B2(G16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1956), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n531), .A2(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(G21), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G1966), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT31), .B(G11), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT89), .B(G28), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(KEYINPUT30), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(new_n654), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n677), .B(new_n678), .C1(new_n680), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n667), .A2(G5), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G171), .B2(new_n667), .ZN(new_n685));
  INV_X1    g260(.A(G1961), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  OAI221_X1 g262(.A(new_n687), .B1(new_n654), .B2(new_n607), .C1(new_n676), .C2(new_n675), .ZN(new_n688));
  INV_X1    g263(.A(G2084), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT84), .B(KEYINPUT24), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G34), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(new_n654), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n483), .B2(new_n654), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n683), .B(new_n688), .C1(new_n689), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n654), .A2(G35), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G162), .B2(new_n654), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT29), .ZN(new_n697));
  INV_X1    g272(.A(G2090), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n693), .A2(new_n689), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT85), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n654), .A2(G27), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G164), .B2(new_n654), .ZN(new_n703));
  INV_X1    g278(.A(G2078), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n694), .A2(new_n699), .A3(new_n701), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n587), .A2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G4), .B2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G1348), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n667), .A2(G19), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n545), .B2(new_n667), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1341), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n481), .A2(G140), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n487), .A2(G128), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n486), .A2(G116), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT81), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n654), .A2(G26), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G2067), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n714), .B(new_n726), .C1(new_n709), .C2(new_n708), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n672), .B(new_n706), .C1(KEYINPUT82), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n487), .A2(G129), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT86), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n481), .A2(G141), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n468), .A2(G105), .ZN(new_n735));
  AND4_X1   g310(.A1(new_n730), .A2(new_n731), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G32), .B(new_n738), .S(G29), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT27), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1996), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n728), .B(new_n741), .C1(KEYINPUT82), .C2(new_n727), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT90), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n667), .A2(G22), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G166), .B2(new_n667), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT79), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G1971), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n667), .A2(G23), .ZN(new_n748));
  INV_X1    g323(.A(G288), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n667), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT33), .ZN(new_n751));
  INV_X1    g326(.A(G1976), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G6), .B(G305), .S(G16), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT78), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT32), .B(G1981), .Z(new_n756));
  XOR2_X1   g331(.A(new_n755), .B(new_n756), .Z(new_n757));
  NOR3_X1   g332(.A1(new_n747), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT34), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n481), .A2(G131), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n487), .A2(G119), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n486), .A2(G107), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G25), .B(new_n766), .S(G29), .Z(new_n767));
  XOR2_X1   g342(.A(KEYINPUT35), .B(G1991), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G24), .B(G290), .S(G16), .Z(new_n770));
  XOR2_X1   g345(.A(KEYINPUT77), .B(G1986), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n760), .A2(new_n761), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT80), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT80), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n774), .A2(KEYINPUT36), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(KEYINPUT36), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n743), .A2(new_n776), .A3(new_n777), .ZN(G150));
  INV_X1    g353(.A(G150), .ZN(G311));
  AOI22_X1  g354(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n519), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT91), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n515), .A2(G93), .B1(new_n509), .B2(G55), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(KEYINPUT91), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G860), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT37), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n545), .B(KEYINPUT92), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(new_n785), .Z(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT38), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n587), .A2(G559), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n790), .B(new_n791), .Z(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT39), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT93), .ZN(new_n795));
  INV_X1    g370(.A(G860), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n793), .B2(KEYINPUT39), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n787), .B1(new_n795), .B2(new_n797), .ZN(G145));
  INV_X1    g373(.A(KEYINPUT40), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n503), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n500), .A2(KEYINPUT94), .A3(new_n502), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n802), .A2(new_n497), .A3(new_n494), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n719), .B(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n736), .B(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(new_n664), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n737), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n737), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n808), .A2(new_n664), .A3(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(new_n800), .B(new_n807), .S(new_n810), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n481), .A2(G142), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n487), .A2(G130), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n486), .A2(G118), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n811), .B(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n766), .B(KEYINPUT96), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(new_n600), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n483), .B(new_n607), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n491), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n811), .A2(new_n816), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n811), .A2(new_n816), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n819), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n821), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G37), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n823), .B1(new_n821), .B2(new_n826), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n799), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n830), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n832), .A2(KEYINPUT40), .A3(new_n828), .A4(new_n827), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(G395));
  XOR2_X1   g409(.A(new_n594), .B(KEYINPUT97), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n789), .ZN(new_n836));
  OR2_X1    g411(.A1(G299), .A2(new_n587), .ZN(new_n837));
  NAND2_X1  g412(.A1(G299), .A2(new_n587), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT98), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n837), .B(KEYINPUT99), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT41), .B1(new_n842), .B2(new_n838), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G299), .B2(new_n587), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n843), .B1(new_n837), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n841), .B1(new_n846), .B2(new_n836), .ZN(new_n847));
  XNOR2_X1  g422(.A(G305), .B(KEYINPUT100), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G303), .ZN(new_n849));
  XNOR2_X1  g424(.A(G290), .B(new_n749), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(KEYINPUT101), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT42), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n847), .B(new_n854), .ZN(new_n855));
  MUX2_X1   g430(.A(new_n785), .B(new_n855), .S(G868), .Z(G295));
  MUX2_X1   g431(.A(new_n785), .B(new_n855), .S(G868), .Z(G331));
  NOR2_X1   g432(.A1(G171), .A2(G168), .ZN(new_n858));
  INV_X1    g433(.A(G286), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(G171), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n789), .B(new_n860), .Z(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n839), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n851), .A2(new_n852), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n863), .B(new_n864), .C1(new_n846), .C2(new_n862), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(new_n828), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n864), .B(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n842), .A2(new_n845), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n839), .A2(new_n844), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n861), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n867), .B(new_n870), .C1(new_n840), .C2(new_n861), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n866), .A2(KEYINPUT43), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n863), .B1(new_n846), .B2(new_n862), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n867), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT43), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT44), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n866), .A2(new_n877), .A3(new_n871), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n866), .B2(new_n874), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n876), .B1(new_n880), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g456(.A(KEYINPUT125), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n482), .A2(G40), .A3(new_n469), .A4(new_n477), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n478), .A2(KEYINPUT104), .A3(G40), .A4(new_n482), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(G164), .A2(G1384), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT50), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n500), .A2(KEYINPUT94), .A3(new_n502), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT94), .B1(new_n500), .B2(new_n502), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(new_n893), .A3(new_n498), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT106), .B1(new_n894), .B2(G1384), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  INV_X1    g471(.A(G1384), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n804), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n889), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(G2084), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT45), .B1(new_n895), .B2(new_n898), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT112), .B1(new_n902), .B2(new_n887), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n894), .A2(KEYINPUT106), .A3(G1384), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n896), .B1(new_n804), .B2(new_n897), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT112), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n885), .A2(new_n886), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n888), .ZN(new_n911));
  XNOR2_X1  g486(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n903), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n901), .B1(new_n915), .B2(new_n676), .ZN(new_n916));
  INV_X1    g491(.A(G8), .ZN(new_n917));
  NOR2_X1   g492(.A1(G168), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n920), .B(KEYINPUT121), .Z(new_n921));
  NOR2_X1   g496(.A1(new_n916), .A2(new_n917), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n922), .A2(KEYINPUT51), .A3(new_n918), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT122), .B1(new_n916), .B2(new_n917), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT122), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n895), .A2(new_n898), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n887), .B1(new_n926), .B2(new_n904), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n913), .B1(new_n927), .B2(new_n908), .ZN(new_n928));
  AOI21_X1  g503(.A(G1966), .B1(new_n928), .B2(new_n903), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n925), .B(G8), .C1(new_n929), .C2(new_n901), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n918), .B(KEYINPUT123), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n924), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT51), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT124), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n923), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(KEYINPUT124), .A3(KEYINPUT51), .ZN(new_n936));
  AOI211_X1 g511(.A(new_n882), .B(new_n921), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n934), .ZN(new_n938));
  INV_X1    g513(.A(new_n923), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n921), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT125), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT62), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n932), .A2(KEYINPUT124), .A3(KEYINPUT51), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT124), .B1(new_n932), .B2(KEYINPUT51), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n944), .A2(new_n945), .A3(new_n923), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n882), .B1(new_n946), .B2(new_n921), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT62), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n940), .A2(KEYINPUT125), .A3(new_n941), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n909), .A2(new_n895), .A3(new_n898), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(G8), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT52), .B1(G288), .B2(new_n752), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n953), .B(new_n954), .C1(new_n752), .C2(G288), .ZN(new_n955));
  NOR2_X1   g530(.A1(G288), .A2(new_n752), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT52), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(G305), .B(G1981), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT109), .B1(new_n959), .B2(KEYINPUT108), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(KEYINPUT49), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n960), .A2(KEYINPUT49), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n955), .B(new_n957), .C1(new_n965), .C2(new_n952), .ZN(new_n966));
  NAND2_X1  g541(.A1(G303), .A2(G8), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT55), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT107), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n804), .A2(KEYINPUT45), .A3(new_n897), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n911), .A2(new_n912), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n909), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n972), .A2(G1971), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n891), .A2(new_n698), .A3(new_n899), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n917), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n911), .A2(KEYINPUT50), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n978), .B(new_n887), .C1(new_n926), .C2(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n698), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n973), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n917), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n982), .B2(new_n981), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n966), .B(new_n977), .C1(new_n984), .C2(new_n968), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT53), .B1(new_n972), .B2(new_n704), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n686), .B2(new_n900), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n704), .A2(KEYINPUT53), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n928), .A2(new_n903), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(G301), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n943), .A2(new_n950), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n966), .B(KEYINPUT110), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n965), .A2(new_n752), .A3(new_n749), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G1981), .B2(G305), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n993), .A2(new_n977), .B1(new_n953), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n922), .A2(new_n859), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT63), .B1(new_n985), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n968), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n975), .A2(new_n1000), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n1001), .A2(new_n976), .A3(KEYINPUT63), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n993), .A2(new_n1002), .A3(new_n998), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n996), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n947), .A2(new_n949), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n912), .B1(new_n894), .B2(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(new_n883), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(new_n970), .A3(new_n1008), .A4(new_n988), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT126), .Z(new_n1010));
  NAND2_X1  g585(.A1(new_n987), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(G171), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1006), .B1(new_n1012), .B2(new_n990), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(G171), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n987), .A2(G301), .A3(new_n989), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(KEYINPUT54), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n985), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n1018));
  AND3_X1   g593(.A1(G299), .A2(new_n1018), .A3(KEYINPUT57), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(KEYINPUT57), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(KEYINPUT57), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(G299), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT56), .B(G2072), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n972), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(G1956), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1024), .B(new_n1026), .C1(new_n979), .C2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n951), .A2(G2067), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1348), .B1(new_n891), .B2(new_n899), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n587), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT115), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n979), .A2(new_n1027), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1026), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1024), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1026), .B(KEYINPUT116), .C1(new_n979), .C2(new_n1027), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1028), .B1(new_n1034), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(KEYINPUT61), .A3(new_n1028), .ZN(new_n1044));
  INV_X1    g619(.A(G1996), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n972), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT58), .B(G1341), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n951), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n545), .A2(KEYINPUT117), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT118), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1053), .A3(new_n1050), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1058), .A2(new_n1059), .A3(new_n587), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1032), .B1(new_n1031), .B2(KEYINPUT60), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1052), .A2(KEYINPUT59), .A3(new_n1054), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1044), .A2(new_n1057), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1039), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1028), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g645(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n1067), .C2(new_n1028), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1043), .B1(new_n1065), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT120), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(new_n1043), .C1(new_n1065), .C2(new_n1072), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1017), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1004), .B1(new_n1005), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n992), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n887), .A2(new_n1007), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1045), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n738), .A2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1082), .B(KEYINPUT105), .Z(new_n1083));
  XNOR2_X1  g658(.A(new_n719), .B(new_n725), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n736), .B2(new_n1045), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1080), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n768), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n766), .B(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1087), .B1(new_n1080), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(G290), .B(G1986), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1080), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1079), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT46), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1081), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT127), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n736), .B(new_n1084), .C1(new_n1095), .C2(G1996), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1080), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(new_n1100), .B(KEYINPUT47), .Z(new_n1101));
  OR3_X1    g676(.A1(new_n1087), .A2(new_n1088), .A3(new_n766), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n719), .A2(G2067), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n887), .B(new_n1007), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G290), .A2(G1986), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1080), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT48), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1101), .B(new_n1104), .C1(new_n1090), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1094), .A2(new_n1108), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g684(.A1(new_n829), .A2(new_n830), .ZN(new_n1111));
  NOR4_X1   g685(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1112));
  OAI21_X1  g686(.A(new_n1112), .B1(new_n878), .B2(new_n879), .ZN(new_n1113));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1113), .ZN(G308));
  OR2_X1    g688(.A1(new_n1111), .A2(new_n1113), .ZN(G225));
endmodule


