//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT2), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G113), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n196), .ZN(new_n198));
  XNOR2_X1  g012(.A(G116), .B(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n197), .A2(new_n200), .A3(KEYINPUT68), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G134), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT67), .B1(new_n209), .B2(G137), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n207), .A2(G134), .ZN(new_n211));
  OAI211_X1 g025(.A(G131), .B(new_n208), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n209), .B2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(G137), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g036(.A(G128), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G143), .ZN(new_n226));
  AOI21_X1  g040(.A(G146), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n223), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n226), .A3(G146), .ZN(new_n231));
  INV_X1    g045(.A(new_n221), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n222), .A3(G128), .A4(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n219), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n205), .A2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n226), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n229), .B1(new_n238), .B2(new_n228), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n237), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT66), .A2(G131), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n235), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n204), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT68), .B1(new_n197), .B2(new_n200), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n243), .A2(KEYINPUT65), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n241), .B1(new_n227), .B2(new_n229), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(new_n237), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n244), .A2(KEYINPUT66), .A3(G131), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n214), .A2(new_n215), .A3(new_n217), .A4(new_n245), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n253), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n230), .A2(new_n233), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n218), .A3(new_n212), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n252), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n246), .B2(new_n243), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n254), .A4(new_n237), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n265), .A2(new_n252), .A3(new_n266), .A4(new_n262), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n235), .A2(KEYINPUT71), .A3(new_n265), .A4(new_n266), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n249), .B1(new_n271), .B2(new_n248), .ZN(new_n272));
  OR2_X1    g086(.A1(KEYINPUT72), .A2(G237), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT72), .A2(G237), .ZN(new_n274));
  AOI21_X1  g088(.A(G953), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G210), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT27), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G101), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n187), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n254), .A2(new_n255), .A3(new_n237), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n255), .B1(new_n254), .B2(new_n237), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n283), .A2(new_n284), .A3(new_n246), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n285), .B2(new_n234), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n265), .A2(KEYINPUT30), .A3(new_n266), .A4(new_n262), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n205), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n269), .A2(new_n270), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n243), .A2(KEYINPUT65), .B1(new_n257), .B2(new_n258), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n234), .B1(new_n291), .B2(new_n256), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n287), .B(new_n205), .C1(new_n292), .C2(KEYINPUT30), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n281), .B1(new_n280), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n265), .A2(new_n262), .A3(new_n266), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n269), .A2(new_n270), .B1(new_n205), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n249), .B1(new_n300), .B2(new_n248), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n279), .A2(KEYINPUT29), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G472), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n272), .A2(new_n280), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n272), .A2(KEYINPUT73), .A3(new_n280), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n295), .A2(new_n279), .A3(new_n288), .A4(new_n289), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT31), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  AOI211_X1 g128(.A(KEYINPUT32), .B(new_n306), .C1(new_n311), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT32), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(KEYINPUT31), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n290), .A2(new_n313), .A3(new_n279), .A4(new_n295), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n272), .A2(KEYINPUT73), .A3(new_n280), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT73), .B1(new_n272), .B2(new_n280), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n316), .B1(new_n321), .B2(new_n305), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n304), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(G475), .A2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G113), .B(G122), .ZN(new_n328));
  INV_X1    g142(.A(G104), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n275), .A2(G143), .A3(G214), .ZN(new_n331));
  INV_X1    g145(.A(G953), .ZN(new_n332));
  AND2_X1   g146(.A1(KEYINPUT72), .A2(G237), .ZN(new_n333));
  NOR2_X1   g147(.A1(KEYINPUT72), .A2(G237), .ZN(new_n334));
  OAI211_X1 g148(.A(G214), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n224), .A2(new_n226), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n216), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G125), .B(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n228), .ZN(new_n340));
  NOR2_X1   g154(.A1(G125), .A2(G140), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n341), .B1(new_n346), .B2(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G146), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n338), .A2(KEYINPUT18), .B1(new_n340), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT18), .A2(G131), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n350), .B(KEYINPUT83), .Z(new_n351));
  NAND3_X1  g165(.A1(new_n331), .A2(new_n337), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n352), .A2(new_n353), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT16), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n344), .A2(G125), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n359));
  OAI21_X1  g173(.A(G140), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n341), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G140), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n346), .A2(new_n357), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n228), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(G146), .B(new_n364), .C1(new_n347), .C2(new_n357), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(KEYINPUT77), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(new_n228), .C1(new_n362), .C2(new_n365), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n338), .A2(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n331), .A2(new_n337), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G131), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n331), .A2(new_n337), .A3(new_n216), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n372), .B1(new_n376), .B2(KEYINPUT17), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n330), .B(new_n356), .C1(new_n371), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n347), .A2(KEYINPUT19), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT19), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n339), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n228), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n367), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n356), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n330), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI211_X1 g200(.A(KEYINPUT20), .B(new_n327), .C1(new_n378), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n378), .A2(new_n386), .A3(KEYINPUT85), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT85), .B1(new_n378), .B2(new_n386), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n389), .A2(new_n390), .A3(new_n327), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G475), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n356), .B1(new_n371), .B2(new_n377), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n385), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n378), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n397), .B2(new_n298), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n393), .A2(KEYINPUT86), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT86), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n378), .A2(new_n386), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n378), .A2(new_n386), .A3(KEYINPUT85), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n326), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n387), .B1(new_n406), .B2(KEYINPUT20), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n401), .B1(new_n407), .B2(new_n398), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  OAI21_X1  g224(.A(G128), .B1(new_n227), .B2(new_n222), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n231), .A2(new_n232), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n413), .A2(new_n233), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n415));
  XNOR2_X1  g229(.A(G104), .B(G107), .ZN(new_n416));
  INV_X1    g230(.A(G101), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G107), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G104), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n329), .A2(G107), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT80), .A3(G101), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT3), .B1(new_n329), .B2(G107), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n419), .A3(G104), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n424), .A2(new_n426), .A3(new_n417), .A4(new_n421), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n410), .B1(new_n414), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n424), .A2(new_n426), .A3(new_n421), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G101), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT4), .A3(new_n427), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n433), .A3(G101), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n435), .A2(new_n243), .ZN(new_n436));
  INV_X1    g250(.A(new_n428), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n261), .A3(KEYINPUT10), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n429), .A2(new_n246), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(new_n261), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n428), .B1(new_n413), .B2(new_n233), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n259), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G140), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT79), .ZN(new_n446));
  INV_X1    g260(.A(G227), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(G953), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n446), .B(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n259), .B(new_n450), .C1(new_n440), .C2(new_n441), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n439), .A2(new_n444), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n438), .B1(new_n435), .B2(new_n243), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n441), .A2(KEYINPUT10), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n259), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n439), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n452), .B1(new_n456), .B2(new_n449), .ZN(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n298), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(new_n298), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n449), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n439), .A2(new_n451), .A3(new_n444), .ZN(new_n463));
  INV_X1    g277(.A(new_n449), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(G469), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n459), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT9), .B(G234), .ZN(new_n468));
  OAI21_X1  g282(.A(G221), .B1(new_n468), .B2(G902), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n332), .A2(G952), .ZN(new_n471));
  NAND2_X1  g285(.A1(G234), .A2(G237), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT21), .B(G898), .Z(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(G902), .A3(G953), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G214), .B1(G237), .B2(G902), .ZN(new_n477));
  XOR2_X1   g291(.A(new_n477), .B(KEYINPUT82), .Z(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G122), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT8), .Z(new_n481));
  NAND2_X1  g295(.A1(new_n199), .A2(KEYINPUT5), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n482), .B(G113), .C1(KEYINPUT5), .C2(new_n189), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n437), .A2(new_n200), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n200), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n428), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n481), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n261), .A2(new_n343), .A3(new_n345), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n254), .A2(new_n237), .A3(new_n346), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n332), .A2(G224), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n488), .B2(new_n489), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n487), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n484), .B(new_n480), .C1(new_n252), .C2(new_n435), .ZN(new_n495));
  AOI21_X1  g309(.A(G902), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n484), .B1(new_n252), .B2(new_n435), .ZN(new_n497));
  INV_X1    g311(.A(new_n480), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(KEYINPUT6), .A3(new_n495), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n488), .A2(new_n489), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(new_n490), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n503), .A3(new_n498), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G210), .B1(G237), .B2(G902), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n496), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n496), .B2(new_n505), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n476), .B(new_n479), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n470), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n220), .A2(G128), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n512), .B(KEYINPUT89), .Z(new_n513));
  NAND2_X1  g327(.A1(new_n336), .A2(G128), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n209), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n513), .A2(G134), .A3(new_n514), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n518), .A3(G134), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n190), .A2(G122), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT87), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n190), .A2(G122), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G107), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n419), .A3(new_n523), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT88), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(KEYINPUT88), .A3(new_n526), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n513), .A2(new_n518), .A3(G134), .A4(new_n514), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n520), .A2(new_n529), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n522), .A2(KEYINPUT14), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n523), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n522), .A2(KEYINPUT14), .ZN(new_n535));
  OAI21_X1  g349(.A(G107), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n536), .A2(new_n526), .A3(new_n516), .A4(new_n517), .ZN(new_n537));
  INV_X1    g351(.A(G217), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n468), .A2(new_n538), .A3(G953), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n532), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n532), .B2(new_n537), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(G902), .ZN(new_n543));
  INV_X1    g357(.A(G478), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n543), .A2(new_n545), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n409), .A2(new_n511), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT74), .B(new_n304), .C1(new_n315), .C2(new_n322), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n538), .B1(G234), .B2(new_n298), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G137), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n332), .A2(G221), .A3(G234), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n554), .B(new_n555), .Z(new_n556));
  XOR2_X1   g370(.A(G119), .B(G128), .Z(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT24), .B(G110), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT75), .B1(new_n188), .B2(G128), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n560), .A2(KEYINPUT23), .B1(new_n188), .B2(G128), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(KEYINPUT23), .B2(new_n560), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n559), .B1(new_n562), .B2(G110), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n368), .A2(new_n370), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT78), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n368), .A2(KEYINPUT78), .A3(new_n370), .A4(new_n563), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n557), .A2(new_n558), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n562), .B2(G110), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n367), .A3(new_n340), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n556), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  INV_X1    g387(.A(new_n556), .ZN(new_n574));
  AOI211_X1 g388(.A(new_n573), .B(new_n574), .C1(new_n566), .C2(new_n567), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT25), .B1(new_n576), .B2(new_n298), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  NOR4_X1   g392(.A1(new_n572), .A2(new_n575), .A3(new_n578), .A4(G902), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n553), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n576), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n553), .A2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n325), .A2(new_n551), .A3(new_n552), .A4(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT90), .B(G101), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G3));
  NOR2_X1   g402(.A1(new_n544), .A2(new_n298), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n543), .B2(new_n544), .ZN(new_n590));
  OR3_X1    g404(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT33), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT33), .B1(new_n540), .B2(new_n541), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(G478), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n409), .A2(new_n510), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT91), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n400), .B2(new_n408), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(KEYINPUT91), .A3(new_n510), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n321), .A2(new_n298), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n321), .A2(new_n305), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n470), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(new_n584), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT34), .B(G104), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  NAND3_X1  g425(.A1(new_n605), .A2(new_n510), .A3(new_n607), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n391), .A2(new_n392), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n406), .A2(KEYINPUT20), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n398), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n550), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT92), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT35), .B(G107), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  NAND2_X1  g434(.A1(new_n603), .A2(new_n604), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT93), .ZN(new_n622));
  INV_X1    g436(.A(new_n553), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n568), .A2(new_n571), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n574), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n568), .A2(new_n571), .A3(new_n556), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n298), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n578), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n576), .A2(KEYINPUT25), .A3(new_n298), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n574), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n624), .B(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n583), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n622), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n633), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n580), .A2(new_n635), .A3(KEYINPUT93), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n621), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n551), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  NOR2_X1   g455(.A1(new_n507), .A2(new_n508), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n478), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n475), .A2(G900), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n473), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n550), .A2(new_n643), .A3(new_n615), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT94), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n637), .A2(new_n606), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(new_n325), .A3(new_n552), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  XNOR2_X1  g465(.A(new_n645), .B(KEYINPUT39), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n470), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT40), .Z(new_n654));
  XOR2_X1   g468(.A(new_n642), .B(KEYINPUT38), .Z(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n580), .A2(new_n635), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n656), .A2(new_n657), .A3(new_n549), .A4(new_n478), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n280), .B1(new_n290), .B2(new_n295), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n300), .A2(new_n280), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n298), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n315), .B2(new_n322), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n654), .A2(new_n658), .A3(new_n409), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n238), .ZN(G45));
  NAND3_X1  g479(.A1(new_n325), .A2(new_n649), .A3(new_n552), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT86), .B1(new_n393), .B2(new_n399), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n407), .A2(new_n401), .A3(new_n398), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n595), .B(new_n645), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT95), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT95), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n599), .A2(new_n671), .A3(new_n645), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n643), .A3(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  AND2_X1   g489(.A1(new_n325), .A2(new_n552), .ZN(new_n676));
  INV_X1    g490(.A(new_n600), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT91), .B1(new_n599), .B2(new_n510), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n439), .A2(new_n444), .A3(new_n449), .A4(new_n451), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n449), .B1(new_n439), .B2(new_n455), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n298), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n459), .A3(new_n469), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n676), .A2(new_n679), .A3(new_n585), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND4_X1  g502(.A1(new_n325), .A2(new_n552), .A3(new_n585), .A4(new_n685), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n550), .A2(new_n510), .A3(new_n615), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n190), .ZN(G18));
  NOR2_X1   g506(.A1(new_n684), .A2(new_n509), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n400), .A2(new_n693), .A3(new_n408), .A4(new_n549), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n637), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n325), .A2(new_n695), .A3(new_n552), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  AOI21_X1  g511(.A(new_n549), .B1(new_n400), .B2(new_n408), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n698), .A2(new_n693), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n301), .A2(new_n280), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n314), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n305), .B(KEYINPUT96), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(G902), .B1(new_n311), .B2(new_n314), .ZN(new_n704));
  INV_X1    g518(.A(G472), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT97), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT97), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n602), .A2(new_n707), .A3(G472), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n699), .A2(new_n585), .A3(new_n703), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  INV_X1    g525(.A(KEYINPUT98), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n671), .A2(new_n409), .A3(new_n595), .A4(new_n645), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n671), .B1(new_n599), .B2(new_n645), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n707), .B1(new_n602), .B2(G472), .ZN(new_n716));
  AOI211_X1 g530(.A(KEYINPUT97), .B(new_n705), .C1(new_n321), .C2(new_n298), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n657), .B(new_n703), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n685), .A2(new_n643), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n670), .A2(KEYINPUT98), .A3(new_n672), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n715), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  NAND2_X1  g537(.A1(new_n715), .A2(new_n721), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n604), .A2(KEYINPUT32), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n321), .A2(new_n316), .A3(new_n305), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n584), .B1(new_n727), .B2(new_n304), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n465), .A2(KEYINPUT99), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n463), .A2(new_n730), .A3(new_n464), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n462), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT100), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(G469), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n459), .A2(new_n461), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT100), .B1(new_n732), .B2(new_n458), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n469), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n642), .A2(new_n479), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n724), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n325), .A2(new_n552), .A3(new_n741), .A4(new_n585), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n745), .B1(new_n724), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT101), .B(G131), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G33));
  NAND3_X1  g564(.A1(new_n550), .A2(new_n615), .A3(new_n645), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  NOR2_X1   g567(.A1(new_n667), .A2(new_n668), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n595), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n621), .A3(new_n657), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT44), .ZN(new_n759));
  INV_X1    g573(.A(new_n740), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n462), .B2(new_n465), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n458), .B(new_n761), .C1(new_n733), .C2(KEYINPUT45), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n460), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n459), .B1(new_n763), .B2(KEYINPUT46), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n469), .B(new_n652), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT102), .Z(new_n767));
  AND3_X1   g581(.A1(new_n759), .A2(new_n760), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n207), .ZN(G39));
  OAI21_X1  g583(.A(new_n469), .B1(new_n764), .B2(new_n765), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n325), .A2(new_n552), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n584), .A3(new_n760), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n771), .A2(new_n713), .A3(new_n714), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n363), .ZN(G42));
  NAND3_X1  g589(.A1(new_n656), .A2(new_n479), .A3(new_n469), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n683), .A2(new_n459), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT49), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n755), .A2(new_n776), .A3(new_n584), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n663), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n690), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n676), .A2(new_n585), .A3(new_n685), .A4(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n710), .A2(new_n696), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n686), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n747), .B2(new_n744), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n605), .A2(new_n510), .A3(new_n599), .A4(new_n607), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n586), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT103), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n586), .A2(KEYINPUT103), .A3(new_n789), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n409), .A2(new_n549), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n639), .B1(new_n612), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n718), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n715), .A2(new_n721), .A3(new_n799), .A4(new_n741), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n549), .A2(new_n760), .A3(new_n615), .A4(new_n645), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n325), .A2(new_n649), .A3(new_n552), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n752), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n696), .B(new_n710), .C1(new_n689), .C2(new_n601), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n691), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n670), .A2(KEYINPUT98), .A3(new_n672), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT98), .B1(new_n670), .B2(new_n672), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n746), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT42), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n806), .B1(new_n811), .B2(new_n743), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT112), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n788), .A2(KEYINPUT53), .A3(new_n804), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT105), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n628), .A2(new_n629), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n633), .B1(new_n816), .B2(new_n553), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n815), .B1(new_n817), .B2(new_n645), .ZN(new_n818));
  INV_X1    g632(.A(new_n645), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n630), .A2(KEYINPUT105), .A3(new_n633), .A4(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n643), .B(new_n698), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n738), .A2(new_n469), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n663), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT106), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n739), .B1(new_n727), .B2(new_n662), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT106), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n698), .A2(new_n643), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT105), .B1(new_n657), .B2(new_n819), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n817), .A2(new_n815), .A3(new_n645), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n674), .A2(new_n832), .A3(new_n722), .A4(new_n650), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT108), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n834), .B1(new_n833), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT107), .B1(new_n833), .B2(new_n835), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n722), .A2(new_n650), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT107), .ZN(new_n842));
  INV_X1    g656(.A(new_n666), .ZN(new_n843));
  INV_X1    g657(.A(new_n673), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n843), .A2(new_n844), .B1(new_n824), .B2(new_n831), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT52), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT109), .B1(new_n838), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n839), .A2(new_n846), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n674), .A2(new_n832), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n835), .B1(new_n850), .B2(new_n840), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT108), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT109), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n849), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n814), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT104), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n786), .A2(new_n858), .A3(new_n804), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n796), .B1(new_n790), .B2(new_n791), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n802), .B1(new_n746), .B2(new_n751), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n860), .A2(new_n862), .A3(new_n793), .A4(new_n800), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT104), .B1(new_n812), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n833), .B(new_n835), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n857), .A2(new_n868), .A3(KEYINPUT54), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n757), .A2(new_n472), .A3(new_n471), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n709), .A2(new_n585), .A3(new_n703), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n478), .A3(new_n656), .A4(new_n685), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT114), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n740), .A2(new_n684), .A3(new_n473), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n757), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT115), .Z(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n799), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n771), .B1(new_n469), .B2(new_n777), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n760), .A3(new_n873), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n780), .A2(new_n585), .A3(new_n880), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n754), .A2(new_n594), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n883), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n870), .B1(new_n879), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT51), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n870), .B(new_n891), .C1(new_n879), .C2(new_n888), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n882), .A2(new_n728), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT48), .Z(new_n894));
  INV_X1    g708(.A(new_n599), .ZN(new_n895));
  INV_X1    g709(.A(new_n873), .ZN(new_n896));
  OAI221_X1 g710(.A(new_n471), .B1(new_n895), .B2(new_n886), .C1(new_n896), .C2(new_n719), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n890), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT110), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n838), .A2(new_n847), .A3(KEYINPUT109), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n855), .B1(new_n849), .B2(new_n854), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n859), .A2(new_n864), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n900), .B(new_n867), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n904), .B1(new_n848), .B2(new_n856), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT110), .B1(new_n906), .B2(KEYINPUT53), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n859), .A2(new_n864), .A3(KEYINPUT53), .A4(new_n865), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT111), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n905), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n869), .B(new_n899), .C1(KEYINPUT54), .C2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n781), .B1(new_n912), .B2(new_n913), .ZN(G75));
  INV_X1    g728(.A(new_n814), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n901), .B2(new_n902), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n866), .A2(new_n867), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n298), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(G210), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n500), .A2(new_n504), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n502), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n332), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n919), .B2(KEYINPUT117), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(KEYINPUT117), .B2(new_n919), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n930), .B2(new_n923), .ZN(G51));
  INV_X1    g745(.A(new_n869), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT54), .B1(new_n857), .B2(new_n868), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n460), .B(KEYINPUT57), .Z(new_n935));
  OAI21_X1  g749(.A(new_n457), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n918), .A2(new_n762), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n926), .B1(new_n936), .B2(new_n937), .ZN(G54));
  NAND3_X1  g752(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n404), .A2(new_n405), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n926), .ZN(G60));
  AND2_X1   g757(.A1(new_n591), .A2(new_n592), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n589), .B(KEYINPUT59), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n927), .B1(new_n934), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n932), .ZN(new_n949));
  INV_X1    g763(.A(new_n945), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n947), .B1(new_n951), .B2(new_n944), .ZN(G63));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT118), .Z(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT60), .Z(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n916), .B2(new_n917), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n576), .ZN(new_n959));
  INV_X1    g773(.A(new_n632), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n960), .B(new_n956), .C1(new_n857), .C2(new_n868), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n927), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n953), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT120), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n956), .B1(new_n857), .B2(new_n868), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n965), .A2(KEYINPUT119), .A3(new_n581), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT119), .B1(new_n965), .B2(new_n581), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n961), .A2(KEYINPUT61), .A3(new_n927), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT119), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n958), .B2(new_n576), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n965), .A2(KEYINPUT119), .A3(new_n581), .ZN(new_n973));
  AND4_X1   g787(.A1(new_n964), .A2(new_n969), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n963), .B1(new_n970), .B2(new_n974), .ZN(G66));
  AOI21_X1  g789(.A(new_n332), .B1(new_n474), .B2(G224), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n798), .A2(new_n785), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n978), .B2(new_n332), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n920), .B1(G898), .B2(new_n332), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT121), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT122), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n979), .B(new_n982), .ZN(G69));
  AND2_X1   g797(.A1(new_n286), .A2(new_n287), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n379), .A2(new_n381), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT123), .Z(new_n986));
  XOR2_X1   g800(.A(new_n984), .B(new_n986), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n653), .B(new_n740), .C1(new_n795), .C2(new_n895), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n989), .A2(new_n676), .A3(new_n585), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n768), .A2(new_n774), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n664), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT124), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n988), .B1(new_n998), .B2(G953), .ZN(new_n999));
  NAND2_X1  g813(.A1(G900), .A2(G953), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n767), .A2(new_n728), .A3(new_n827), .ZN(new_n1001));
  INV_X1    g815(.A(new_n752), .ZN(new_n1002));
  NOR4_X1   g816(.A1(new_n768), .A2(new_n1001), .A3(new_n1002), .A4(new_n774), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n748), .A3(new_n992), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n987), .B(new_n1000), .C1(new_n1004), .C2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n999), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n999), .A2(KEYINPUT126), .ZN(new_n1007));
  INV_X1    g821(.A(G900), .ZN(new_n1008));
  OAI21_X1  g822(.A(G953), .B1(new_n447), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1010), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n999), .B(new_n1005), .C1(KEYINPUT126), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(G72));
  XNOR2_X1  g828(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n705), .A2(new_n298), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1015), .B(new_n1016), .Z(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n1004), .B2(new_n978), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n296), .A2(new_n279), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n926), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1017), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n998), .B2(new_n977), .ZN(new_n1022));
  INV_X1    g836(.A(new_n659), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1019), .A2(new_n659), .A3(new_n1021), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n911), .B2(new_n1025), .ZN(G57));
endmodule


