//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(new_n207), .A2(new_n208), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G50), .A2(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI211_X1 g0021(.A(new_n218), .B(new_n221), .C1(G116), .C2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n224), .A2(KEYINPUT66), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(KEYINPUT66), .B1(new_n224), .B2(new_n225), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n205), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n214), .B1(new_n208), .B2(new_n207), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT67), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(G1), .B(G13), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G232), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n255), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G226), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n251), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G41), .A2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n262), .A2(G1), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT69), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n251), .B1(new_n270), .B2(new_n262), .ZN(new_n271));
  INV_X1    g0071(.A(G238), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n265), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n261), .A2(KEYINPUT13), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G97), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n260), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n211), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(KEYINPUT69), .A2(G1), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT69), .A2(G1), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n262), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n264), .B1(new_n286), .B2(G238), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n275), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(G169), .B1(new_n274), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(KEYINPUT14), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT13), .B1(new_n261), .B2(new_n273), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n281), .A2(new_n275), .A3(new_n287), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(new_n292), .A3(G179), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n291), .B2(new_n292), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT14), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n268), .A2(G13), .A3(G20), .A4(new_n269), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G68), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT12), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n249), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G77), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G50), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n302), .B1(new_n212), .B2(G68), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n211), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT11), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(KEYINPUT11), .A3(new_n308), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n308), .B1(new_n284), .B2(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G68), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n290), .A2(new_n297), .B1(new_n300), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n300), .ZN(new_n316));
  AOI21_X1  g0116(.A(G200), .B1(new_n291), .B2(new_n292), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n274), .A2(new_n288), .A3(G190), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n258), .B2(G20), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n220), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G58), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n220), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n330), .B2(new_n201), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n303), .A2(G159), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT16), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT7), .B1(new_n326), .B2(new_n212), .ZN(new_n335));
  NOR4_X1   g0135(.A1(new_n324), .A2(new_n325), .A3(new_n322), .A4(G20), .ZN(new_n336));
  OAI21_X1  g0136(.A(G68), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n332), .A4(new_n331), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n308), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n258), .A2(G223), .A3(new_n259), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n258), .A2(G226), .A3(G1698), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G87), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n280), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n264), .B1(new_n286), .B2(G232), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT74), .B(G190), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n265), .B1(new_n271), .B2(new_n252), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n280), .B2(new_n345), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n351), .B2(G200), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n312), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n353), .B2(new_n298), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n341), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT17), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n307), .A2(new_n211), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n334), .B2(new_n339), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(new_n355), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(KEYINPUT17), .A3(new_n352), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n346), .A2(G179), .A3(new_n347), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n351), .B2(new_n294), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n361), .B2(new_n355), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT18), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT18), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n366), .B(new_n369), .C1(new_n361), .C2(new_n355), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n312), .A2(G77), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G77), .B2(new_n298), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT15), .B(G87), .Z(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n301), .B1(G20), .B2(G77), .ZN(new_n376));
  INV_X1    g0176(.A(new_n353), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n303), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n360), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  OR3_X1    g0180(.A1(new_n326), .A2(KEYINPUT70), .A3(new_n259), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT70), .B1(new_n326), .B2(new_n259), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n219), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n256), .A2(new_n259), .ZN(new_n384));
  INV_X1    g0184(.A(G107), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n258), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n280), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n264), .B1(new_n286), .B2(G244), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(G190), .ZN(new_n390));
  AOI21_X1  g0190(.A(G200), .B1(new_n387), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n380), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n380), .ZN(new_n393));
  INV_X1    g0193(.A(G179), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n294), .B1(new_n387), .B2(new_n388), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n321), .A2(new_n372), .A3(new_n392), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  INV_X1    g0199(.A(G223), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n381), .B2(new_n382), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n258), .A2(new_n259), .ZN(new_n402));
  INV_X1    g0202(.A(G222), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n402), .A2(new_n403), .B1(new_n216), .B2(new_n258), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n280), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n264), .B1(new_n286), .B2(G226), .ZN(new_n406));
  AOI211_X1 g0206(.A(KEYINPUT73), .B(new_n399), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n405), .ZN(new_n408));
  INV_X1    g0208(.A(new_n406), .ZN(new_n409));
  OAI21_X1  g0209(.A(G200), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(G190), .A3(new_n406), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT73), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n407), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT10), .B1(new_n414), .B2(KEYINPUT72), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n298), .A2(new_n305), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n312), .B2(new_n305), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT71), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n417), .B(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n420));
  INV_X1    g0220(.A(G150), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n304), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n353), .A2(G20), .A3(new_n249), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n308), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n425), .A2(KEYINPUT9), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(KEYINPUT9), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n414), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n415), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n408), .A2(new_n409), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G179), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n294), .B2(new_n430), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n414), .B1(KEYINPUT72), .B2(KEYINPUT10), .C1(new_n426), .C2(new_n427), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n398), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G116), .ZN(new_n437));
  OAI21_X1  g0237(.A(G244), .B1(new_n324), .B2(new_n325), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n437), .B1(new_n438), .B2(new_n259), .C1(new_n402), .C2(new_n272), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n280), .ZN(new_n440));
  INV_X1    g0240(.A(G45), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n270), .A2(new_n441), .A3(new_n263), .ZN(new_n442));
  INV_X1    g0242(.A(G250), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n284), .B2(G45), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n251), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G169), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n394), .B2(new_n446), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n268), .A2(G33), .A3(new_n269), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n298), .A2(new_n360), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n375), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n212), .B(G68), .C1(new_n324), .C2(new_n325), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n258), .A2(KEYINPUT79), .A3(new_n212), .A4(G68), .ZN(new_n458));
  NOR3_X1   g0258(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n459));
  AOI21_X1  g0259(.A(G20), .B1(G33), .B2(G97), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT19), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OR3_X1    g0261(.A1(new_n277), .A2(KEYINPUT19), .A3(G20), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n457), .A2(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n360), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  AOI21_X1  g0266(.A(G20), .B1(new_n254), .B2(new_n255), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT79), .B1(new_n467), .B2(G68), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n455), .A2(new_n456), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT80), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n298), .A2(new_n375), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT81), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  AOI211_X1 g0276(.A(new_n476), .B(new_n473), .C1(new_n465), .C2(new_n471), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n454), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n449), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n308), .B1(new_n470), .B2(KEYINPUT80), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n463), .A2(new_n464), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n474), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n476), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n472), .A2(KEYINPUT81), .A3(new_n474), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n453), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT82), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n399), .B1(new_n440), .B2(new_n445), .ZN(new_n488));
  INV_X1    g0288(.A(G87), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n451), .A2(new_n489), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n488), .B(new_n490), .C1(new_n484), .C2(new_n485), .ZN(new_n491));
  INV_X1    g0291(.A(new_n446), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G190), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT83), .ZN(new_n494));
  INV_X1    g0294(.A(G190), .ZN(new_n495));
  OR3_X1    g0295(.A1(new_n446), .A2(KEYINPUT83), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n480), .A2(new_n487), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT76), .B1(new_n499), .B2(G41), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT76), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n250), .A3(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(G274), .B1(new_n279), .B2(new_n211), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(G41), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n268), .A2(new_n506), .A3(G45), .A4(new_n269), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT75), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT75), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n284), .A2(new_n509), .A3(G45), .A4(new_n506), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n505), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(G257), .B(new_n251), .C1(new_n507), .C2(new_n503), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT77), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT77), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n515), .A3(new_n512), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(G1698), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(G244), .C1(new_n325), .C2(new_n324), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n217), .B1(new_n254), .B2(new_n255), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(KEYINPUT4), .ZN(new_n522));
  OAI21_X1  g0322(.A(G250), .B1(new_n324), .B2(new_n325), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n259), .B1(new_n523), .B2(KEYINPUT4), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n280), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n514), .A2(new_n394), .A3(new_n516), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G97), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n298), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(G97), .B2(new_n451), .ZN(new_n529));
  OAI21_X1  g0329(.A(G107), .B1(new_n335), .B2(new_n336), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  AND2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n385), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(G20), .B1(G77), .B2(new_n303), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n529), .B1(new_n538), .B2(new_n308), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n525), .A2(new_n512), .A3(new_n511), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n294), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n526), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT78), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n514), .A2(new_n516), .A3(new_n525), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n525), .A2(G190), .A3(new_n512), .A4(new_n511), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n443), .B1(new_n254), .B2(new_n255), .ZN(new_n550));
  OAI21_X1  g0350(.A(G1698), .B1(new_n550), .B2(new_n517), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n438), .A2(new_n517), .B1(G33), .B2(G283), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n519), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n513), .A2(KEYINPUT77), .B1(new_n280), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n399), .B1(new_n554), .B2(new_n516), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n539), .A2(new_n547), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n555), .A2(KEYINPUT78), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n543), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n550), .A2(new_n259), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n258), .A2(G257), .A3(G1698), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G294), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n280), .ZN(new_n563));
  OAI211_X1 g0363(.A(G264), .B(new_n251), .C1(new_n507), .C2(new_n503), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n511), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n399), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n563), .A2(new_n495), .A3(new_n511), .A4(new_n564), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR3_X1    g0368(.A1(new_n298), .A2(KEYINPUT25), .A3(G107), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n298), .A2(new_n450), .A3(new_n360), .A4(G107), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT25), .B1(new_n298), .B2(G107), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n569), .A2(KEYINPUT86), .A3(new_n570), .A4(new_n571), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(new_n385), .A3(G20), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n576), .B(new_n578), .C1(G20), .C2(new_n437), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n212), .B(G87), .C1(new_n324), .C2(new_n325), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT22), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n258), .A2(new_n582), .A3(new_n212), .A4(G87), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n584), .A2(KEYINPUT24), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n360), .B1(new_n584), .B2(KEYINPUT24), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n574), .A2(new_n575), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT87), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n568), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n568), .B2(new_n587), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT20), .ZN(new_n592));
  INV_X1    g0392(.A(G116), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n212), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n520), .B1(new_n527), .B2(G33), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(new_n212), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n596), .B2(new_n360), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n249), .A2(G97), .ZN(new_n598));
  AOI21_X1  g0398(.A(G20), .B1(new_n598), .B2(new_n520), .ZN(new_n599));
  OAI211_X1 g0399(.A(KEYINPUT20), .B(new_n308), .C1(new_n599), .C2(new_n594), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n298), .A2(new_n450), .A3(new_n360), .A4(G116), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n284), .A2(G13), .A3(G20), .A4(new_n593), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT85), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT85), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT21), .ZN(new_n609));
  OAI211_X1 g0409(.A(G270), .B(new_n251), .C1(new_n507), .C2(new_n503), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n511), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G264), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n612));
  OAI211_X1 g0412(.A(G257), .B(new_n259), .C1(new_n324), .C2(new_n325), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n254), .A2(G303), .A3(new_n255), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n612), .A2(new_n613), .A3(new_n617), .A4(new_n614), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n280), .A3(new_n618), .ZN(new_n619));
  AOI211_X1 g0419(.A(new_n609), .B(new_n294), .C1(new_n611), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n611), .A2(new_n619), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n394), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n608), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT85), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n624), .A2(new_n605), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(G169), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n609), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n611), .A2(new_n348), .A3(new_n619), .ZN(new_n628));
  AOI21_X1  g0428(.A(G200), .B1(new_n611), .B2(new_n619), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n574), .A2(new_n575), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n585), .A2(new_n586), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n565), .A2(G169), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n563), .A2(G179), .A3(new_n511), .A4(new_n564), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n623), .A2(new_n627), .A3(new_n630), .A4(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n558), .A2(new_n591), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n436), .A2(new_n498), .A3(new_n639), .ZN(G372));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n484), .A2(new_n485), .ZN(new_n642));
  INV_X1    g0442(.A(new_n488), .ZN(new_n643));
  INV_X1    g0443(.A(new_n490), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .A4(new_n493), .ZN(new_n645));
  INV_X1    g0445(.A(new_n543), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n478), .A2(new_n448), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n641), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n497), .A2(new_n642), .A3(new_n643), .A4(new_n644), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n448), .B1(new_n486), .B2(KEYINPUT82), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n478), .A2(new_n479), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n649), .B(new_n646), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n648), .B1(KEYINPUT26), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT78), .B1(new_n555), .B2(new_n556), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n546), .A2(new_n548), .A3(new_n544), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n646), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n568), .A2(new_n587), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT87), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n568), .A2(new_n587), .A3(new_n588), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n623), .A2(new_n627), .A3(new_n637), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n656), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n662), .A2(new_n645), .B1(new_n478), .B2(new_n448), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n653), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n436), .ZN(new_n665));
  INV_X1    g0465(.A(new_n371), .ZN(new_n666));
  INV_X1    g0466(.A(new_n315), .ZN(new_n667));
  INV_X1    g0467(.A(new_n397), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT17), .B1(new_n362), .B2(new_n352), .ZN(new_n670));
  AND4_X1   g0470(.A1(KEYINPUT17), .A2(new_n341), .A3(new_n356), .A4(new_n352), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n319), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n666), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n429), .A2(new_n434), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(new_n425), .B2(new_n432), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n665), .A2(new_n676), .ZN(G369));
  AND2_X1   g0477(.A1(new_n623), .A2(new_n627), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n212), .A2(G13), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n284), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n678), .A2(new_n630), .B1(new_n608), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n685), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n625), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n686), .B1(new_n678), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n587), .A2(new_n687), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT88), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n637), .B1(new_n692), .B2(new_n591), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n637), .B2(new_n685), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n637), .A2(new_n685), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n678), .A2(new_n685), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n206), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G1), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n489), .A2(new_n527), .A3(new_n385), .A4(new_n593), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n704), .A2(new_n705), .B1(new_n209), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n563), .A2(new_n564), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n446), .A2(new_n708), .A3(new_n394), .ZN(new_n709));
  INV_X1    g0509(.A(new_n541), .ZN(new_n710));
  INV_X1    g0510(.A(new_n621), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g0512(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n492), .A2(G179), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n545), .A3(new_n565), .A4(new_n621), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n685), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n639), .A2(new_n498), .A3(new_n687), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n685), .A2(KEYINPUT31), .ZN(new_n724));
  INV_X1    g0524(.A(new_n717), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n719), .B1(new_n725), .B2(KEYINPUT90), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G330), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n498), .A2(new_n641), .A3(new_n646), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n645), .A2(new_n647), .A3(new_n646), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT26), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n663), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .A3(new_n687), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n685), .B1(new_n653), .B2(new_n663), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n731), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n707), .B1(new_n739), .B2(G1), .ZN(G364));
  AOI21_X1  g0540(.A(new_n704), .B1(G45), .B2(new_n679), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n690), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n689), .A2(G330), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n689), .A2(G20), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n211), .B1(G20), .B2(new_n294), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n244), .A2(new_n441), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n209), .A2(new_n441), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n701), .B(new_n258), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n701), .A2(new_n326), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G355), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G116), .B2(new_n206), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n750), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n212), .A2(new_n394), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(new_n348), .A3(new_n399), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n212), .B1(new_n761), .B2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n760), .A2(G326), .B1(G294), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT91), .Z(new_n765));
  NOR2_X1   g0565(.A1(new_n399), .A2(G179), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n212), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n767), .A2(new_n761), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n258), .B(new_n770), .C1(G329), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n759), .A2(new_n348), .A3(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G322), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n759), .A2(new_n399), .A3(G190), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(G311), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n766), .A2(G20), .A3(G190), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT92), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G303), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n773), .A2(new_n775), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n763), .A2(G97), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n772), .A2(G159), .ZN(new_n785));
  INV_X1    g0585(.A(new_n778), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n784), .B1(new_n785), .B2(KEYINPUT32), .C1(new_n786), .C2(new_n216), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n768), .A2(new_n385), .ZN(new_n788));
  INV_X1    g0588(.A(new_n780), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n326), .B(new_n788), .C1(G87), .C2(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G58), .A2(new_n774), .B1(new_n776), .B2(G68), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n760), .A2(G50), .B1(new_n785), .B2(KEYINPUT32), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n765), .A2(new_n783), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n742), .B1(new_n794), .B2(new_n749), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n757), .A2(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n743), .A2(new_n744), .B1(new_n747), .B2(new_n796), .ZN(G396));
  OAI211_X1 g0597(.A(new_n392), .B(new_n397), .C1(new_n380), .C2(new_n687), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(new_n397), .B2(new_n687), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n737), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(KEYINPUT97), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n737), .A2(new_n802), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n741), .B1(new_n808), .B2(new_n731), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n731), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n749), .A2(new_n745), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n742), .B1(new_n216), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n258), .B1(new_n781), .B2(G107), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT93), .ZN(new_n814));
  INV_X1    g0614(.A(new_n768), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G87), .B1(new_n772), .B2(G311), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  INV_X1    g0617(.A(new_n774), .ZN(new_n818));
  INV_X1    g0618(.A(new_n760), .ZN(new_n819));
  INV_X1    g0619(.A(G303), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n817), .A2(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n776), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n786), .A2(new_n593), .B1(new_n822), .B2(new_n769), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n814), .A2(new_n784), .A3(new_n816), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n768), .A2(new_n220), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n781), .B2(G50), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT94), .Z(new_n828));
  AOI21_X1  g0628(.A(new_n326), .B1(new_n772), .B2(G132), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n329), .C2(new_n762), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G137), .A2(new_n760), .B1(new_n778), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n832), .B2(new_n818), .C1(new_n421), .C2(new_n822), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT34), .Z(new_n834));
  OAI21_X1  g0634(.A(new_n825), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(KEYINPUT95), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n749), .B1(new_n835), .B2(KEYINPUT95), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n812), .B1(new_n836), .B2(new_n837), .C1(new_n802), .C2(new_n746), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n810), .A2(new_n838), .ZN(G384));
  NAND3_X1  g0639(.A1(new_n738), .A2(new_n436), .A3(new_n736), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n676), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT99), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n397), .A2(new_n685), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n737), .B2(new_n802), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n316), .A2(new_n687), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n315), .A2(new_n319), .A3(KEYINPUT98), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT98), .B1(new_n315), .B2(new_n319), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT98), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n320), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n846), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n315), .A2(new_n319), .A3(KEYINPUT98), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  INV_X1    g0656(.A(new_n683), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n361), .B2(new_n355), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n666), .B2(new_n672), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n357), .A2(new_n367), .A3(new_n858), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n856), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n860), .B(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(new_n858), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n364), .B2(new_n371), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n845), .A2(new_n855), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n868), .B(KEYINPUT39), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n667), .A2(new_n687), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n870), .A2(new_n872), .B1(new_n371), .B2(new_n683), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n842), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n722), .A2(KEYINPUT31), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n720), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT31), .B(new_n685), .C1(new_n717), .C2(new_n719), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT100), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT101), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n868), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT40), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n868), .A2(new_n855), .A3(new_n802), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n868), .B2(new_n883), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n723), .A2(new_n880), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n868), .A2(new_n855), .A3(new_n802), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n890), .A2(new_n435), .A3(new_n398), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n730), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n876), .A2(new_n896), .B1(new_n284), .B2(new_n679), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n876), .B2(new_n896), .ZN(new_n898));
  OR3_X1    g0698(.A1(new_n209), .A2(new_n216), .A3(new_n330), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n305), .A2(G68), .ZN(new_n900));
  AOI211_X1 g0700(.A(G13), .B(new_n284), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(G116), .B(new_n213), .C1(new_n536), .C2(KEYINPUT35), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(KEYINPUT35), .B2(new_n536), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT36), .ZN(new_n904));
  OR3_X1    g0704(.A1(new_n898), .A2(new_n901), .A3(new_n904), .ZN(G367));
  NOR3_X1   g0705(.A1(new_n694), .A2(new_n678), .A3(new_n685), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n540), .A2(new_n685), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n656), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT103), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n646), .A2(new_n685), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n543), .B1(new_n910), .B2(new_n637), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n913), .A2(KEYINPUT42), .B1(new_n687), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n642), .A2(new_n644), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n685), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n919), .A2(new_n647), .A3(new_n645), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT102), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n647), .B2(new_n919), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(KEYINPUT102), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT43), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT43), .B1(new_n922), .B2(new_n923), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n917), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n914), .A2(new_n916), .A3(new_n925), .A4(new_n924), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n695), .A2(new_n912), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n702), .B(KEYINPUT41), .Z(new_n933));
  NAND2_X1  g0733(.A1(new_n912), .A2(new_n699), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT45), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n912), .A2(KEYINPUT44), .A3(new_n699), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT44), .B1(new_n912), .B2(new_n699), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n695), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT45), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n934), .B(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n941), .A2(new_n696), .A3(new_n937), .A4(new_n936), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n694), .B(new_n698), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(new_n690), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n939), .A2(new_n942), .A3(new_n739), .A4(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n933), .B1(new_n945), .B2(new_n739), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n267), .B1(new_n679), .B2(G45), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n932), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n924), .A2(new_n748), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n701), .A2(new_n258), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n239), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n750), .B1(new_n206), .B2(new_n452), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n741), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G283), .A2(new_n778), .B1(new_n776), .B2(G294), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n780), .B2(new_n593), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(new_n820), .C2(new_n818), .ZN(new_n958));
  INV_X1    g0758(.A(new_n781), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n959), .A2(new_n956), .A3(new_n593), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n258), .B1(new_n772), .B2(G317), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n527), .B2(new_n768), .ZN(new_n962));
  XNOR2_X1  g0762(.A(KEYINPUT104), .B(G311), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n760), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n385), .B2(new_n762), .ZN(new_n965));
  NOR4_X1   g0765(.A1(new_n958), .A2(new_n960), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G150), .A2(new_n774), .B1(new_n778), .B2(G50), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n832), .B2(new_n819), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n768), .A2(new_n216), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT105), .B(G137), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n969), .B1(new_n772), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(new_n258), .C1(new_n329), .C2(new_n780), .ZN(new_n973));
  INV_X1    g0773(.A(G159), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n822), .A2(new_n974), .B1(new_n762), .B2(new_n220), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n968), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n966), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT47), .ZN(new_n978));
  INV_X1    g0778(.A(new_n749), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n977), .B2(KEYINPUT47), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n954), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n950), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n949), .A2(new_n982), .ZN(G387));
  AOI22_X1  g0783(.A1(new_n754), .A2(new_n705), .B1(new_n385), .B2(new_n701), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n236), .A2(new_n441), .ZN(new_n985));
  AOI211_X1 g0785(.A(G45), .B(new_n705), .C1(G68), .C2(G77), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n377), .A2(KEYINPUT50), .A3(new_n305), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT50), .B1(new_n377), .B2(new_n305), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n951), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n984), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n742), .B1(new_n991), .B2(new_n750), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G50), .A2(new_n774), .B1(new_n778), .B2(G68), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n452), .B2(new_n762), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n789), .A2(G77), .B1(new_n772), .B2(G150), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n995), .B(new_n258), .C1(new_n527), .C2(new_n768), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n819), .A2(new_n974), .B1(new_n822), .B2(new_n353), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n789), .A2(G294), .B1(new_n763), .B2(G283), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n774), .A2(G317), .B1(new_n776), .B2(new_n963), .ZN(new_n1000));
  INV_X1    g0800(.A(G322), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n820), .B2(new_n786), .C1(new_n1001), .C2(new_n819), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT48), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1006));
  INV_X1    g0806(.A(G326), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n326), .B1(new_n771), .B2(new_n1007), .C1(new_n593), .C2(new_n768), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n1005), .B2(KEYINPUT49), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n998), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n992), .B1(new_n1010), .B2(new_n979), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n694), .B2(new_n748), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n944), .B2(new_n948), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n739), .A2(new_n944), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n702), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n739), .A2(new_n944), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(G393));
  NAND2_X1  g0817(.A1(new_n939), .A2(new_n942), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n1014), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(new_n702), .A3(new_n945), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT107), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT107), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1022), .A3(new_n702), .A4(new_n945), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1018), .A2(new_n947), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n910), .A2(new_n748), .A3(new_n911), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n750), .B1(new_n527), .B2(new_n206), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n247), .B2(new_n951), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G311), .A2(new_n774), .B1(new_n760), .B2(G317), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT52), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n780), .A2(new_n769), .B1(new_n771), .B2(new_n1001), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1030), .A2(new_n258), .A3(new_n788), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n776), .A2(G303), .B1(G116), .B2(new_n763), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n817), .C2(new_n786), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G150), .A2(new_n760), .B1(new_n774), .B2(G159), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT51), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n789), .A2(G68), .B1(new_n772), .B2(G143), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n258), .C1(new_n489), .C2(new_n768), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n762), .A2(new_n216), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n305), .A2(new_n822), .B1(new_n786), .B2(new_n353), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1034), .B1(new_n1042), .B2(KEYINPUT106), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(KEYINPUT106), .B2(new_n1042), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n742), .B(new_n1027), .C1(new_n1044), .C2(new_n749), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1024), .B1(new_n1025), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1021), .A2(new_n1023), .A3(new_n1046), .ZN(G390));
  NOR2_X1   g0847(.A1(new_n800), .A2(new_n801), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n735), .A2(new_n1048), .A3(new_n687), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n843), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1052), .A2(new_n799), .B1(new_n668), .B2(new_n685), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n849), .B2(new_n854), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1051), .B1(new_n731), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(G330), .B1(new_n723), .B2(new_n880), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT109), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT109), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(G330), .C1(new_n723), .C2(new_n880), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1053), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1055), .B1(new_n1060), .B2(new_n855), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT108), .ZN(new_n1062));
  OAI211_X1 g0862(.A(G330), .B(new_n802), .C1(new_n723), .C2(new_n728), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n855), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1054), .B(G330), .C1(new_n723), .C2(new_n880), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1062), .B1(new_n1067), .B2(new_n845), .ZN(new_n1068));
  AOI211_X1 g0868(.A(KEYINPUT108), .B(new_n844), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1061), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n894), .A2(G330), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n676), .A3(new_n840), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n871), .B1(new_n844), .B2(new_n1064), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n870), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1051), .A2(new_n855), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n872), .B1(new_n863), .B2(new_n867), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1075), .A2(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n731), .A2(new_n1054), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1079), .B2(new_n1066), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n703), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1074), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1082), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n948), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n258), .B(new_n826), .C1(G294), .C2(new_n772), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1039), .B1(new_n774), .B2(G116), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n489), .C2(new_n959), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G283), .A2(new_n760), .B1(new_n776), .B2(G107), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n527), .B2(new_n786), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT54), .B(G143), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n760), .A2(G128), .B1(new_n778), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n789), .A2(G150), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1095), .A2(new_n1096), .B1(G159), .B2(new_n763), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n815), .A2(G50), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n326), .B1(new_n772), .B2(G125), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1094), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n776), .A2(new_n971), .ZN(new_n1101));
  INV_X1    g0901(.A(G132), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1101), .B1(new_n1095), .B2(new_n1096), .C1(new_n818), .C2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1089), .A2(new_n1091), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n749), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n742), .B1(new_n353), .B2(new_n811), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n870), .C2(new_n746), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1084), .A2(new_n1086), .A3(new_n1107), .ZN(G378));
  INV_X1    g0908(.A(KEYINPUT117), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n425), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n683), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n435), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1111), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n429), .A2(new_n434), .A3(new_n433), .A4(new_n1113), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n893), .B2(G330), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n730), .B(new_n1119), .C1(new_n887), .C2(new_n892), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1109), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n885), .B1(new_n882), .B2(new_n886), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n890), .A2(new_n889), .A3(new_n891), .ZN(new_n1125));
  OAI21_X1  g0925(.A(G330), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1119), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n893), .A2(G330), .A3(new_n1120), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(KEYINPUT117), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1123), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1060), .A2(new_n855), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1056), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n1054), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT108), .B1(new_n1137), .B2(new_n844), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1067), .A2(new_n1062), .A3(new_n845), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1135), .A2(new_n1055), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1073), .B1(new_n1082), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT57), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n875), .B1(new_n1122), .B2(new_n1121), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1127), .A2(new_n874), .A3(new_n1128), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT57), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n702), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n742), .B1(new_n305), .B2(new_n811), .ZN(new_n1149));
  AOI211_X1 g0949(.A(G41), .B(new_n258), .C1(new_n772), .C2(G283), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n329), .B2(new_n768), .C1(new_n216), .C2(new_n780), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G116), .A2(new_n760), .B1(new_n776), .B2(G97), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n452), .B2(new_n786), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n818), .A2(new_n385), .B1(new_n220), .B2(new_n762), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT112), .Z(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT58), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(KEYINPUT58), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(G33), .A2(G41), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT111), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n305), .C1(G41), .C2(new_n258), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(G124), .B2(new_n772), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n974), .B2(new_n768), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT114), .Z(new_n1164));
  AOI22_X1  g0964(.A1(G128), .A2(new_n774), .B1(new_n776), .B2(G132), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n760), .A2(G125), .B1(G150), .B2(new_n763), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n778), .A2(G137), .B1(new_n789), .B2(new_n1093), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT113), .B(KEYINPUT59), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1164), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AND4_X1   g0972(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .A4(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1149), .B1(new_n979), .B2(new_n1173), .C1(new_n1120), .C2(new_n746), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT115), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1134), .B2(new_n948), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1148), .A2(new_n1176), .ZN(G375));
  INV_X1    g0977(.A(new_n933), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1061), .B(new_n1072), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1074), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1064), .A2(new_n745), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n819), .A2(new_n817), .B1(new_n822), .B2(new_n593), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G107), .B2(new_n778), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n781), .A2(G97), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n258), .B(new_n969), .C1(G303), .C2(new_n772), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n774), .A2(G283), .B1(new_n375), .B2(new_n763), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n819), .A2(new_n1102), .B1(new_n786), .B2(new_n421), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G50), .B2(new_n763), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n781), .A2(G159), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n258), .B1(new_n768), .B2(new_n329), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G128), .B2(new_n772), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n774), .A2(new_n971), .B1(new_n776), .B2(new_n1093), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n979), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n742), .B(new_n1195), .C1(new_n220), .C2(new_n811), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1070), .A2(new_n948), .B1(new_n1181), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1180), .A2(new_n1197), .ZN(G381));
  NOR2_X1   g0998(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1176), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1199), .A2(new_n1200), .A3(G378), .ZN(new_n1201));
  OR3_X1    g1001(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(G387), .A2(new_n1202), .A3(G390), .A4(G381), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(G407));
  INV_X1    g1004(.A(G213), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(G343), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1207), .A2(KEYINPUT118), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(KEYINPUT118), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G213), .B(G407), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT119), .ZN(G409));
  AND3_X1   g1011(.A1(new_n1021), .A2(new_n1023), .A3(new_n1046), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(G387), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(G390), .A2(new_n949), .A3(new_n982), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(G390), .A2(new_n949), .A3(KEYINPUT124), .A4(new_n982), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(G393), .B(G396), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(KEYINPUT125), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1219), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT125), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT60), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1179), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1074), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT122), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT123), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT122), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1228), .A2(new_n1232), .A3(new_n1074), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n702), .B1(new_n1179), .B2(new_n1227), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1197), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1234), .B1(new_n1229), .B2(KEYINPUT122), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1231), .B1(new_n1238), .B2(new_n1233), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1226), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1230), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT123), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1242), .A2(G384), .A3(new_n1197), .A4(new_n1236), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1206), .ZN(new_n1245));
  INV_X1    g1045(.A(G2897), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1084), .A2(new_n1086), .A3(new_n1107), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT121), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1144), .A2(new_n1145), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n948), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1130), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1121), .A2(new_n1122), .A3(new_n1109), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT117), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1141), .A2(new_n1257), .A3(new_n1178), .A4(new_n1131), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1174), .B(new_n1253), .C1(new_n1258), .C2(KEYINPUT120), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1258), .A2(KEYINPUT120), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1249), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1176), .C1(new_n1142), .C2(new_n1147), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1245), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1240), .B(new_n1243), .C1(new_n1246), .C2(new_n1245), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1248), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(KEYINPUT126), .A3(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1263), .A2(new_n1245), .A3(new_n1240), .A4(new_n1243), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1244), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1272), .A2(KEYINPUT62), .A3(new_n1245), .A4(new_n1263), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT126), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1225), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1225), .A2(KEYINPUT61), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1269), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT63), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1266), .A2(KEYINPUT63), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1278), .B(new_n1280), .C1(new_n1281), .C2(new_n1279), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1282), .ZN(G405));
  NAND3_X1  g1083(.A1(new_n1148), .A2(new_n1249), .A3(new_n1176), .ZN(new_n1284));
  OAI21_X1  g1084(.A(G378), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1244), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1244), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(new_n1225), .A2(KEYINPUT127), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1288), .A2(new_n1292), .A3(new_n1293), .ZN(G402));
endmodule


