

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  XNOR2_X1 U325 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n418) );
  XNOR2_X1 U326 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U327 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U328 ( .A(n376), .B(n375), .ZN(n379) );
  XNOR2_X1 U329 ( .A(n409), .B(n382), .ZN(n383) );
  XNOR2_X1 U330 ( .A(n408), .B(n383), .ZN(n588) );
  XNOR2_X1 U331 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U332 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(G85GAT), .B(G162GAT), .Z(n295) );
  XNOR2_X1 U334 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n293), .B(KEYINPUT2), .ZN(n422) );
  XNOR2_X1 U336 ( .A(G29GAT), .B(n422), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n318) );
  XOR2_X1 U338 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n297) );
  XNOR2_X1 U339 ( .A(KEYINPUT5), .B(KEYINPUT97), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U341 ( .A(KEYINPUT96), .B(n298), .Z(n300) );
  NAND2_X1 U342 ( .A1(G225GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U344 ( .A(n301), .B(KEYINPUT94), .Z(n307) );
  XNOR2_X1 U345 ( .A(G120GAT), .B(KEYINPUT81), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n302), .B(KEYINPUT0), .ZN(n303) );
  XOR2_X1 U347 ( .A(n303), .B(KEYINPUT82), .Z(n305) );
  XNOR2_X1 U348 ( .A(G113GAT), .B(G134GAT), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n305), .B(n304), .ZN(n452) );
  XNOR2_X1 U350 ( .A(n452), .B(KEYINPUT92), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n315) );
  XOR2_X1 U352 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n309) );
  XNOR2_X1 U353 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U355 ( .A(KEYINPUT91), .B(G57GAT), .Z(n311) );
  XNOR2_X1 U356 ( .A(G127GAT), .B(G148GAT), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U358 ( .A(n313), .B(n312), .Z(n314) );
  XNOR2_X1 U359 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U360 ( .A(G155GAT), .B(n316), .Z(n317) );
  XNOR2_X1 U361 ( .A(n318), .B(n317), .ZN(n499) );
  XOR2_X1 U362 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n320) );
  XNOR2_X1 U363 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n319) );
  XNOR2_X1 U364 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(n321), .ZN(n457) );
  XOR2_X1 U366 ( .A(G197GAT), .B(KEYINPUT21), .Z(n423) );
  XOR2_X1 U367 ( .A(KEYINPUT98), .B(n423), .Z(n323) );
  NAND2_X1 U368 ( .A1(G226GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n323), .B(n322), .ZN(n325) );
  XNOR2_X1 U370 ( .A(G8GAT), .B(G183GAT), .ZN(n324) );
  XNOR2_X1 U371 ( .A(n324), .B(G211GAT), .ZN(n350) );
  XOR2_X1 U372 ( .A(n325), .B(n350), .Z(n331) );
  XOR2_X1 U373 ( .A(G92GAT), .B(G64GAT), .Z(n327) );
  XNOR2_X1 U374 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U376 ( .A(G176GAT), .B(n328), .Z(n345) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(G190GAT), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n329), .B(G218GAT), .ZN(n363) );
  XNOR2_X1 U379 ( .A(n345), .B(n363), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n457), .B(n332), .ZN(n529) );
  INV_X1 U382 ( .A(n529), .ZN(n502) );
  XOR2_X1 U383 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n334) );
  XNOR2_X1 U384 ( .A(G71GAT), .B(G57GAT), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n353) );
  XOR2_X1 U386 ( .A(KEYINPUT33), .B(n353), .Z(n336) );
  XOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .Z(n377) );
  XNOR2_X1 U388 ( .A(G120GAT), .B(n377), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n341) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(G78GAT), .ZN(n337) );
  XOR2_X1 U391 ( .A(n337), .B(G148GAT), .Z(n421) );
  XNOR2_X1 U392 ( .A(n421), .B(KEYINPUT76), .ZN(n339) );
  NAND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U395 ( .A(n341), .B(n340), .Z(n347) );
  XOR2_X1 U396 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n343) );
  XNOR2_X1 U397 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n582) );
  XOR2_X1 U401 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n349) );
  XNOR2_X1 U402 ( .A(KEYINPUT79), .B(KEYINPUT14), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n362) );
  XOR2_X1 U404 ( .A(n350), .B(KEYINPUT15), .Z(n352) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U408 ( .A(G15GAT), .B(G127GAT), .Z(n443) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G155GAT), .Z(n424) );
  XOR2_X1 U410 ( .A(n443), .B(n424), .Z(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n358) );
  INV_X1 U412 ( .A(G64GAT), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U414 ( .A(G1GAT), .B(KEYINPUT70), .Z(n397) );
  XNOR2_X1 U415 ( .A(n397), .B(G78GAT), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n411) );
  INV_X1 U418 ( .A(n411), .ZN(n493) );
  XOR2_X1 U419 ( .A(G50GAT), .B(G162GAT), .Z(n427) );
  XNOR2_X1 U420 ( .A(n363), .B(n427), .ZN(n367) );
  INV_X1 U421 ( .A(n367), .ZN(n365) );
  AND2_X1 U422 ( .A1(G232GAT), .A2(G233GAT), .ZN(n366) );
  INV_X1 U423 ( .A(n366), .ZN(n364) );
  NAND2_X1 U424 ( .A1(n365), .A2(n364), .ZN(n369) );
  NAND2_X1 U425 ( .A1(n367), .A2(n366), .ZN(n368) );
  NAND2_X1 U426 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n370), .B(G92GAT), .ZN(n376) );
  XOR2_X1 U428 ( .A(G29GAT), .B(G43GAT), .Z(n372) );
  XNOR2_X1 U429 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n398) );
  XOR2_X1 U431 ( .A(n398), .B(G134GAT), .Z(n374) );
  INV_X1 U432 ( .A(KEYINPUT10), .ZN(n373) );
  XNOR2_X1 U433 ( .A(G106GAT), .B(n377), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n408) );
  XOR2_X1 U435 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT11), .B(KEYINPUT77), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n409) );
  XNOR2_X1 U438 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n382) );
  NOR2_X1 U439 ( .A1(n493), .A2(n588), .ZN(n384) );
  XOR2_X1 U440 ( .A(KEYINPUT45), .B(n384), .Z(n385) );
  NOR2_X1 U441 ( .A1(n582), .A2(n385), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n386), .B(KEYINPUT116), .ZN(n407) );
  XOR2_X1 U443 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n388) );
  XNOR2_X1 U444 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n406) );
  XOR2_X1 U446 ( .A(G141GAT), .B(G197GAT), .Z(n390) );
  XNOR2_X1 U447 ( .A(G50GAT), .B(G36GAT), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U449 ( .A(G113GAT), .B(G15GAT), .Z(n392) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(G22GAT), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U452 ( .A(n394), .B(n393), .Z(n404) );
  XOR2_X1 U453 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n396) );
  XNOR2_X1 U454 ( .A(KEYINPUT67), .B(KEYINPUT71), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n402) );
  XOR2_X1 U456 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U457 ( .A1(G229GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n565) );
  INV_X1 U462 ( .A(n565), .ZN(n577) );
  NAND2_X1 U463 ( .A1(n407), .A2(n577), .ZN(n416) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n563) );
  XOR2_X1 U465 ( .A(n582), .B(KEYINPUT41), .Z(n567) );
  NAND2_X1 U466 ( .A1(n567), .A2(n565), .ZN(n410) );
  XNOR2_X1 U467 ( .A(KEYINPUT46), .B(n410), .ZN(n412) );
  XNOR2_X1 U468 ( .A(KEYINPUT115), .B(n411), .ZN(n573) );
  NAND2_X1 U469 ( .A1(n412), .A2(n573), .ZN(n413) );
  NOR2_X1 U470 ( .A1(n563), .A2(n413), .ZN(n414) );
  XNOR2_X1 U471 ( .A(KEYINPUT47), .B(n414), .ZN(n415) );
  NAND2_X1 U472 ( .A1(n416), .A2(n415), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n417), .B(KEYINPUT48), .ZN(n536) );
  NAND2_X1 U474 ( .A1(n502), .A2(n536), .ZN(n419) );
  NOR2_X1 U475 ( .A1(n499), .A2(n420), .ZN(n576) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n438) );
  XOR2_X1 U477 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U480 ( .A(n428), .B(n427), .Z(n436) );
  XOR2_X1 U481 ( .A(KEYINPUT24), .B(G204GAT), .Z(n430) );
  XNOR2_X1 U482 ( .A(G218GAT), .B(KEYINPUT90), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U484 ( .A(KEYINPUT22), .B(G211GAT), .Z(n432) );
  XNOR2_X1 U485 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n476) );
  NAND2_X1 U490 ( .A1(n576), .A2(n476), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n439), .B(KEYINPUT55), .ZN(n459) );
  XOR2_X1 U492 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n441) );
  XNOR2_X1 U493 ( .A(G190GAT), .B(G71GAT), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U495 ( .A(n442), .B(G99GAT), .Z(n445) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n456) );
  XOR2_X1 U498 ( .A(KEYINPUT65), .B(KEYINPUT83), .Z(n447) );
  XNOR2_X1 U499 ( .A(G183GAT), .B(G176GAT), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT88), .B(n448), .Z(n450) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U504 ( .A(n451), .B(KEYINPUT87), .Z(n454) );
  XNOR2_X1 U505 ( .A(n452), .B(KEYINPUT86), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n458) );
  XNOR2_X1 U508 ( .A(n458), .B(n457), .ZN(n518) );
  NAND2_X1 U509 ( .A1(n459), .A2(n518), .ZN(n460) );
  XNOR2_X1 U510 ( .A(n460), .B(KEYINPUT123), .ZN(n571) );
  NAND2_X1 U511 ( .A1(n571), .A2(n563), .ZN(n464) );
  XNOR2_X1 U512 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n462) );
  XOR2_X1 U513 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n461) );
  XNOR2_X1 U514 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n483) );
  NOR2_X1 U515 ( .A1(n577), .A2(n582), .ZN(n497) );
  NOR2_X1 U516 ( .A1(n493), .A2(n563), .ZN(n466) );
  XNOR2_X1 U517 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n466), .B(n465), .ZN(n480) );
  INV_X1 U519 ( .A(n499), .ZN(n526) );
  NAND2_X1 U520 ( .A1(n518), .A2(n502), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n476), .A2(n467), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n468), .Z(n472) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(n502), .ZN(n474) );
  NOR2_X1 U524 ( .A1(n518), .A2(n476), .ZN(n470) );
  XNOR2_X1 U525 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n470), .B(n469), .ZN(n575) );
  NAND2_X1 U527 ( .A1(n474), .A2(n575), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n526), .A2(n473), .ZN(n479) );
  NAND2_X1 U530 ( .A1(n474), .A2(n499), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n475), .B(KEYINPUT99), .ZN(n537) );
  XOR2_X1 U532 ( .A(KEYINPUT28), .B(n476), .Z(n541) );
  NOR2_X1 U533 ( .A1(n518), .A2(n541), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n537), .A2(n477), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n492) );
  AND2_X1 U536 ( .A1(n480), .A2(n492), .ZN(n513) );
  NAND2_X1 U537 ( .A1(n497), .A2(n513), .ZN(n481) );
  XNOR2_X1 U538 ( .A(KEYINPUT101), .B(n481), .ZN(n488) );
  NAND2_X1 U539 ( .A1(n499), .A2(n488), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n502), .A2(n488), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n486) );
  NAND2_X1 U544 ( .A1(n488), .A2(n518), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n541), .A2(n488), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n491) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n501) );
  NAND2_X1 U552 ( .A1(n493), .A2(n492), .ZN(n494) );
  NOR2_X1 U553 ( .A1(n588), .A2(n494), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT37), .B(n495), .Z(n496) );
  XNOR2_X1 U555 ( .A(KEYINPUT104), .B(n496), .ZN(n524) );
  NAND2_X1 U556 ( .A1(n524), .A2(n497), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT38), .B(n498), .Z(n507) );
  NAND2_X1 U558 ( .A1(n507), .A2(n499), .ZN(n500) );
  XOR2_X1 U559 ( .A(n501), .B(n500), .Z(G1328GAT) );
  NAND2_X1 U560 ( .A1(n507), .A2(n502), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n505) );
  NAND2_X1 U563 ( .A1(n507), .A2(n518), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n509) );
  NAND2_X1 U567 ( .A1(n507), .A2(n541), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n512) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  XNOR2_X1 U572 ( .A(n512), .B(n511), .ZN(n515) );
  AND2_X1 U573 ( .A1(n577), .A2(n567), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n513), .A2(n525), .ZN(n520) );
  NOR2_X1 U575 ( .A1(n526), .A2(n520), .ZN(n514) );
  XOR2_X1 U576 ( .A(n515), .B(n514), .Z(n516) );
  XNOR2_X1 U577 ( .A(KEYINPUT110), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n529), .A2(n520), .ZN(n517) );
  XOR2_X1 U579 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  INV_X1 U580 ( .A(n518), .ZN(n538) );
  NOR2_X1 U581 ( .A1(n538), .A2(n520), .ZN(n519) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n519), .Z(G1334GAT) );
  INV_X1 U583 ( .A(n541), .ZN(n533) );
  NOR2_X1 U584 ( .A1(n533), .A2(n520), .ZN(n522) );
  XNOR2_X1 U585 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U587 ( .A(G78GAT), .B(n523), .Z(G1335GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n532) );
  NOR2_X1 U589 ( .A1(n526), .A2(n532), .ZN(n527) );
  XOR2_X1 U590 ( .A(G85GAT), .B(n527), .Z(n528) );
  XNOR2_X1 U591 ( .A(KEYINPUT114), .B(n528), .ZN(G1336GAT) );
  NOR2_X1 U592 ( .A1(n529), .A2(n532), .ZN(n530) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n530), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n538), .A2(n532), .ZN(n531) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n531), .Z(G1338GAT) );
  NOR2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U597 ( .A(G106GAT), .B(n534), .Z(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT44), .B(n535), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n537), .ZN(n555) );
  NOR2_X1 U600 ( .A1(n538), .A2(n555), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n539), .B(KEYINPUT117), .ZN(n540) );
  NOR2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT118), .B(n542), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n551), .A2(n565), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U607 ( .A1(n567), .A2(n551), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n547) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(KEYINPUT120), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n550) );
  INV_X1 U612 ( .A(n551), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n573), .A2(n548), .ZN(n549) );
  XOR2_X1 U614 ( .A(n550), .B(n549), .Z(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U616 ( .A1(n551), .A2(n563), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  XOR2_X1 U618 ( .A(G141GAT), .B(KEYINPUT121), .Z(n557) );
  INV_X1 U619 ( .A(n575), .ZN(n554) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n562), .A2(n565), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U624 ( .A1(n562), .A2(n567), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n411), .A2(n562), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n571), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n571), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G176GAT), .ZN(G1349GAT) );
  INV_X1 U637 ( .A(n571), .ZN(n572) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n581) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n587) );
  NOR2_X1 U642 ( .A1(n577), .A2(n587), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U647 ( .A(n587), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n411), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

