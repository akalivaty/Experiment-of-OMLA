

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779;

  INV_X1 U370 ( .A(n658), .ZN(n349) );
  NOR2_X1 U371 ( .A1(n421), .A2(G953), .ZN(n420) );
  AND2_X2 U372 ( .A1(n432), .A2(n430), .ZN(n429) );
  XNOR2_X2 U373 ( .A(n641), .B(KEYINPUT62), .ZN(n642) );
  XNOR2_X2 U374 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X2 U375 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n583) );
  AND2_X2 U376 ( .A1(n644), .A2(G953), .ZN(n749) );
  XNOR2_X1 U377 ( .A(n348), .B(KEYINPUT87), .ZN(n596) );
  NAND2_X1 U378 ( .A1(n408), .A2(n410), .ZN(n348) );
  NAND2_X1 U379 ( .A1(n350), .A2(n349), .ZN(n572) );
  INV_X1 U380 ( .A(n674), .ZN(n350) );
  AND2_X2 U381 ( .A1(n565), .A2(n580), .ZN(n365) );
  NOR2_X4 U382 ( .A1(n569), .A2(n560), .ZN(n355) );
  XNOR2_X2 U383 ( .A(n405), .B(KEYINPUT0), .ZN(n569) );
  NAND2_X1 U384 ( .A1(n617), .A2(n354), .ZN(n628) );
  XNOR2_X1 U385 ( .A(n611), .B(n612), .ZN(n354) );
  INV_X2 U386 ( .A(G131), .ZN(n456) );
  BUF_X2 U387 ( .A(n603), .Z(n698) );
  XNOR2_X1 U388 ( .A(G107), .B(G110), .ZN(n522) );
  XNOR2_X2 U389 ( .A(n533), .B(n532), .ZN(n534) );
  INV_X1 U390 ( .A(n668), .ZN(n671) );
  NAND2_X1 U391 ( .A1(n571), .A2(n570), .ZN(n668) );
  XNOR2_X1 U392 ( .A(n607), .B(KEYINPUT40), .ZN(n779) );
  XNOR2_X1 U393 ( .A(n626), .B(n625), .ZN(n776) );
  XNOR2_X1 U394 ( .A(n390), .B(KEYINPUT19), .ZN(n609) );
  NAND2_X1 U395 ( .A1(n554), .A2(n682), .ZN(n390) );
  XNOR2_X1 U396 ( .A(n552), .B(n551), .ZN(n554) );
  INV_X2 U397 ( .A(G110), .ZN(n356) );
  NAND2_X1 U398 ( .A1(n428), .A2(n738), .ZN(n427) );
  AND2_X1 U399 ( .A1(n364), .A2(n637), .ZN(n723) );
  NOR2_X1 U400 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U401 ( .A(n406), .B(KEYINPUT32), .ZN(n778) );
  AND2_X1 U402 ( .A1(n630), .A2(n671), .ZN(n607) );
  AND2_X1 U403 ( .A1(n604), .A2(n447), .ZN(n619) );
  XNOR2_X1 U404 ( .A(n490), .B(n640), .ZN(n603) );
  XNOR2_X1 U405 ( .A(n550), .B(KEYINPUT93), .ZN(n551) );
  XNOR2_X1 U406 ( .A(n420), .B(n422), .ZN(n493) );
  NAND2_X1 U407 ( .A1(n549), .A2(G214), .ZN(n682) );
  XNOR2_X1 U408 ( .A(n455), .B(G137), .ZN(n454) );
  NAND2_X1 U409 ( .A1(G237), .A2(G234), .ZN(n510) );
  INV_X2 U410 ( .A(KEYINPUT4), .ZN(n455) );
  XOR2_X2 U411 ( .A(G140), .B(G104), .Z(n523) );
  XNOR2_X1 U412 ( .A(G116), .B(G119), .ZN(n486) );
  XNOR2_X2 U413 ( .A(n355), .B(KEYINPUT22), .ZN(n589) );
  XNOR2_X2 U414 ( .A(n356), .B(G119), .ZN(n542) );
  BUF_X1 U415 ( .A(n372), .Z(n357) );
  BUF_X1 U416 ( .A(n554), .Z(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n743), .ZN(n452) );
  NOR2_X1 U418 ( .A1(n742), .A2(n387), .ZN(n359) );
  BUF_X1 U419 ( .A(n745), .Z(n360) );
  BUF_X1 U420 ( .A(n409), .Z(n361) );
  XNOR2_X1 U421 ( .A(n441), .B(n561), .ZN(n409) );
  INV_X1 U422 ( .A(n569), .ZN(n565) );
  INV_X4 U423 ( .A(G953), .ZN(n769) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n482) );
  NOR2_X1 U425 ( .A1(n426), .A2(n505), .ZN(n425) );
  XNOR2_X1 U426 ( .A(n480), .B(n479), .ZN(n582) );
  NOR2_X1 U427 ( .A1(G902), .A2(n650), .ZN(n479) );
  XNOR2_X1 U428 ( .A(n608), .B(KEYINPUT46), .ZN(n444) );
  AND2_X1 U429 ( .A1(n574), .A2(n573), .ZN(n408) );
  XNOR2_X1 U430 ( .A(G902), .B(KEYINPUT92), .ZN(n504) );
  XNOR2_X1 U431 ( .A(n466), .B(G125), .ZN(n535) );
  INV_X1 U432 ( .A(G234), .ZN(n421) );
  XOR2_X1 U433 ( .A(KEYINPUT7), .B(G122), .Z(n461) );
  XNOR2_X1 U434 ( .A(KEYINPUT9), .B(KEYINPUT104), .ZN(n457) );
  XOR2_X1 U435 ( .A(KEYINPUT105), .B(KEYINPUT103), .Z(n458) );
  INV_X1 U436 ( .A(G134), .ZN(n460) );
  XNOR2_X1 U437 ( .A(KEYINPUT99), .B(KEYINPUT97), .ZN(n473) );
  XOR2_X1 U438 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n474) );
  XOR2_X1 U439 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n472) );
  XNOR2_X1 U440 ( .A(n376), .B(n543), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n481), .B(n377), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n775), .B(n378), .ZN(n377) );
  INV_X1 U443 ( .A(KEYINPUT11), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n448), .B(KEYINPUT30), .ZN(n447) );
  INV_X1 U445 ( .A(n682), .ZN(n449) );
  INV_X1 U446 ( .A(KEYINPUT1), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n413), .B(n412), .ZN(n508) );
  XNOR2_X1 U448 ( .A(n507), .B(KEYINPUT96), .ZN(n412) );
  XNOR2_X1 U449 ( .A(n435), .B(n540), .ZN(n434) );
  XNOR2_X1 U450 ( .A(n485), .B(n436), .ZN(n435) );
  XNOR2_X1 U451 ( .A(n486), .B(n437), .ZN(n436) );
  XOR2_X1 U452 ( .A(G116), .B(G107), .Z(n544) );
  XNOR2_X1 U453 ( .A(n468), .B(n467), .ZN(n762) );
  XOR2_X1 U454 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n468) );
  XNOR2_X1 U455 ( .A(n535), .B(G140), .ZN(n467) );
  XNOR2_X1 U456 ( .A(n542), .B(G128), .ZN(n492) );
  INV_X1 U457 ( .A(n723), .ZN(n414) );
  XNOR2_X1 U458 ( .A(n528), .B(n403), .ZN(n740) );
  NAND2_X1 U459 ( .A1(n599), .A2(n394), .ZN(n393) );
  INV_X1 U460 ( .A(n689), .ZN(n394) );
  NOR2_X1 U461 ( .A1(n668), .A2(n622), .ZN(n379) );
  AND2_X1 U462 ( .A1(n373), .A2(n450), .ZN(n610) );
  XNOR2_X1 U463 ( .A(n374), .B(KEYINPUT28), .ZN(n373) );
  NOR2_X1 U464 ( .A1(n698), .A2(n598), .ZN(n374) );
  XNOR2_X1 U465 ( .A(n603), .B(n491), .ZN(n576) );
  BUF_X1 U466 ( .A(n740), .Z(n389) );
  INV_X1 U467 ( .A(G237), .ZN(n519) );
  XNOR2_X1 U468 ( .A(n506), .B(KEYINPUT20), .ZN(n516) );
  INV_X1 U469 ( .A(G902), .ZN(n520) );
  NAND2_X1 U470 ( .A1(n516), .A2(G217), .ZN(n413) );
  INV_X1 U471 ( .A(KEYINPUT78), .ZN(n437) );
  INV_X1 U472 ( .A(KEYINPUT48), .ZN(n442) );
  XNOR2_X1 U473 ( .A(n481), .B(n454), .ZN(n453) );
  XNOR2_X1 U474 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n494) );
  INV_X1 U475 ( .A(KEYINPUT65), .ZN(n416) );
  INV_X1 U476 ( .A(KEYINPUT66), .ZN(n489) );
  XNOR2_X1 U477 ( .A(KEYINPUT18), .B(KEYINPUT91), .ZN(n536) );
  XOR2_X1 U478 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n511) );
  INV_X1 U479 ( .A(KEYINPUT3), .ZN(n487) );
  XNOR2_X1 U480 ( .A(n396), .B(n395), .ZN(n743) );
  XNOR2_X1 U481 ( .A(n462), .B(n366), .ZN(n395) );
  XNOR2_X1 U482 ( .A(n478), .B(n391), .ZN(n650) );
  INV_X1 U483 ( .A(n762), .ZN(n391) );
  XNOR2_X1 U484 ( .A(n477), .B(n375), .ZN(n478) );
  BUF_X1 U485 ( .A(n681), .Z(n715) );
  NAND2_X1 U486 ( .A1(n400), .A2(KEYINPUT34), .ZN(n399) );
  AND2_X1 U487 ( .A1(n699), .A2(n450), .ZN(n604) );
  XNOR2_X1 U488 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U489 ( .A(G478), .ZN(n387) );
  NOR2_X1 U490 ( .A1(n431), .A2(n749), .ZN(n430) );
  NOR2_X1 U491 ( .A1(n440), .A2(G210), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n392), .B(n601), .ZN(n774) );
  XNOR2_X1 U493 ( .A(n381), .B(n380), .ZN(n615) );
  INV_X1 U494 ( .A(KEYINPUT36), .ZN(n380) );
  AND2_X1 U495 ( .A1(n584), .A2(n576), .ZN(n407) );
  INV_X1 U496 ( .A(G143), .ZN(n469) );
  INV_X1 U497 ( .A(KEYINPUT109), .ZN(n625) );
  INV_X1 U498 ( .A(KEYINPUT86), .ZN(n561) );
  XNOR2_X1 U499 ( .A(n424), .B(n423), .ZN(n741) );
  XNOR2_X1 U500 ( .A(n389), .B(n739), .ZN(n423) );
  XOR2_X1 U501 ( .A(n621), .B(KEYINPUT81), .Z(n362) );
  AND2_X1 U502 ( .A1(n521), .A2(n682), .ZN(n363) );
  AND2_X1 U503 ( .A1(n638), .A2(KEYINPUT2), .ZN(n364) );
  XOR2_X1 U504 ( .A(n461), .B(n544), .Z(n366) );
  AND2_X1 U505 ( .A1(n576), .A2(n563), .ZN(n367) );
  XNOR2_X1 U506 ( .A(KEYINPUT90), .B(KEYINPUT33), .ZN(n368) );
  INV_X1 U507 ( .A(KEYINPUT34), .ZN(n580) );
  OR2_X1 U508 ( .A1(n505), .A2(n719), .ZN(n369) );
  AND2_X1 U509 ( .A1(n440), .A2(G210), .ZN(n370) );
  INV_X1 U510 ( .A(n749), .ZN(n439) );
  AND2_X1 U511 ( .A1(n371), .A2(n425), .ZN(n634) );
  XNOR2_X2 U512 ( .A(n443), .B(n442), .ZN(n371) );
  NAND2_X1 U513 ( .A1(n371), .A2(n633), .ZN(n765) );
  XNOR2_X2 U514 ( .A(n453), .B(n372), .ZN(n763) );
  XNOR2_X1 U515 ( .A(n463), .B(n357), .ZN(n396) );
  XNOR2_X2 U516 ( .A(n537), .B(n460), .ZN(n372) );
  AND2_X1 U517 ( .A1(n609), .A2(n610), .ZN(n665) );
  XNOR2_X2 U518 ( .A(n470), .B(G113), .ZN(n543) );
  XNOR2_X2 U519 ( .A(n456), .B(KEYINPUT70), .ZN(n481) );
  NAND2_X1 U520 ( .A1(n363), .A2(n671), .ZN(n614) );
  NAND2_X1 U521 ( .A1(n363), .A2(n379), .ZN(n381) );
  NAND2_X1 U522 ( .A1(n744), .A2(G469), .ZN(n424) );
  BUF_X1 U523 ( .A(n737), .Z(n382) );
  NOR2_X1 U524 ( .A1(n603), .A2(n449), .ZN(n448) );
  XNOR2_X1 U525 ( .A(n411), .B(n583), .ZN(n383) );
  XNOR2_X1 U526 ( .A(n411), .B(n583), .ZN(n777) );
  NAND2_X1 U527 ( .A1(n695), .A2(n694), .ZN(n564) );
  XNOR2_X1 U528 ( .A(n501), .B(n500), .ZN(n502) );
  NAND2_X1 U529 ( .A1(n361), .A2(n562), .ZN(n384) );
  NAND2_X1 U530 ( .A1(n409), .A2(n562), .ZN(n574) );
  INV_X1 U531 ( .A(n565), .ZN(n385) );
  INV_X1 U532 ( .A(n585), .ZN(n563) );
  NAND2_X1 U533 ( .A1(n699), .A2(n585), .ZN(n575) );
  XNOR2_X2 U534 ( .A(n567), .B(n388), .ZN(n585) );
  XNOR2_X2 U535 ( .A(G122), .B(G104), .ZN(n470) );
  NAND2_X1 U536 ( .A1(n493), .A2(G221), .ZN(n499) );
  XNOR2_X2 U537 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n532) );
  NAND2_X1 U538 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U539 ( .A(n502), .B(n762), .ZN(n745) );
  XNOR2_X1 U540 ( .A(n534), .B(n535), .ZN(n539) );
  AND2_X2 U541 ( .A1(n398), .A2(n397), .ZN(n401) );
  NOR2_X2 U542 ( .A1(n645), .A2(n749), .ZN(n647) );
  NOR2_X2 U543 ( .A1(n653), .A2(n749), .ZN(n655) );
  NAND2_X1 U544 ( .A1(n716), .A2(n610), .ZN(n392) );
  XNOR2_X2 U545 ( .A(n393), .B(KEYINPUT41), .ZN(n716) );
  NOR2_X1 U546 ( .A1(n565), .A2(n580), .ZN(n402) );
  NAND2_X1 U547 ( .A1(n365), .A2(n681), .ZN(n397) );
  NOR2_X1 U548 ( .A1(n402), .A2(n362), .ZN(n398) );
  NAND2_X2 U549 ( .A1(n401), .A2(n399), .ZN(n411) );
  INV_X1 U550 ( .A(n681), .ZN(n400) );
  XNOR2_X2 U551 ( .A(n579), .B(n368), .ZN(n681) );
  NOR2_X2 U552 ( .A1(n740), .A2(G902), .ZN(n404) );
  XNOR2_X1 U553 ( .A(n527), .B(n526), .ZN(n403) );
  XNOR2_X2 U554 ( .A(n763), .B(G146), .ZN(n528) );
  XNOR2_X2 U555 ( .A(n404), .B(n529), .ZN(n567) );
  NAND2_X1 U556 ( .A1(n609), .A2(n559), .ZN(n405) );
  NAND2_X1 U557 ( .A1(n589), .A2(n407), .ZN(n406) );
  NAND2_X1 U558 ( .A1(n777), .A2(KEYINPUT44), .ZN(n410) );
  NAND2_X1 U559 ( .A1(n415), .A2(n414), .ZN(n639) );
  XNOR2_X1 U560 ( .A(n417), .B(n416), .ZN(n415) );
  NAND2_X1 U561 ( .A1(n418), .A2(n369), .ZN(n417) );
  XNOR2_X1 U562 ( .A(n635), .B(n419), .ZN(n418) );
  INV_X1 U563 ( .A(KEYINPUT85), .ZN(n419) );
  XNOR2_X2 U564 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n422) );
  INV_X1 U565 ( .A(n633), .ZN(n426) );
  INV_X1 U566 ( .A(n665), .ZN(n669) );
  NAND2_X1 U567 ( .A1(n665), .A2(n687), .ZN(n611) );
  NAND2_X1 U568 ( .A1(n429), .A2(n427), .ZN(n433) );
  INV_X1 U569 ( .A(n744), .ZN(n428) );
  NAND2_X1 U570 ( .A1(n744), .A2(n370), .ZN(n432) );
  XNOR2_X1 U571 ( .A(n433), .B(n438), .ZN(G51) );
  XNOR2_X1 U572 ( .A(n528), .B(n434), .ZN(n641) );
  INV_X1 U573 ( .A(KEYINPUT56), .ZN(n438) );
  INV_X1 U574 ( .A(n738), .ZN(n440) );
  NAND2_X1 U575 ( .A1(n589), .A2(n367), .ZN(n441) );
  NAND2_X1 U576 ( .A1(n445), .A2(n444), .ZN(n443) );
  XNOR2_X1 U577 ( .A(n629), .B(n446), .ZN(n445) );
  INV_X1 U578 ( .A(KEYINPUT71), .ZN(n446) );
  XNOR2_X2 U579 ( .A(n564), .B(KEYINPUT67), .ZN(n699) );
  INV_X1 U580 ( .A(n567), .ZN(n450) );
  XNOR2_X1 U581 ( .A(n451), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U582 ( .A1(n452), .A2(n439), .ZN(n451) );
  XNOR2_X2 U583 ( .A(n459), .B(G128), .ZN(n537) );
  XNOR2_X1 U584 ( .A(n606), .B(KEYINPUT39), .ZN(n630) );
  XNOR2_X1 U585 ( .A(n776), .B(KEYINPUT83), .ZN(n627) );
  BUF_X1 U586 ( .A(n585), .Z(n700) );
  INV_X1 U587 ( .A(n586), .ZN(n562) );
  XNOR2_X1 U588 ( .A(G478), .B(KEYINPUT106), .ZN(n465) );
  XNOR2_X1 U589 ( .A(n458), .B(n457), .ZN(n462) );
  INV_X2 U590 ( .A(G143), .ZN(n459) );
  NAND2_X1 U591 ( .A1(G217), .A2(n493), .ZN(n463) );
  NOR2_X1 U592 ( .A1(n743), .A2(G902), .ZN(n464) );
  XOR2_X1 U593 ( .A(n465), .B(n464), .Z(n581) );
  INV_X1 U594 ( .A(n581), .ZN(n571) );
  XNOR2_X1 U595 ( .A(KEYINPUT13), .B(G475), .ZN(n480) );
  INV_X1 U596 ( .A(G146), .ZN(n466) );
  INV_X1 U597 ( .A(n469), .ZN(n775) );
  NAND2_X1 U598 ( .A1(n482), .A2(G214), .ZN(n471) );
  XNOR2_X1 U599 ( .A(n472), .B(n471), .ZN(n476) );
  XNOR2_X1 U600 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U601 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U602 ( .A(KEYINPUT102), .B(n582), .ZN(n570) );
  XOR2_X1 U603 ( .A(G113), .B(KEYINPUT5), .Z(n484) );
  NAND2_X1 U604 ( .A1(n482), .A2(G210), .ZN(n483) );
  XNOR2_X1 U605 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U606 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n488) );
  XNOR2_X1 U607 ( .A(n488), .B(n487), .ZN(n750) );
  XNOR2_X1 U608 ( .A(n489), .B(G101), .ZN(n525) );
  XNOR2_X1 U609 ( .A(n750), .B(n525), .ZN(n540) );
  NAND2_X1 U610 ( .A1(n641), .A2(n520), .ZN(n490) );
  INV_X1 U611 ( .A(G472), .ZN(n640) );
  INV_X1 U612 ( .A(KEYINPUT6), .ZN(n491) );
  XNOR2_X1 U613 ( .A(n492), .B(G137), .ZN(n501) );
  INV_X1 U614 ( .A(n494), .ZN(n496) );
  XNOR2_X1 U615 ( .A(KEYINPUT95), .B(KEYINPUT75), .ZN(n495) );
  XNOR2_X1 U616 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U617 ( .A(n497), .ZN(n498) );
  NOR2_X2 U618 ( .A1(n745), .A2(G902), .ZN(n509) );
  XOR2_X1 U619 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n507) );
  INV_X1 U620 ( .A(KEYINPUT15), .ZN(n503) );
  XNOR2_X1 U621 ( .A(n504), .B(n503), .ZN(n548) );
  INV_X1 U622 ( .A(n548), .ZN(n505) );
  NAND2_X1 U623 ( .A1(n505), .A2(G234), .ZN(n506) );
  XNOR2_X2 U624 ( .A(n509), .B(n508), .ZN(n695) );
  XNOR2_X1 U625 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U626 ( .A1(G952), .A2(n512), .ZN(n714) );
  NOR2_X1 U627 ( .A1(n714), .A2(G953), .ZN(n556) );
  NAND2_X1 U628 ( .A1(n512), .A2(G902), .ZN(n513) );
  XOR2_X1 U629 ( .A(KEYINPUT94), .B(n513), .Z(n555) );
  NAND2_X1 U630 ( .A1(G953), .A2(n555), .ZN(n514) );
  NOR2_X1 U631 ( .A1(G900), .A2(n514), .ZN(n515) );
  NOR2_X1 U632 ( .A1(n556), .A2(n515), .ZN(n602) );
  NOR2_X1 U633 ( .A1(n695), .A2(n602), .ZN(n518) );
  NAND2_X1 U634 ( .A1(G221), .A2(n516), .ZN(n517) );
  XOR2_X1 U635 ( .A(KEYINPUT21), .B(n517), .Z(n694) );
  NAND2_X1 U636 ( .A1(n518), .A2(n694), .ZN(n598) );
  NOR2_X1 U637 ( .A1(n576), .A2(n598), .ZN(n521) );
  NAND2_X1 U638 ( .A1(n520), .A2(n519), .ZN(n549) );
  XOR2_X1 U639 ( .A(KEYINPUT108), .B(n614), .Z(n530) );
  XNOR2_X1 U640 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U641 ( .A(n525), .B(n524), .Z(n527) );
  NAND2_X1 U642 ( .A1(G227), .A2(n769), .ZN(n526) );
  XNOR2_X1 U643 ( .A(KEYINPUT72), .B(G469), .ZN(n529) );
  NAND2_X1 U644 ( .A1(n530), .A2(n563), .ZN(n531) );
  XNOR2_X1 U645 ( .A(n531), .B(KEYINPUT43), .ZN(n553) );
  NAND2_X1 U646 ( .A1(n769), .A2(G224), .ZN(n533) );
  XNOR2_X1 U647 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U648 ( .A(n539), .B(n538), .ZN(n541) );
  XNOR2_X1 U649 ( .A(n541), .B(n540), .ZN(n547) );
  XOR2_X1 U650 ( .A(n542), .B(n543), .Z(n546) );
  XNOR2_X1 U651 ( .A(n544), .B(KEYINPUT16), .ZN(n545) );
  XNOR2_X1 U652 ( .A(n546), .B(n545), .ZN(n752) );
  XNOR2_X1 U653 ( .A(n547), .B(n752), .ZN(n737) );
  NAND2_X1 U654 ( .A1(n737), .A2(n505), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n549), .A2(G210), .ZN(n550) );
  INV_X1 U656 ( .A(n358), .ZN(n622) );
  AND2_X1 U657 ( .A1(n553), .A2(n622), .ZN(n632) );
  XOR2_X1 U658 ( .A(n632), .B(G140), .Z(G42) );
  NOR2_X1 U659 ( .A1(G898), .A2(n769), .ZN(n753) );
  NAND2_X1 U660 ( .A1(n555), .A2(n753), .ZN(n558) );
  INV_X1 U661 ( .A(n556), .ZN(n557) );
  NAND2_X1 U662 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U663 ( .A1(n581), .A2(n582), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n599), .A2(n694), .ZN(n560) );
  INV_X1 U665 ( .A(n695), .ZN(n586) );
  XNOR2_X1 U666 ( .A(n384), .B(G101), .ZN(G3) );
  NOR2_X1 U667 ( .A1(n575), .A2(n698), .ZN(n705) );
  NAND2_X1 U668 ( .A1(n565), .A2(n705), .ZN(n566) );
  XNOR2_X1 U669 ( .A(n566), .B(KEYINPUT31), .ZN(n674) );
  NAND2_X1 U670 ( .A1(n604), .A2(n698), .ZN(n568) );
  NOR2_X1 U671 ( .A1(n385), .A2(n568), .ZN(n658) );
  NOR2_X1 U672 ( .A1(n571), .A2(n570), .ZN(n673) );
  OR2_X1 U673 ( .A1(n673), .A2(n671), .ZN(n687) );
  NAND2_X1 U674 ( .A1(n572), .A2(n687), .ZN(n573) );
  XNOR2_X1 U675 ( .A(n575), .B(KEYINPUT107), .ZN(n578) );
  INV_X1 U676 ( .A(n576), .ZN(n577) );
  NAND2_X1 U677 ( .A1(n582), .A2(n581), .ZN(n621) );
  INV_X1 U678 ( .A(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U679 ( .A1(n383), .A2(n590), .ZN(n594) );
  NOR2_X1 U680 ( .A1(n563), .A2(n562), .ZN(n584) );
  NAND2_X1 U681 ( .A1(n586), .A2(n698), .ZN(n587) );
  NOR2_X1 U682 ( .A1(n700), .A2(n587), .ZN(n588) );
  NAND2_X1 U683 ( .A1(n589), .A2(n588), .ZN(n663) );
  NAND2_X1 U684 ( .A1(n778), .A2(n663), .ZN(n592) );
  NAND2_X1 U685 ( .A1(KEYINPUT88), .A2(n590), .ZN(n591) );
  XNOR2_X1 U686 ( .A(n592), .B(n591), .ZN(n593) );
  NAND2_X1 U687 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U688 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X2 U689 ( .A(n597), .B(KEYINPUT45), .ZN(n636) );
  XOR2_X1 U690 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n601) );
  INV_X1 U691 ( .A(n599), .ZN(n685) );
  INV_X1 U692 ( .A(KEYINPUT38), .ZN(n600) );
  XNOR2_X1 U693 ( .A(n358), .B(n600), .ZN(n683) );
  NAND2_X1 U694 ( .A1(n683), .A2(n682), .ZN(n689) );
  INV_X1 U695 ( .A(n602), .ZN(n620) );
  AND2_X1 U696 ( .A1(n620), .A2(n683), .ZN(n605) );
  NAND2_X1 U697 ( .A1(n605), .A2(n619), .ZN(n606) );
  NOR2_X1 U698 ( .A1(n774), .A2(n779), .ZN(n608) );
  INV_X1 U699 ( .A(KEYINPUT76), .ZN(n613) );
  NOR2_X1 U700 ( .A1(n613), .A2(KEYINPUT47), .ZN(n612) );
  NAND2_X1 U701 ( .A1(n613), .A2(KEYINPUT47), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n615), .A2(n700), .ZN(n676) );
  AND2_X1 U703 ( .A1(n616), .A2(n676), .ZN(n617) );
  AND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n624) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n630), .A2(n673), .ZN(n679) );
  INV_X1 U708 ( .A(n679), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n636), .A2(n634), .ZN(n635) );
  INV_X1 U711 ( .A(KEYINPUT2), .ZN(n719) );
  BUF_X1 U712 ( .A(n636), .Z(n637) );
  INV_X1 U713 ( .A(n765), .ZN(n638) );
  XNOR2_X2 U714 ( .A(n639), .B(KEYINPUT64), .ZN(n742) );
  NOR2_X1 U715 ( .A1(n742), .A2(n640), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(n645) );
  INV_X1 U717 ( .A(G952), .ZN(n644) );
  XNOR2_X1 U718 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n647), .B(n646), .ZN(G57) );
  INV_X1 U720 ( .A(G475), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n742), .A2(n648), .ZN(n652) );
  XOR2_X1 U722 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n649) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U724 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(G60) );
  NAND2_X1 U726 ( .A1(n658), .A2(n671), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT112), .ZN(n657) );
  XNOR2_X1 U728 ( .A(G104), .B(n657), .ZN(G6) );
  XOR2_X1 U729 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n660) );
  NAND2_X1 U730 ( .A1(n658), .A2(n673), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n660), .B(n659), .ZN(n662) );
  XOR2_X1 U732 ( .A(G107), .B(KEYINPUT27), .Z(n661) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(G9) );
  XNOR2_X1 U734 ( .A(G110), .B(KEYINPUT114), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n664), .B(n663), .ZN(G12) );
  XOR2_X1 U736 ( .A(G128), .B(KEYINPUT29), .Z(n667) );
  NAND2_X1 U737 ( .A1(n665), .A2(n673), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n667), .B(n666), .ZN(G30) );
  OR2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n670), .B(G146), .ZN(G48) );
  NAND2_X1 U741 ( .A1(n671), .A2(n674), .ZN(n672) );
  XNOR2_X1 U742 ( .A(G113), .B(n672), .ZN(G15) );
  NAND2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n675), .B(G116), .ZN(G18) );
  XNOR2_X1 U745 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U747 ( .A(G125), .B(n678), .ZN(G27) );
  XNOR2_X1 U748 ( .A(G134), .B(KEYINPUT116), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(G36) );
  XOR2_X1 U750 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n734) );
  INV_X1 U751 ( .A(n715), .ZN(n693) );
  NOR2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U754 ( .A(KEYINPUT119), .B(n686), .Z(n691) );
  INV_X1 U755 ( .A(n687), .ZN(n688) );
  NOR2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n711) );
  NOR2_X1 U759 ( .A1(n562), .A2(n694), .ZN(n696) );
  XNOR2_X1 U760 ( .A(n696), .B(KEYINPUT49), .ZN(n697) );
  NAND2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n703) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U763 ( .A(n701), .B(KEYINPUT50), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U766 ( .A(KEYINPUT51), .B(n706), .Z(n707) );
  XNOR2_X1 U767 ( .A(KEYINPUT117), .B(n707), .ZN(n708) );
  NAND2_X1 U768 ( .A1(n708), .A2(n716), .ZN(n709) );
  XOR2_X1 U769 ( .A(KEYINPUT118), .B(n709), .Z(n710) );
  NOR2_X1 U770 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U771 ( .A(n712), .B(KEYINPUT52), .ZN(n713) );
  NOR2_X1 U772 ( .A1(n714), .A2(n713), .ZN(n731) );
  NAND2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n729) );
  XNOR2_X1 U774 ( .A(KEYINPUT82), .B(KEYINPUT2), .ZN(n717) );
  NOR2_X1 U775 ( .A1(n638), .A2(n717), .ZN(n718) );
  XOR2_X1 U776 ( .A(KEYINPUT84), .B(n718), .Z(n727) );
  INV_X1 U777 ( .A(KEYINPUT82), .ZN(n720) );
  NOR2_X1 U778 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n637), .A2(n721), .ZN(n722) );
  NOR2_X1 U780 ( .A1(n723), .A2(n722), .ZN(n725) );
  NOR2_X1 U781 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n724) );
  OR2_X1 U782 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U783 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U785 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U786 ( .A1(n732), .A2(n769), .ZN(n733) );
  XNOR2_X1 U787 ( .A(n734), .B(n733), .ZN(G75) );
  INV_X1 U788 ( .A(n742), .ZN(n744) );
  XOR2_X1 U789 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n735) );
  XNOR2_X1 U790 ( .A(n735), .B(KEYINPUT89), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n382), .B(n736), .ZN(n738) );
  XOR2_X1 U792 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n739) );
  NOR2_X1 U793 ( .A1(n749), .A2(n741), .ZN(G54) );
  NAND2_X1 U794 ( .A1(n744), .A2(G217), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n360), .B(KEYINPUT124), .ZN(n746) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U797 ( .A1(n749), .A2(n748), .ZN(G66) );
  XOR2_X1 U798 ( .A(G101), .B(n750), .Z(n751) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(n754) );
  NOR2_X1 U800 ( .A1(n754), .A2(n753), .ZN(n761) );
  NAND2_X1 U801 ( .A1(n637), .A2(n769), .ZN(n759) );
  XOR2_X1 U802 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n756) );
  NAND2_X1 U803 ( .A1(G224), .A2(G953), .ZN(n755) );
  XNOR2_X1 U804 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U805 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U807 ( .A(n761), .B(n760), .ZN(G69) );
  XOR2_X1 U808 ( .A(n763), .B(n762), .Z(n764) );
  XOR2_X1 U809 ( .A(KEYINPUT126), .B(n764), .Z(n767) );
  XOR2_X1 U810 ( .A(n767), .B(n765), .Z(n766) );
  NAND2_X1 U811 ( .A1(n766), .A2(n769), .ZN(n772) );
  XOR2_X1 U812 ( .A(G227), .B(n767), .Z(n768) );
  NOR2_X1 U813 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U814 ( .A1(G900), .A2(n770), .ZN(n771) );
  NAND2_X1 U815 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U816 ( .A(KEYINPUT127), .B(n773), .ZN(G72) );
  XOR2_X1 U817 ( .A(G137), .B(n774), .Z(G39) );
  XNOR2_X1 U818 ( .A(n776), .B(n775), .ZN(G45) );
  XOR2_X1 U819 ( .A(n383), .B(G122), .Z(G24) );
  XNOR2_X1 U820 ( .A(G119), .B(n778), .ZN(G21) );
  XOR2_X1 U821 ( .A(n779), .B(G131), .Z(G33) );
endmodule

