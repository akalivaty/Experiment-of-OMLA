//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(new_n218), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  NOR2_X1   g0035(.A1(new_n201), .A2(new_n202), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(new_n203), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT64), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G97), .B(G107), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  XNOR2_X1  g0045(.A(KEYINPUT3), .B(G33), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT7), .ZN(new_n247));
  NOR3_X1   g0047(.A1(new_n246), .A2(new_n247), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(KEYINPUT7), .B1(new_n253), .B2(new_n213), .ZN(new_n254));
  OAI21_X1  g0054(.A(G68), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n217), .A2(new_n201), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G58), .A2(G68), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G159), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n255), .A2(KEYINPUT16), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT16), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n247), .B1(new_n246), .B2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n201), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n267), .B2(new_n261), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n212), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT68), .B1(new_n269), .B2(new_n212), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n263), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n274), .A2(new_n213), .A3(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n269), .A2(new_n212), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n212), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n213), .A2(G1), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n280), .A2(new_n283), .B1(new_n275), .B2(new_n281), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n273), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n273), .A2(KEYINPUT74), .A3(new_n284), .ZN(new_n288));
  AND2_X1   g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  OAI21_X1  g0089(.A(G274), .B1(new_n289), .B2(new_n212), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT65), .ZN(new_n294));
  INV_X1    g0094(.A(G1), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G41), .B2(G45), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT65), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n290), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G1), .A3(G13), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G232), .A3(new_n296), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT75), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G274), .ZN(new_n305));
  INV_X1    g0105(.A(new_n212), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n300), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n291), .A2(new_n292), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT65), .B1(new_n308), .B2(new_n295), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n296), .A2(new_n297), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT75), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n302), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G1698), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT66), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT66), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(new_n246), .A3(G223), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n246), .A2(G226), .A3(G1698), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G87), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n301), .ZN(new_n324));
  AOI21_X1  g0124(.A(G179), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n299), .A2(new_n303), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n314), .A2(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n287), .A2(new_n288), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT76), .A2(KEYINPUT18), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n326), .A2(new_n304), .A3(new_n313), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(G200), .B1(new_n326), .B2(new_n327), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n273), .B(new_n284), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n337), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n335), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(KEYINPUT77), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n343), .A2(new_n273), .A3(new_n284), .A4(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n331), .A2(new_n333), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(KEYINPUT76), .A2(KEYINPUT18), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n333), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n287), .A2(new_n288), .A3(new_n330), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(KEYINPUT78), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G226), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n301), .A2(new_n296), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n311), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n246), .A2(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(G223), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n356), .A2(new_n357), .B1(new_n202), .B2(new_n246), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n319), .A2(new_n246), .ZN(new_n359));
  INV_X1    g0159(.A(G222), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT67), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n301), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OR3_X1    g0164(.A1(new_n358), .A2(new_n361), .A3(new_n363), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n355), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n329), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n282), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n280), .A2(G50), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n213), .A2(G33), .ZN(new_n373));
  INV_X1    g0173(.A(G150), .ZN(new_n374));
  INV_X1    g0174(.A(new_n259), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n281), .A2(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(G50), .A2(G58), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n213), .B1(new_n377), .B2(new_n201), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n272), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n274), .A2(G1), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G20), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n372), .B(new_n379), .C1(G50), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n368), .A2(new_n370), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT69), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n368), .A2(KEYINPUT69), .A3(new_n370), .A4(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n366), .A2(G190), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT71), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n382), .B(KEYINPUT9), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G200), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n366), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT10), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n390), .A2(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n367), .A2(G200), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT10), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .A4(new_n388), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n253), .A2(G107), .ZN(new_n400));
  INV_X1    g0200(.A(G238), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n400), .B1(new_n356), .B2(new_n401), .C1(new_n218), .C2(new_n359), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n324), .ZN(new_n403));
  INV_X1    g0203(.A(new_n354), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n299), .B1(G244), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n329), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n280), .A2(G77), .A3(new_n371), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT15), .B(G87), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT70), .ZN(new_n410));
  OR3_X1    g0210(.A1(new_n409), .A2(new_n410), .A3(new_n373), .ZN(new_n411));
  XOR2_X1   g0211(.A(KEYINPUT8), .B(G58), .Z(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n410), .B1(new_n409), .B2(new_n373), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n278), .A2(new_n279), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n408), .B1(G77), .B2(new_n381), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n407), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n406), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n369), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n417), .B1(new_n419), .B2(G190), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n392), .B2(new_n419), .ZN(new_n423));
  AND4_X1   g0223(.A1(new_n387), .A2(new_n399), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n331), .A2(new_n333), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n341), .A2(new_n347), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n351), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT78), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n280), .A2(G68), .A3(new_n371), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT72), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n201), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n202), .B2(new_n373), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n272), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT11), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n275), .A2(new_n201), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT12), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n272), .A2(new_n433), .A3(KEYINPUT11), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n431), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT66), .B(G1698), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n442), .A2(new_n353), .B1(new_n218), .B2(new_n315), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(new_n246), .B1(G33), .B2(G97), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n301), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n311), .B1(new_n401), .B2(new_n354), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT13), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n299), .B1(G238), .B2(new_n404), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT13), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n448), .B(new_n449), .C1(new_n301), .C2(new_n444), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n441), .B1(new_n451), .B2(new_n334), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n392), .B1(new_n447), .B2(new_n450), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n447), .A2(new_n450), .A3(G179), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT73), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n447), .A2(new_n450), .A3(KEYINPUT73), .A4(G179), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n451), .A2(G169), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT14), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT14), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n451), .A2(new_n462), .A3(G169), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n441), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n454), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND4_X1   g0266(.A1(new_n352), .A2(new_n424), .A3(new_n429), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT85), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n250), .A2(new_n252), .A3(G257), .A4(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT84), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT84), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n246), .A2(new_n471), .A3(G257), .A4(G1698), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n319), .A2(new_n246), .A3(G250), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G294), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n470), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n324), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n295), .A2(G45), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n480), .A2(G264), .A3(new_n301), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n307), .A2(new_n479), .A3(new_n477), .ZN(new_n483));
  AND4_X1   g0283(.A1(G179), .A2(new_n476), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n475), .B2(new_n324), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n329), .B1(new_n485), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n468), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(G179), .A3(new_n483), .ZN(new_n488));
  INV_X1    g0288(.A(new_n483), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n489), .B(new_n481), .C1(new_n475), .C2(new_n324), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n488), .B(KEYINPUT85), .C1(new_n490), .C2(new_n329), .ZN(new_n491));
  INV_X1    g0291(.A(G107), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n492), .A2(KEYINPUT23), .A3(G20), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT23), .B1(new_n492), .B2(G20), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n493), .A2(new_n494), .B1(G20), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n246), .A2(new_n213), .A3(G87), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT22), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT22), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n246), .A2(new_n499), .A3(new_n213), .A4(G87), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT24), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(KEYINPUT24), .B(new_n496), .C1(new_n498), .C2(new_n500), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n272), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n213), .A2(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n380), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g0308(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n509));
  AND4_X1   g0309(.A1(new_n380), .A2(new_n507), .A3(new_n509), .A4(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n295), .A2(G33), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n381), .B(new_n511), .C1(new_n270), .C2(new_n271), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI211_X1 g0313(.A(new_n508), .B(new_n510), .C1(new_n513), .C2(G107), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n487), .A2(new_n491), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT86), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n487), .A2(new_n491), .A3(KEYINPUT86), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n490), .A2(G190), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n485), .A2(new_n483), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n520), .A2(new_n522), .A3(new_n505), .A4(new_n514), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n518), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT87), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT87), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n518), .A2(new_n526), .A3(new_n519), .A4(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n380), .A2(G20), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n269), .A2(new_n212), .B1(G20), .B2(new_n529), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(new_n213), .C1(G33), .C2(new_n219), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n531), .A2(KEYINPUT20), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT20), .B1(new_n531), .B2(new_n533), .ZN(new_n535));
  OAI221_X1 g0335(.A(new_n530), .B1(new_n534), .B2(new_n535), .C1(new_n529), .C2(new_n512), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n246), .A2(G264), .A3(G1698), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n253), .A2(G303), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n359), .C2(new_n220), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n324), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n480), .A2(G270), .A3(new_n301), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n483), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n536), .B1(new_n542), .B2(G200), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n334), .B2(new_n542), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n536), .A3(G169), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n541), .A2(new_n483), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n539), .B2(new_n324), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n536), .A3(G179), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n542), .A2(new_n536), .A3(KEYINPUT21), .A4(G169), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n544), .A2(new_n547), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT82), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n319), .A2(new_n246), .A3(G244), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n250), .A2(new_n252), .A3(G250), .A4(G1698), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n557), .A2(new_n532), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n319), .A2(new_n246), .A3(KEYINPUT4), .A4(G244), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n324), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n480), .A2(G257), .A3(new_n301), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n483), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n565), .A2(new_n219), .A3(G107), .ZN(new_n566));
  XNOR2_X1  g0366(.A(G97), .B(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n568), .A2(new_n213), .B1(new_n202), .B2(new_n375), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n492), .B1(new_n265), .B2(new_n266), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n272), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n512), .A2(G97), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n275), .A2(G97), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(KEYINPUT79), .B(new_n574), .C1(new_n512), .C2(G97), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n562), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n560), .B2(new_n324), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(G190), .A3(new_n483), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n564), .A2(new_n571), .A3(new_n578), .A4(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n571), .B1(new_n576), .B2(new_n577), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n561), .A2(new_n369), .A3(new_n483), .A4(new_n562), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n489), .B(new_n579), .C1(new_n560), .C2(new_n324), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(G169), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n250), .A2(new_n252), .A3(new_n213), .A4(G68), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n373), .B2(new_n219), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G97), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n213), .B1(new_n592), .B2(new_n589), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT80), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(KEYINPUT80), .B(new_n213), .C1(new_n592), .C2(new_n589), .ZN(new_n596));
  OR2_X1    g0396(.A1(KEYINPUT81), .A2(G87), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G97), .A2(G107), .ZN(new_n598));
  NAND2_X1  g0398(.A1(KEYINPUT81), .A2(G87), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n416), .B1(new_n591), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G87), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n512), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n409), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n381), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n602), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n250), .A2(new_n252), .A3(G244), .A4(G1698), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n495), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n319), .A2(new_n246), .A3(G238), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n301), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n301), .A2(G250), .A3(new_n478), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n290), .B2(new_n478), .ZN(new_n613));
  OAI21_X1  g0413(.A(G200), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n495), .A3(new_n608), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(new_n324), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G190), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n607), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n591), .A2(new_n601), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n272), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n513), .A2(new_n605), .ZN(new_n621));
  INV_X1    g0421(.A(new_n606), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n329), .B1(new_n611), .B2(new_n613), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n616), .A2(new_n369), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n553), .B1(new_n587), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n618), .A2(new_n626), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n582), .A2(new_n629), .A3(KEYINPUT82), .A4(new_n586), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n552), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n467), .A2(new_n528), .A3(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n586), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(KEYINPUT89), .A3(new_n629), .A4(KEYINPUT26), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT88), .B1(new_n616), .B2(new_n392), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n636), .B(G200), .C1(new_n611), .C2(new_n613), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n635), .A2(new_n607), .A3(new_n637), .A4(new_n617), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(new_n626), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(new_n523), .A3(new_n586), .A4(new_n582), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n641));
  INV_X1    g0441(.A(new_n486), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n488), .B1(new_n505), .B2(new_n514), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n626), .B(new_n634), .C1(new_n640), .C2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n584), .ZN(new_n646));
  AOI21_X1  g0446(.A(G169), .B1(new_n580), .B2(new_n483), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n629), .A2(new_n648), .A3(KEYINPUT26), .A4(new_n583), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n638), .A2(new_n626), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n586), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n467), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n426), .ZN(new_n657));
  INV_X1    g0457(.A(new_n421), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n453), .B2(new_n452), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n464), .A2(new_n465), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT18), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n285), .A2(new_n330), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n285), .B2(new_n330), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n399), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n387), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n656), .A2(new_n668), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n380), .A2(new_n213), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT27), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n671), .A2(KEYINPUT90), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT90), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n670), .B2(KEYINPUT27), .ZN(new_n675));
  OAI221_X1 g0475(.A(G213), .B1(KEYINPUT27), .B2(new_n670), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G343), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n515), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT91), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n525), .B2(new_n527), .ZN(new_n682));
  INV_X1    g0482(.A(new_n516), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n679), .ZN(new_n684));
  INV_X1    g0484(.A(new_n641), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n679), .A2(new_n536), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n544), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n685), .A2(new_n679), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n682), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n643), .B2(new_n678), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n207), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G1), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n597), .A2(new_n599), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(new_n529), .A3(new_n598), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n699), .A2(new_n701), .B1(new_n210), .B2(new_n698), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n563), .A2(new_n705), .A3(new_n521), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT93), .B(new_n483), .C1(new_n580), .C2(new_n485), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n549), .A2(G179), .A3(new_n616), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n580), .A2(new_n549), .A3(G179), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n485), .A2(new_n616), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT92), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n485), .A2(KEYINPUT92), .A3(new_n616), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n709), .B1(new_n715), .B2(KEYINPUT30), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n717), .B(new_n710), .C1(new_n713), .C2(new_n714), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n679), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI211_X1 g0521(.A(new_n552), .B(new_n679), .C1(new_n628), .C2(new_n630), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n528), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(new_n720), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n704), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n655), .A2(new_n678), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n626), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n651), .A2(new_n586), .A3(new_n650), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(KEYINPUT94), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n639), .A2(new_n633), .A3(KEYINPUT26), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT94), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n650), .B1(new_n586), .B2(new_n627), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n518), .A2(new_n519), .A3(new_n685), .ZN(new_n737));
  INV_X1    g0537(.A(new_n640), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n679), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT29), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n725), .B1(new_n728), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n703), .B1(new_n742), .B2(G1), .ZN(G364));
  NOR2_X1   g0543(.A1(new_n688), .A2(G330), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT95), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n274), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n295), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OR3_X1    g0548(.A1(new_n697), .A2(new_n748), .A3(KEYINPUT96), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT96), .B1(new_n697), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n689), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n751), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n696), .A2(new_n253), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G355), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G116), .B2(new_n207), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n241), .A2(G45), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n696), .A2(new_n246), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n292), .B2(new_n211), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n756), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n212), .B1(G20), .B2(new_n329), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n753), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n765), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n334), .A2(new_n392), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n213), .A2(G179), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n253), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n213), .A2(new_n369), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G190), .A3(new_n392), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n770), .A2(new_n775), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n777), .A2(G322), .B1(new_n779), .B2(G326), .ZN(new_n780));
  INV_X1    g0580(.A(G329), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n771), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n334), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n213), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n774), .B(new_n784), .C1(G294), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT97), .ZN(new_n789));
  AND3_X1   g0589(.A1(new_n775), .A2(new_n789), .A3(new_n782), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n775), .B2(new_n782), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G311), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n392), .A2(G190), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n771), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT99), .Z(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G283), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n775), .A2(new_n795), .A3(KEYINPUT100), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(KEYINPUT100), .B1(new_n775), .B2(new_n795), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT101), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n788), .A2(new_n794), .A3(new_n798), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n783), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT98), .B(KEYINPUT32), .Z(new_n810));
  XNOR2_X1  g0610(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G77), .B2(new_n793), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n246), .B1(new_n700), .B2(new_n772), .ZN(new_n813));
  INV_X1    g0613(.A(G50), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n776), .A2(new_n217), .B1(new_n778), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(G97), .C2(new_n787), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n797), .A2(G107), .B1(new_n803), .B2(G68), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n812), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n769), .B1(new_n807), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n768), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n764), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n688), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n752), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  AND3_X1   g0624(.A1(new_n418), .A2(new_n420), .A3(new_n678), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n679), .A2(new_n417), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n423), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n825), .B1(new_n827), .B2(new_n421), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n726), .B(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n725), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n753), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n725), .B2(new_n829), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n769), .A2(new_n763), .ZN(new_n835));
  INV_X1    g0635(.A(G311), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n253), .B1(new_n783), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n772), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n777), .A2(G294), .B1(new_n838), .B2(G107), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n773), .B2(new_n778), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n837), .B(new_n840), .C1(G97), .C2(new_n787), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n797), .A2(G87), .B1(new_n793), .B2(G116), .ZN(new_n842));
  INV_X1    g0642(.A(G283), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n802), .A2(KEYINPUT102), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n802), .A2(KEYINPUT102), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n777), .A2(G143), .B1(new_n779), .B2(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n849), .B1(new_n792), .B2(new_n808), .C1(new_n374), .C2(new_n802), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT34), .Z(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n246), .B1(new_n783), .B2(new_n852), .C1(new_n786), .C2(new_n217), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n797), .A2(G68), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n814), .B2(new_n772), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT103), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n848), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT104), .Z(new_n860));
  OAI221_X1 g0660(.A(new_n753), .B1(G77), .B2(new_n835), .C1(new_n860), .C2(new_n769), .ZN(new_n861));
  INV_X1    g0661(.A(new_n828), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n762), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT105), .Z(new_n864));
  NOR2_X1   g0664(.A1(new_n834), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n746), .A2(new_n295), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n528), .A2(new_n722), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n719), .A2(KEYINPUT110), .A3(new_n720), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT110), .B1(new_n719), .B2(new_n720), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n721), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n441), .A2(new_n678), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n466), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n465), .B(new_n679), .C1(new_n464), .C2(new_n454), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n828), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n676), .B1(new_n273), .B2(new_n284), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n348), .B2(new_n351), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n338), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n287), .A2(new_n288), .A3(new_n677), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n331), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n285), .A2(new_n330), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n338), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n890), .B2(new_n882), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n881), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT107), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n427), .A2(new_n882), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n888), .A2(new_n891), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n873), .B(new_n880), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n886), .A2(new_n331), .A3(new_n887), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n889), .A2(new_n338), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n885), .B1(new_n904), .B2(new_n887), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT109), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n273), .A2(KEYINPUT74), .A3(new_n284), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT74), .B1(new_n273), .B2(new_n284), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(new_n676), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n909), .B2(new_n890), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT109), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n911), .A3(new_n888), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n887), .B1(new_n665), .B2(new_n426), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n906), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n881), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n897), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n917), .A2(new_n873), .A3(new_n880), .A4(KEYINPUT40), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n902), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n467), .A2(new_n873), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(G330), .A3(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT111), .Z(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n910), .A2(new_n888), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n913), .B1(new_n927), .B2(KEYINPUT109), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n928), .B2(new_n912), .ZN(new_n929));
  AOI221_X4 g0729(.A(new_n881), .B1(new_n888), .B2(new_n891), .C1(new_n427), .C2(new_n882), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n464), .A2(new_n465), .A3(new_n678), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT108), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n877), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n874), .B(new_n454), .C1(new_n464), .C2(new_n465), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n678), .B(new_n828), .C1(new_n645), .C2(new_n654), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n825), .B(KEYINPUT106), .Z(new_n940));
  AOI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n898), .B2(new_n899), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n666), .A2(new_n676), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n935), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n467), .A2(new_n728), .A3(new_n741), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n668), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n867), .B1(new_n925), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n925), .B2(new_n947), .ZN(new_n949));
  INV_X1    g0749(.A(new_n568), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT35), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT35), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n951), .A2(G116), .A3(new_n214), .A4(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT36), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n256), .A2(new_n210), .A3(new_n202), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n201), .A2(G50), .ZN(new_n956));
  OAI211_X1 g0756(.A(G1), .B(new_n274), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n954), .A3(new_n957), .ZN(G367));
  NAND2_X1  g0758(.A1(new_n679), .A2(new_n583), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(new_n582), .A3(new_n586), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n586), .B2(new_n678), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n693), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n518), .B2(new_n519), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n678), .B1(new_n964), .B2(new_n633), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(KEYINPUT113), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(KEYINPUT113), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n626), .A2(new_n678), .A3(new_n607), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT112), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT112), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n678), .A2(new_n607), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n972), .B(new_n973), .C1(new_n651), .C2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT43), .Z(new_n976));
  OR3_X1    g0776(.A1(new_n968), .A2(new_n969), .A3(new_n976), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n968), .A2(new_n969), .B1(KEYINPUT43), .B2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n690), .A2(new_n961), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n697), .B(KEYINPUT41), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n694), .A2(new_n961), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT45), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n694), .A2(new_n961), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n690), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n691), .A3(new_n986), .ZN(new_n989));
  INV_X1    g0789(.A(new_n692), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n693), .B1(new_n684), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(new_n689), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n988), .A2(new_n742), .A3(new_n989), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n982), .B1(new_n993), .B2(new_n742), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n981), .B1(new_n994), .B2(new_n748), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n772), .A2(new_n529), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT46), .ZN(new_n997));
  INV_X1    g0797(.A(new_n847), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(new_n998), .B2(G294), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT114), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(KEYINPUT114), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n253), .B1(new_n796), .B2(new_n219), .C1(new_n786), .C2(new_n492), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n777), .A2(G303), .B1(new_n779), .B2(G311), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n783), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1002), .B(new_n1005), .C1(G283), .C2(new_n793), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1000), .A2(new_n1001), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT115), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(KEYINPUT115), .ZN(new_n1010));
  INV_X1    g0810(.A(G143), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n246), .B1(new_n778), .B2(new_n1011), .C1(new_n786), .C2(new_n201), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n776), .A2(new_n374), .B1(new_n796), .B2(new_n202), .ZN(new_n1013));
  INV_X1    g0813(.A(G137), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n772), .A2(new_n217), .B1(new_n783), .B2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n814), .B2(new_n792), .C1(new_n847), .C2(new_n808), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT116), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1009), .A2(new_n1010), .A3(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT117), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT47), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n769), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n1021), .B2(new_n1020), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n234), .A2(new_n758), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n767), .B1(new_n696), .B2(new_n605), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n751), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1023), .B(new_n1026), .C1(new_n821), .C2(new_n975), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n995), .A2(new_n1027), .ZN(G387));
  AOI21_X1  g0828(.A(new_n698), .B1(new_n992), .B2(new_n742), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n742), .B2(new_n992), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n231), .A2(new_n292), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1031), .A2(new_n758), .B1(new_n701), .B2(new_n754), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n412), .A2(new_n814), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n1034), .A2(G45), .A3(new_n236), .A4(new_n701), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1032), .A2(new_n1035), .B1(G107), .B2(new_n207), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n751), .B1(new_n1036), .B2(new_n766), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n778), .A2(new_n808), .B1(new_n783), .B2(new_n374), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G50), .B2(new_n777), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n253), .B1(new_n838), .B2(G77), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n409), .C2(new_n786), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n802), .A2(new_n281), .B1(new_n792), .B2(new_n201), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT118), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(G97), .C2(new_n797), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n792), .A2(new_n773), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(KEYINPUT119), .B(G322), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n776), .A2(new_n1004), .B1(new_n778), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1045), .B(new_n1047), .C1(new_n998), .C2(G311), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT48), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(KEYINPUT48), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n787), .A2(G283), .B1(new_n838), .B2(G294), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT49), .ZN(new_n1054));
  INV_X1    g0854(.A(G326), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n253), .B1(new_n783), .B2(new_n1055), .C1(new_n529), .C2(new_n796), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1053), .B2(KEYINPUT49), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1044), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1037), .B1(new_n1058), .B2(new_n769), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n684), .B2(new_n764), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n992), .B2(new_n748), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1030), .A2(new_n1061), .ZN(G393));
  NAND2_X1  g0862(.A1(new_n992), .A2(new_n742), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n989), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n691), .B1(new_n984), .B2(new_n986), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n993), .A3(new_n697), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n961), .A2(new_n821), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n766), .B1(new_n219), .B2(new_n207), .C1(new_n244), .C2(new_n759), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n753), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n847), .A2(new_n773), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n797), .A2(G107), .B1(new_n793), .B2(G294), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n776), .A2(new_n836), .B1(new_n778), .B2(new_n1004), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n253), .B1(new_n783), .B2(new_n1046), .C1(new_n843), .C2(new_n772), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G116), .B2(new_n787), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n847), .A2(new_n814), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n797), .A2(G87), .B1(new_n793), .B2(new_n412), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n246), .B1(new_n783), .B2(new_n1011), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n786), .A2(new_n202), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(G68), .C2(new_n838), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n776), .A2(new_n808), .B1(new_n778), .B2(new_n374), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT51), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1080), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1072), .A2(new_n1078), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1071), .B1(new_n1087), .B2(new_n765), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1068), .A2(new_n748), .B1(new_n1069), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1067), .A2(new_n1089), .ZN(G390));
  AOI21_X1  g0890(.A(new_n704), .B1(new_n723), .B2(new_n871), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n880), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n939), .A2(new_n940), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n933), .B1(new_n1094), .B2(new_n878), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n931), .B2(new_n934), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n933), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n929), .B2(new_n930), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n827), .A2(new_n421), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n737), .A2(new_n738), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n731), .A2(new_n735), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n678), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n825), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n938), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1093), .B1(new_n1096), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT39), .B1(new_n916), .B2(new_n897), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n934), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1107), .A2(new_n1108), .B1(new_n941), .B2(new_n933), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n825), .B1(new_n740), .B2(new_n1099), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n917), .B(new_n1097), .C1(new_n1110), .C2(new_n938), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n868), .A2(new_n724), .A3(new_n872), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1112), .A2(G330), .A3(new_n828), .A4(new_n878), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1109), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n762), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n753), .B1(new_n412), .B2(new_n835), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n847), .A2(new_n492), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n783), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n246), .B(new_n1082), .C1(G294), .C2(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n776), .A2(new_n529), .B1(new_n772), .B2(new_n603), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G283), .B2(new_n779), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n793), .A2(G97), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n854), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n847), .A2(new_n1014), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n772), .A2(new_n374), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1128));
  XNOR2_X1  g0928(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n792), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n246), .B1(new_n776), .B2(new_n852), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G159), .B2(new_n787), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  INV_X1    g0934(.A(G125), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n778), .A2(new_n1134), .B1(new_n783), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n796), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(G50), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1129), .A2(new_n1131), .A3(new_n1133), .A4(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1119), .A2(new_n1125), .B1(new_n1126), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1118), .B1(new_n1140), .B2(new_n765), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT121), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1116), .A2(new_n748), .B1(new_n1117), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n704), .B(new_n862), .C1(new_n723), .C2(new_n724), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1092), .B1(new_n1144), .B2(new_n878), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1094), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1113), .A2(new_n1110), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1091), .A2(new_n828), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n938), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n467), .A2(new_n1091), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n945), .A2(new_n1152), .A3(new_n668), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n1115), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n697), .B1(new_n1157), .B2(new_n1116), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1143), .B1(new_n1156), .B2(new_n1158), .ZN(G378));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1153), .B1(new_n1116), .B2(new_n1151), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n902), .A2(G330), .A3(new_n918), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n677), .A2(new_n382), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT124), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n399), .A2(new_n383), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n399), .B2(new_n383), .ZN(new_n1167));
  XOR2_X1   g0967(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OR3_X1    g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT125), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n944), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT38), .B1(new_n895), .B2(new_n896), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT107), .B1(new_n930), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1179), .A2(new_n941), .B1(new_n666), .B2(new_n676), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1173), .B1(new_n1180), .B2(new_n935), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1162), .B1(new_n1175), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n944), .A2(new_n1174), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n902), .A2(G330), .A3(new_n918), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n935), .A3(new_n1173), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1160), .B1(new_n1161), .B2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1094), .A2(new_n1145), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1154), .B1(new_n1189), .B2(new_n1115), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1190), .A2(KEYINPUT57), .A3(new_n1182), .A4(new_n1186), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n697), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1182), .A2(new_n748), .A3(new_n1186), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1170), .A2(new_n762), .A3(new_n1172), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n753), .B1(G50), .B2(new_n835), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n802), .A2(new_n852), .B1(new_n792), .B2(new_n1014), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n779), .A2(G125), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n1134), .B2(new_n776), .C1(new_n772), .C2(new_n1130), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G150), .C2(new_n787), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1137), .A2(G159), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n1120), .C2(G124), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G41), .B(new_n246), .C1(new_n838), .C2(G77), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n217), .B2(new_n796), .C1(new_n843), .C2(new_n783), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT122), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n802), .A2(new_n219), .B1(new_n792), .B2(new_n409), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT123), .Z(new_n1210));
  OAI22_X1  g1010(.A1(new_n776), .A2(new_n492), .B1(new_n778), .B2(new_n529), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G68), .B2(new_n787), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT58), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(G50), .B1(new_n249), .B2(new_n291), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n246), .B2(G41), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1205), .A2(new_n1215), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1195), .B1(new_n1219), .B2(new_n765), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1194), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1193), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1192), .A2(new_n1223), .ZN(G375));
  NAND2_X1  g1024(.A1(new_n938), .A2(new_n762), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n753), .B1(G68), .B2(new_n835), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n847), .A2(new_n529), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n797), .A2(G77), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n793), .A2(G107), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n772), .A2(new_n219), .B1(new_n783), .B2(new_n773), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G294), .B2(new_n779), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n253), .B1(new_n776), .B2(new_n843), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n605), .B2(new_n787), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1228), .A2(new_n1229), .A3(new_n1231), .A4(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n847), .A2(new_n1130), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n246), .B1(new_n796), .B2(new_n217), .C1(new_n786), .C2(new_n814), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n776), .A2(new_n1014), .B1(new_n783), .B2(new_n1134), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n778), .A2(new_n852), .B1(new_n772), .B2(new_n808), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n374), .B2(new_n792), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1227), .A2(new_n1234), .B1(new_n1235), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1226), .B1(new_n1241), .B2(new_n765), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1151), .A2(new_n748), .B1(new_n1225), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n982), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1155), .A2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1243), .B1(new_n1245), .B2(new_n1246), .ZN(G381));
  NOR2_X1   g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n865), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(G390), .A2(G381), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  OR3_X1    g1052(.A1(new_n1252), .A2(G387), .A3(G375), .ZN(G407));
  INV_X1    g1053(.A(G213), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1254), .A2(G343), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G407), .B(G213), .C1(G375), .C2(new_n1256), .ZN(G409));
  AOI21_X1  g1057(.A(new_n823), .B1(new_n1030), .B2(new_n1061), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1248), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G390), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1067), .B(new_n1089), .C1(new_n1248), .C2(new_n1258), .ZN(new_n1261));
  AND4_X1   g1061(.A1(new_n1027), .A2(new_n1260), .A3(new_n995), .A4(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1260), .A2(new_n1261), .B1(new_n995), .B2(new_n1027), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1189), .A2(KEYINPUT60), .A3(new_n1153), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n697), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1246), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1155), .A2(KEYINPUT60), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1267), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1243), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n865), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1246), .B1(KEYINPUT60), .B2(new_n1155), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G384), .B(new_n1243), .C1(new_n1273), .C2(new_n1267), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1255), .A2(G2897), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1184), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1244), .A3(new_n1190), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1222), .B1(new_n1282), .B2(KEYINPUT127), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(new_n1284), .A3(new_n1244), .A4(new_n1190), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1191), .A2(new_n697), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT57), .B1(new_n1281), .B2(new_n1190), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1223), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT126), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1192), .A2(new_n1291), .A3(G378), .A4(new_n1223), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1286), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1278), .B1(new_n1293), .B2(new_n1255), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1293), .A2(new_n1255), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1265), .B(new_n1294), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1286), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1255), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1295), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1304), .A2(KEYINPUT62), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1264), .B1(new_n1298), .B2(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1294), .A2(new_n1265), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1304), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1296), .A2(KEYINPUT63), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1306), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(G375), .A2(new_n1251), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1299), .A2(new_n1314), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1315), .B(new_n1295), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1316), .B(new_n1308), .ZN(G402));
endmodule


