

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U552 ( .A(n690), .Z(n733) );
  XNOR2_X1 U553 ( .A(KEYINPUT71), .B(n589), .ZN(n950) );
  AND2_X1 U554 ( .A1(n763), .A2(n762), .ZN(n764) );
  OR2_X1 U555 ( .A1(n686), .A2(n685), .ZN(n689) );
  NOR2_X2 U556 ( .A1(G2104), .A2(n524), .ZN(n879) );
  XNOR2_X1 U557 ( .A(n703), .B(KEYINPUT29), .ZN(n704) );
  AND2_X2 U558 ( .A1(n524), .A2(G2104), .ZN(n874) );
  XNOR2_X1 U559 ( .A(n766), .B(KEYINPUT101), .ZN(n770) );
  NAND2_X1 U560 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U561 ( .A(n701), .B(KEYINPUT28), .Z(n518) );
  OR2_X1 U562 ( .A1(n769), .A2(n768), .ZN(n519) );
  NAND2_X2 U563 ( .A1(n573), .A2(n572), .ZN(n959) );
  NOR2_X2 U564 ( .A1(n558), .A2(n557), .ZN(G160) );
  XOR2_X1 U565 ( .A(KEYINPUT12), .B(n562), .Z(n520) );
  INV_X1 U566 ( .A(KEYINPUT27), .ZN(n692) );
  XNOR2_X1 U567 ( .A(n693), .B(n692), .ZN(n694) );
  INV_X1 U568 ( .A(KEYINPUT30), .ZN(n715) );
  XNOR2_X1 U569 ( .A(n715), .B(KEYINPUT97), .ZN(n716) );
  XNOR2_X1 U570 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U571 ( .A(n740), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U572 ( .A1(G160), .A2(G40), .ZN(n772) );
  INV_X1 U573 ( .A(KEYINPUT13), .ZN(n566) );
  XNOR2_X1 U574 ( .A(n566), .B(KEYINPUT69), .ZN(n567) );
  AND2_X1 U575 ( .A1(n770), .A2(n519), .ZN(n803) );
  XNOR2_X1 U576 ( .A(n568), .B(n567), .ZN(n569) );
  NOR2_X1 U577 ( .A1(G651), .A2(n649), .ZN(n643) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n636) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n537), .Z(n648) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n521), .Z(n873) );
  NAND2_X1 U582 ( .A1(G138), .A2(n873), .ZN(n523) );
  NAND2_X1 U583 ( .A1(G102), .A2(n874), .ZN(n522) );
  NAND2_X1 U584 ( .A1(n523), .A2(n522), .ZN(n528) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U586 ( .A1(G114), .A2(n878), .ZN(n526) );
  INV_X1 U587 ( .A(G2105), .ZN(n524) );
  NAND2_X1 U588 ( .A1(G126), .A2(n879), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n528), .A2(n527), .ZN(G164) );
  AND2_X1 U591 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U592 ( .A1(G135), .A2(n873), .ZN(n530) );
  NAND2_X1 U593 ( .A1(G111), .A2(n878), .ZN(n529) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n879), .A2(G123), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT18), .B(n531), .Z(n532) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n874), .A2(G99), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n1009) );
  XNOR2_X1 U600 ( .A(G2096), .B(n1009), .ZN(n536) );
  OR2_X1 U601 ( .A1(G2100), .A2(n536), .ZN(G156) );
  INV_X1 U602 ( .A(G651), .ZN(n540) );
  NOR2_X1 U603 ( .A1(G543), .A2(n540), .ZN(n537) );
  NAND2_X1 U604 ( .A1(G65), .A2(n648), .ZN(n539) );
  XOR2_X1 U605 ( .A(G543), .B(KEYINPUT0), .Z(n649) );
  NAND2_X1 U606 ( .A1(G53), .A2(n643), .ZN(n538) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n544) );
  NOR2_X1 U608 ( .A1(n649), .A2(n540), .ZN(n563) );
  NAND2_X1 U609 ( .A1(G78), .A2(n563), .ZN(n542) );
  NAND2_X1 U610 ( .A1(G91), .A2(n636), .ZN(n541) );
  NAND2_X1 U611 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n700) );
  INV_X1 U613 ( .A(n700), .ZN(G299) );
  INV_X1 U614 ( .A(G132), .ZN(G219) );
  INV_X1 U615 ( .A(G82), .ZN(G220) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  NAND2_X1 U617 ( .A1(G75), .A2(n563), .ZN(n546) );
  NAND2_X1 U618 ( .A1(G88), .A2(n636), .ZN(n545) );
  NAND2_X1 U619 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U620 ( .A1(G62), .A2(n648), .ZN(n548) );
  NAND2_X1 U621 ( .A1(G50), .A2(n643), .ZN(n547) );
  NAND2_X1 U622 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U623 ( .A1(n550), .A2(n549), .ZN(G166) );
  NAND2_X1 U624 ( .A1(G125), .A2(n879), .ZN(n551) );
  XNOR2_X1 U625 ( .A(n551), .B(KEYINPUT64), .ZN(n554) );
  NAND2_X1 U626 ( .A1(G101), .A2(n874), .ZN(n552) );
  XOR2_X1 U627 ( .A(KEYINPUT23), .B(n552), .Z(n553) );
  NAND2_X1 U628 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U629 ( .A1(G137), .A2(n873), .ZN(n556) );
  NAND2_X1 U630 ( .A1(G113), .A2(n878), .ZN(n555) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U632 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n822) );
  NAND2_X1 U634 ( .A1(n822), .A2(G567), .ZN(n560) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U636 ( .A1(n648), .A2(G56), .ZN(n561) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(n561), .Z(n570) );
  NAND2_X1 U638 ( .A1(n636), .A2(G81), .ZN(n562) );
  NAND2_X1 U639 ( .A1(n563), .A2(G68), .ZN(n564) );
  XOR2_X1 U640 ( .A(n564), .B(KEYINPUT68), .Z(n565) );
  NOR2_X1 U641 ( .A1(n520), .A2(n565), .ZN(n568) );
  NOR2_X1 U642 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U643 ( .A(n571), .B(KEYINPUT70), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G43), .A2(n643), .ZN(n572) );
  INV_X1 U645 ( .A(G860), .ZN(n608) );
  OR2_X1 U646 ( .A1(n959), .A2(n608), .ZN(G153) );
  NAND2_X1 U647 ( .A1(n563), .A2(G77), .ZN(n574) );
  XOR2_X1 U648 ( .A(KEYINPUT67), .B(n574), .Z(n576) );
  NAND2_X1 U649 ( .A1(n636), .A2(G90), .ZN(n575) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U651 ( .A(KEYINPUT9), .B(n577), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G64), .A2(n648), .ZN(n579) );
  NAND2_X1 U653 ( .A1(G52), .A2(n643), .ZN(n578) );
  AND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G79), .A2(n563), .ZN(n583) );
  NAND2_X1 U657 ( .A1(G66), .A2(n648), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G92), .A2(n636), .ZN(n585) );
  NAND2_X1 U660 ( .A1(G54), .A2(n643), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n588), .Z(n589) );
  INV_X1 U664 ( .A(G868), .ZN(n661) );
  NAND2_X1 U665 ( .A1(n950), .A2(n661), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n590), .B(KEYINPUT72), .ZN(n592) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U669 ( .A1(n636), .A2(G89), .ZN(n593) );
  XNOR2_X1 U670 ( .A(n593), .B(KEYINPUT4), .ZN(n595) );
  NAND2_X1 U671 ( .A1(G76), .A2(n563), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U673 ( .A(KEYINPUT5), .B(n596), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n643), .A2(G51), .ZN(n597) );
  XOR2_X1 U675 ( .A(KEYINPUT73), .B(n597), .Z(n599) );
  NAND2_X1 U676 ( .A1(n648), .A2(G63), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U678 ( .A(KEYINPUT6), .B(n600), .Z(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U680 ( .A(KEYINPUT7), .B(n603), .ZN(G168) );
  XOR2_X1 U681 ( .A(G168), .B(KEYINPUT8), .Z(n604) );
  XNOR2_X1 U682 ( .A(KEYINPUT74), .B(n604), .ZN(G286) );
  XNOR2_X1 U683 ( .A(KEYINPUT75), .B(G868), .ZN(n605) );
  NOR2_X1 U684 ( .A1(G286), .A2(n605), .ZN(n607) );
  NOR2_X1 U685 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U686 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n608), .A2(G559), .ZN(n609) );
  INV_X1 U688 ( .A(n950), .ZN(n894) );
  NAND2_X1 U689 ( .A1(n609), .A2(n894), .ZN(n610) );
  XNOR2_X1 U690 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U691 ( .A1(n950), .A2(n661), .ZN(n611) );
  XOR2_X1 U692 ( .A(KEYINPUT76), .B(n611), .Z(n612) );
  NOR2_X1 U693 ( .A1(G559), .A2(n612), .ZN(n614) );
  NOR2_X1 U694 ( .A1(G868), .A2(n959), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U696 ( .A1(G559), .A2(n894), .ZN(n615) );
  XNOR2_X1 U697 ( .A(n615), .B(n959), .ZN(n658) );
  NOR2_X1 U698 ( .A1(G860), .A2(n658), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G80), .A2(n563), .ZN(n617) );
  NAND2_X1 U700 ( .A1(G93), .A2(n636), .ZN(n616) );
  NAND2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G67), .A2(n648), .ZN(n619) );
  NAND2_X1 U703 ( .A1(G55), .A2(n643), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U705 ( .A(KEYINPUT77), .B(n620), .Z(n621) );
  OR2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n662) );
  XOR2_X1 U707 ( .A(n662), .B(KEYINPUT78), .Z(n623) );
  XNOR2_X1 U708 ( .A(n624), .B(n623), .ZN(G145) );
  NAND2_X1 U709 ( .A1(G73), .A2(n563), .ZN(n625) );
  XNOR2_X1 U710 ( .A(n625), .B(KEYINPUT2), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G86), .A2(n636), .ZN(n627) );
  NAND2_X1 U712 ( .A1(G48), .A2(n643), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U714 ( .A1(G61), .A2(n648), .ZN(n628) );
  XNOR2_X1 U715 ( .A(KEYINPUT81), .B(n628), .ZN(n629) );
  NOR2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U718 ( .A1(n563), .A2(G72), .ZN(n633) );
  XNOR2_X1 U719 ( .A(KEYINPUT66), .B(n633), .ZN(n641) );
  NAND2_X1 U720 ( .A1(G60), .A2(n648), .ZN(n635) );
  NAND2_X1 U721 ( .A1(G47), .A2(n643), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U723 ( .A1(G85), .A2(n636), .ZN(n637) );
  XNOR2_X1 U724 ( .A(KEYINPUT65), .B(n637), .ZN(n638) );
  NOR2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U727 ( .A1(G651), .A2(G74), .ZN(n642) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n642), .Z(n645) );
  NAND2_X1 U729 ( .A1(n643), .A2(G49), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U731 ( .A(KEYINPUT80), .B(n646), .ZN(n647) );
  NOR2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n649), .A2(G87), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(G288) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n653) );
  XNOR2_X1 U736 ( .A(G305), .B(n700), .ZN(n652) );
  XNOR2_X1 U737 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U738 ( .A(n662), .B(n654), .Z(n656) );
  XNOR2_X1 U739 ( .A(G290), .B(G166), .ZN(n655) );
  XNOR2_X1 U740 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U741 ( .A(n657), .B(G288), .ZN(n893) );
  XNOR2_X1 U742 ( .A(n893), .B(n658), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n659), .A2(G868), .ZN(n660) );
  XOR2_X1 U744 ( .A(KEYINPUT83), .B(n660), .Z(n664) );
  NAND2_X1 U745 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U751 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U753 ( .A1(G69), .A2(G120), .ZN(n669) );
  NOR2_X1 U754 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U755 ( .A1(G108), .A2(n670), .ZN(n827) );
  NAND2_X1 U756 ( .A1(n827), .A2(G567), .ZN(n676) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U759 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G96), .A2(n673), .ZN(n826) );
  NAND2_X1 U761 ( .A1(G2106), .A2(n826), .ZN(n674) );
  XNOR2_X1 U762 ( .A(KEYINPUT84), .B(n674), .ZN(n675) );
  NAND2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n849) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U765 ( .A1(n849), .A2(n677), .ZN(n825) );
  NAND2_X1 U766 ( .A1(n825), .A2(G36), .ZN(G176) );
  INV_X1 U767 ( .A(G166), .ZN(G303) );
  INV_X1 U768 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U769 ( .A(KEYINPUT89), .B(n772), .ZN(n678) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NAND2_X1 U771 ( .A1(n678), .A2(n771), .ZN(n690) );
  NAND2_X1 U772 ( .A1(G8), .A2(n733), .ZN(n769) );
  NOR2_X1 U773 ( .A1(G1966), .A2(n769), .ZN(n713) );
  INV_X1 U774 ( .A(n713), .ZN(n726) );
  INV_X1 U775 ( .A(G1996), .ZN(n847) );
  NOR2_X1 U776 ( .A1(n733), .A2(n847), .ZN(n679) );
  XOR2_X1 U777 ( .A(n679), .B(KEYINPUT26), .Z(n681) );
  NAND2_X1 U778 ( .A1(n733), .A2(G1341), .ZN(n680) );
  NAND2_X1 U779 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U780 ( .A1(n959), .A2(n682), .ZN(n686) );
  NAND2_X1 U781 ( .A1(G1348), .A2(n733), .ZN(n684) );
  NAND2_X1 U782 ( .A1(G2067), .A2(n691), .ZN(n683) );
  NAND2_X1 U783 ( .A1(n684), .A2(n683), .ZN(n687) );
  NOR2_X1 U784 ( .A1(n950), .A2(n687), .ZN(n685) );
  NAND2_X1 U785 ( .A1(n950), .A2(n687), .ZN(n688) );
  NAND2_X1 U786 ( .A1(n689), .A2(n688), .ZN(n698) );
  XNOR2_X1 U787 ( .A(G1956), .B(KEYINPUT92), .ZN(n980) );
  NAND2_X1 U788 ( .A1(n733), .A2(n980), .ZN(n695) );
  INV_X1 U789 ( .A(n690), .ZN(n691) );
  NAND2_X1 U790 ( .A1(n691), .A2(G2072), .ZN(n693) );
  NAND2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U792 ( .A(n696), .B(KEYINPUT93), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n518), .ZN(n705) );
  XNOR2_X1 U797 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n703) );
  XNOR2_X1 U798 ( .A(n705), .B(n704), .ZN(n711) );
  XOR2_X1 U799 ( .A(G2078), .B(KEYINPUT90), .Z(n706) );
  XNOR2_X1 U800 ( .A(KEYINPUT25), .B(n706), .ZN(n923) );
  NAND2_X1 U801 ( .A1(n923), .A2(n691), .ZN(n708) );
  NAND2_X1 U802 ( .A1(G1961), .A2(n733), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U804 ( .A(n709), .B(KEYINPUT91), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n719), .A2(G171), .ZN(n710) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U807 ( .A(n712), .B(KEYINPUT96), .ZN(n724) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n733), .ZN(n728) );
  NOR2_X1 U809 ( .A1(n728), .A2(n713), .ZN(n714) );
  NAND2_X1 U810 ( .A1(G8), .A2(n714), .ZN(n717) );
  NOR2_X1 U811 ( .A1(G168), .A2(n718), .ZN(n721) );
  NOR2_X1 U812 ( .A1(G171), .A2(n719), .ZN(n720) );
  NOR2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U814 ( .A(KEYINPUT31), .B(n722), .Z(n723) );
  NAND2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U816 ( .A(n725), .B(KEYINPUT98), .ZN(n731) );
  AND2_X1 U817 ( .A1(n726), .A2(n731), .ZN(n727) );
  XOR2_X1 U818 ( .A(KEYINPUT99), .B(n727), .Z(n730) );
  NAND2_X1 U819 ( .A1(G8), .A2(n728), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n755) );
  NAND2_X1 U821 ( .A1(n731), .A2(G286), .ZN(n738) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n769), .ZN(n732) );
  XNOR2_X1 U823 ( .A(n732), .B(KEYINPUT100), .ZN(n735) );
  NOR2_X1 U824 ( .A1(n733), .A2(G2090), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n736), .A2(G303), .ZN(n737) );
  NAND2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n739), .A2(G8), .ZN(n740) );
  AND2_X1 U829 ( .A1(n753), .A2(n769), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n755), .A2(n741), .ZN(n745) );
  NOR2_X1 U831 ( .A1(G2090), .A2(G303), .ZN(n742) );
  NAND2_X1 U832 ( .A1(G8), .A2(n742), .ZN(n743) );
  OR2_X1 U833 ( .A1(n746), .A2(n743), .ZN(n744) );
  AND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n765) );
  INV_X1 U835 ( .A(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n946) );
  INV_X1 U837 ( .A(n769), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n946), .A2(n746), .ZN(n747) );
  AND2_X1 U839 ( .A1(n758), .A2(n747), .ZN(n752) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n944) );
  NAND2_X1 U841 ( .A1(n944), .A2(KEYINPUT33), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n748), .A2(n769), .ZN(n750) );
  XOR2_X1 U843 ( .A(G1981), .B(G305), .Z(n941) );
  INV_X1 U844 ( .A(n941), .ZN(n749) );
  OR2_X1 U845 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U846 ( .A1(n752), .A2(n751), .ZN(n756) );
  AND2_X1 U847 ( .A1(n753), .A2(n756), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n763) );
  INV_X1 U849 ( .A(n756), .ZN(n761) );
  NOR2_X1 U850 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U851 ( .A1(n944), .A2(n757), .ZN(n759) );
  AND2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n760) );
  OR2_X1 U853 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U856 ( .A(n767), .B(KEYINPUT24), .Z(n768) );
  NOR2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U858 ( .A(n773), .B(KEYINPUT86), .Z(n800) );
  INV_X1 U859 ( .A(n800), .ZN(n817) );
  NAND2_X1 U860 ( .A1(G140), .A2(n873), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G104), .A2(n874), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n777) );
  XOR2_X1 U863 ( .A(KEYINPUT34), .B(KEYINPUT87), .Z(n776) );
  XNOR2_X1 U864 ( .A(n777), .B(n776), .ZN(n782) );
  NAND2_X1 U865 ( .A1(G116), .A2(n878), .ZN(n779) );
  NAND2_X1 U866 ( .A1(G128), .A2(n879), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U868 ( .A(KEYINPUT35), .B(n780), .Z(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U870 ( .A(KEYINPUT36), .B(n783), .ZN(n890) );
  XNOR2_X1 U871 ( .A(G2067), .B(KEYINPUT37), .ZN(n807) );
  NOR2_X1 U872 ( .A1(n890), .A2(n807), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n784), .B(KEYINPUT88), .ZN(n1011) );
  NAND2_X1 U874 ( .A1(n817), .A2(n1011), .ZN(n814) );
  NAND2_X1 U875 ( .A1(G131), .A2(n873), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G107), .A2(n878), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U878 ( .A1(G95), .A2(n874), .ZN(n788) );
  NAND2_X1 U879 ( .A1(G119), .A2(n879), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  OR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n885) );
  AND2_X1 U882 ( .A1(n885), .A2(G1991), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G141), .A2(n873), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G117), .A2(n878), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n874), .A2(G105), .ZN(n793) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n793), .Z(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n879), .A2(G129), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n857) );
  AND2_X1 U891 ( .A1(G1996), .A2(n857), .ZN(n798) );
  NOR2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n1006) );
  NOR2_X1 U893 ( .A1(n800), .A2(n1006), .ZN(n811) );
  INV_X1 U894 ( .A(n811), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n814), .A2(n801), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n806) );
  XOR2_X1 U897 ( .A(G1986), .B(KEYINPUT85), .Z(n804) );
  XNOR2_X1 U898 ( .A(G290), .B(n804), .ZN(n956) );
  NAND2_X1 U899 ( .A1(n956), .A2(n817), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n820) );
  NAND2_X1 U901 ( .A1(n890), .A2(n807), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n808), .B(KEYINPUT102), .ZN(n1015) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n857), .ZN(n1003) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n885), .ZN(n1008) );
  NOR2_X1 U906 ( .A1(n809), .A2(n1008), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n1003), .A2(n812), .ZN(n813) );
  XNOR2_X1 U909 ( .A(n813), .B(KEYINPUT39), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n1015), .A2(n816), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U914 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U917 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XOR2_X1 U926 ( .A(G2678), .B(KEYINPUT43), .Z(n829) );
  XNOR2_X1 U927 ( .A(KEYINPUT106), .B(KEYINPUT105), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U929 ( .A(KEYINPUT42), .B(G2072), .Z(n831) );
  XNOR2_X1 U930 ( .A(G2067), .B(G2090), .ZN(n830) );
  XNOR2_X1 U931 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U932 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U933 ( .A(G2096), .B(G2100), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n837) );
  XOR2_X1 U935 ( .A(G2084), .B(G2078), .Z(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U937 ( .A(G1971), .B(G1981), .Z(n839) );
  XNOR2_X1 U938 ( .A(G1991), .B(G1986), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(G1976), .B(G1956), .Z(n841) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1961), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U944 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U946 ( .A(G2474), .B(n846), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(G229) );
  INV_X1 U948 ( .A(n849), .ZN(G319) );
  NAND2_X1 U949 ( .A1(G124), .A2(n879), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n878), .A2(G112), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G136), .A2(n873), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G100), .A2(n874), .ZN(n853) );
  NAND2_X1 U955 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U956 ( .A1(n856), .A2(n855), .ZN(G162) );
  XNOR2_X1 U957 ( .A(G160), .B(n857), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n858), .B(n1009), .ZN(n859) );
  XNOR2_X1 U959 ( .A(G164), .B(n859), .ZN(n889) );
  XOR2_X1 U960 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n861) );
  XNOR2_X1 U961 ( .A(G162), .B(KEYINPUT48), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n872) );
  NAND2_X1 U963 ( .A1(G118), .A2(n878), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G130), .A2(n879), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n870) );
  NAND2_X1 U966 ( .A1(n874), .A2(G106), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n864), .B(KEYINPUT108), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G142), .A2(n873), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(KEYINPUT109), .B(n867), .ZN(n868) );
  XNOR2_X1 U971 ( .A(KEYINPUT45), .B(n868), .ZN(n869) );
  NOR2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(n872), .B(n871), .Z(n887) );
  NAND2_X1 U974 ( .A1(G139), .A2(n873), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G103), .A2(n874), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(KEYINPUT110), .B(n877), .ZN(n884) );
  NAND2_X1 U978 ( .A1(G115), .A2(n878), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G127), .A2(n879), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n998) );
  XOR2_X1 U983 ( .A(n885), .B(n998), .Z(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U986 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U987 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U988 ( .A(G286), .B(n893), .ZN(n896) );
  XNOR2_X1 U989 ( .A(G171), .B(n894), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U991 ( .A(n897), .B(n959), .Z(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G397) );
  NOR2_X1 U993 ( .A1(G227), .A2(G229), .ZN(n900) );
  XNOR2_X1 U994 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n913) );
  XNOR2_X1 U996 ( .A(G2451), .B(G2435), .ZN(n910) );
  XOR2_X1 U997 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n902) );
  XNOR2_X1 U998 ( .A(G2454), .B(G2430), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1000 ( .A(G2446), .B(G2438), .Z(n904) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1003 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G2443), .B(G2427), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n911), .A2(G14), .ZN(n916) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n916), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n916), .ZN(G401) );
  XNOR2_X1 U1015 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1029) );
  XOR2_X1 U1016 ( .A(G29), .B(KEYINPUT120), .Z(n939) );
  XOR2_X1 U1017 ( .A(KEYINPUT119), .B(G34), .Z(n918) );
  XNOR2_X1 U1018 ( .A(G2084), .B(KEYINPUT54), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(n918), .B(n917), .ZN(n936) );
  XOR2_X1 U1020 ( .A(G2090), .B(G35), .Z(n934) );
  XOR2_X1 U1021 ( .A(G25), .B(G1991), .Z(n919) );
  NAND2_X1 U1022 ( .A1(n919), .A2(G28), .ZN(n929) );
  XNOR2_X1 U1023 ( .A(G2067), .B(G26), .ZN(n921) );
  XNOR2_X1 U1024 ( .A(G2072), .B(G33), .ZN(n920) );
  NOR2_X1 U1025 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1026 ( .A(KEYINPUT116), .B(n922), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(n923), .B(G27), .ZN(n925) );
  XNOR2_X1 U1028 ( .A(G32), .B(G1996), .ZN(n924) );
  NOR2_X1 U1029 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(n931), .B(n930), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(n932), .B(KEYINPUT53), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(KEYINPUT55), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(G11), .A2(n940), .ZN(n996) );
  XNOR2_X1 U1040 ( .A(G16), .B(KEYINPUT56), .ZN(n965) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G168), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT57), .ZN(n963) );
  INV_X1 U1044 ( .A(n944), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1046 ( .A(KEYINPUT121), .B(n947), .Z(n949) );
  XNOR2_X1 U1047 ( .A(G1961), .B(G301), .ZN(n948) );
  NOR2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G166), .B(G1971), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n950), .B(G1348), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(G299), .B(G1956), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G1341), .B(n959), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n994) );
  INV_X1 U1060 ( .A(G16), .ZN(n992) );
  XOR2_X1 U1061 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n972) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G22), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(G23), .B(G1976), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n970) );
  XOR2_X1 U1065 ( .A(G1986), .B(KEYINPUT124), .Z(n968) );
  XNOR2_X1 U1066 ( .A(G24), .B(n968), .ZN(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(n972), .B(n971), .ZN(n989) );
  XNOR2_X1 U1069 ( .A(G1981), .B(G6), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(KEYINPUT122), .B(n975), .ZN(n979) );
  XOR2_X1 U1073 ( .A(G4), .B(KEYINPUT123), .Z(n977) );
  XNOR2_X1 U1074 ( .A(G1348), .B(KEYINPUT59), .ZN(n976) );
  XNOR2_X1 U1075 ( .A(n977), .B(n976), .ZN(n978) );
  NAND2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(G20), .B(n980), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(KEYINPUT60), .B(n983), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G21), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(G5), .B(G1961), .ZN(n984) );
  NOR2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(KEYINPUT61), .B(n990), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(KEYINPUT126), .ZN(n1027) );
  XNOR2_X1 U1090 ( .A(KEYINPUT52), .B(KEYINPUT114), .ZN(n1022) );
  XOR2_X1 U1091 ( .A(G2072), .B(n998), .Z(n1000) );
  XOR2_X1 U1092 ( .A(G164), .B(G2078), .Z(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(KEYINPUT50), .B(n1001), .ZN(n1019) );
  XOR2_X1 U1095 ( .A(G2090), .B(G162), .Z(n1002) );
  NOR2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1097 ( .A(KEYINPUT51), .B(n1004), .Z(n1005) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1017) );
  XOR2_X1 U1099 ( .A(G160), .B(G2084), .Z(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1103 ( .A(KEYINPUT113), .B(n1013), .Z(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(n1020), .B(KEYINPUT115), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1022), .B(n1021), .ZN(n1024) );
  INV_X1 U1109 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(n1029), .B(n1028), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

