

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772;

  XOR2_X1 U375 ( .A(G122), .B(G104), .Z(n447) );
  XNOR2_X1 U376 ( .A(G101), .B(G146), .ZN(n483) );
  BUF_X1 U377 ( .A(G143), .Z(n353) );
  BUF_X1 U378 ( .A(G113), .Z(n675) );
  NAND2_X1 U379 ( .A1(n352), .A2(n374), .ZN(n402) );
  XNOR2_X2 U380 ( .A(n405), .B(n404), .ZN(n352) );
  XNOR2_X2 U381 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X2 U382 ( .A(n647), .B(KEYINPUT62), .ZN(n648) );
  XNOR2_X2 U383 ( .A(n436), .B(KEYINPUT0), .ZN(n437) );
  XNOR2_X2 U384 ( .A(KEYINPUT15), .B(G902), .ZN(n635) );
  AND2_X2 U385 ( .A1(n653), .A2(KEYINPUT44), .ZN(n557) );
  XNOR2_X2 U386 ( .A(n480), .B(n479), .ZN(n497) );
  XNOR2_X2 U387 ( .A(n497), .B(n500), .ZN(n757) );
  XNOR2_X1 U388 ( .A(G134), .B(G116), .ZN(n455) );
  NOR2_X2 U389 ( .A1(n684), .A2(n642), .ZN(n730) );
  NOR2_X2 U390 ( .A1(n684), .A2(n642), .ZN(n385) );
  XNOR2_X2 U391 ( .A(n440), .B(KEYINPUT10), .ZN(n756) );
  AND2_X2 U392 ( .A1(n398), .A2(n397), .ZN(n396) );
  XNOR2_X2 U393 ( .A(n438), .B(n437), .ZN(n542) );
  XNOR2_X2 U394 ( .A(n399), .B(G128), .ZN(n465) );
  XNOR2_X2 U395 ( .A(KEYINPUT65), .B(G143), .ZN(n399) );
  XNOR2_X2 U396 ( .A(G116), .B(G113), .ZN(n412) );
  INV_X1 U397 ( .A(n538), .ZN(n551) );
  INV_X2 U398 ( .A(G953), .ZN(n765) );
  OR2_X1 U399 ( .A1(n515), .A2(n689), .ZN(n516) );
  OR2_X1 U400 ( .A1(n647), .A2(G902), .ZN(n498) );
  INV_X1 U401 ( .A(G146), .ZN(n418) );
  NOR2_X1 U402 ( .A1(G953), .A2(n721), .ZN(n723) );
  OR2_X1 U403 ( .A1(n685), .A2(n686), .ZN(n373) );
  AND2_X1 U404 ( .A1(n550), .A2(n559), .ZN(n366) );
  XNOR2_X1 U405 ( .A(n695), .B(KEYINPUT6), .ZN(n550) );
  OR2_X1 U406 ( .A1(n556), .A2(n555), .ZN(n706) );
  NOR2_X1 U407 ( .A1(n726), .A2(G902), .ZN(n365) );
  XNOR2_X1 U408 ( .A(n757), .B(n487), .ZN(n726) );
  XNOR2_X1 U409 ( .A(n421), .B(n420), .ZN(n391) );
  XNOR2_X1 U410 ( .A(n465), .B(n375), .ZN(n480) );
  XNOR2_X1 U411 ( .A(n418), .B(G125), .ZN(n439) );
  XOR2_X1 U412 ( .A(KEYINPUT23), .B(G110), .Z(n502) );
  XNOR2_X2 U413 ( .A(G110), .B(G104), .ZN(n416) );
  BUF_X2 U414 ( .A(n537), .Z(n477) );
  XNOR2_X1 U415 ( .A(n354), .B(KEYINPUT32), .ZN(n654) );
  NAND2_X1 U416 ( .A1(n654), .A2(n560), .ZN(n407) );
  NAND2_X1 U417 ( .A1(n537), .A2(n366), .ZN(n354) );
  XNOR2_X2 U418 ( .A(n476), .B(n475), .ZN(n537) );
  NAND2_X1 U419 ( .A1(n355), .A2(n369), .ZN(n392) );
  XNOR2_X1 U420 ( .A(n356), .B(n563), .ZN(n355) );
  NAND2_X1 U421 ( .A1(n358), .A2(n357), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n562), .B(KEYINPUT66), .ZN(n357) );
  NOR2_X1 U423 ( .A1(n558), .A2(n557), .ZN(n358) );
  INV_X1 U424 ( .A(n565), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n402), .B(KEYINPUT35), .ZN(n653) );
  AND2_X1 U426 ( .A1(n538), .A2(n550), .ZN(n360) );
  OR2_X2 U427 ( .A1(n741), .A2(n391), .ZN(n362) );
  NAND2_X1 U428 ( .A1(n741), .A2(n391), .ZN(n361) );
  NAND2_X1 U429 ( .A1(n362), .A2(n361), .ZN(n390) );
  BUF_X1 U430 ( .A(n548), .Z(n363) );
  NAND2_X1 U431 ( .A1(n400), .A2(n573), .ZN(n548) );
  XNOR2_X1 U432 ( .A(n540), .B(n383), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n540), .B(n383), .ZN(n554) );
  XNOR2_X2 U434 ( .A(n365), .B(G469), .ZN(n580) );
  BUF_X2 U435 ( .A(n542), .Z(n540) );
  XNOR2_X2 U436 ( .A(n580), .B(KEYINPUT1), .ZN(n538) );
  NAND2_X1 U437 ( .A1(n396), .A2(n394), .ZN(n367) );
  NAND2_X1 U438 ( .A1(n396), .A2(n394), .ZN(n595) );
  INV_X1 U439 ( .A(n604), .ZN(n368) );
  XNOR2_X1 U440 ( .A(KEYINPUT3), .B(G119), .ZN(n413) );
  XNOR2_X1 U441 ( .A(KEYINPUT71), .B(G131), .ZN(n478) );
  INV_X1 U442 ( .A(KEYINPUT72), .ZN(n481) );
  NOR2_X1 U443 ( .A1(n569), .A2(KEYINPUT19), .ZN(n395) );
  XNOR2_X1 U444 ( .A(G128), .B(G119), .ZN(n501) );
  XNOR2_X1 U445 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n461) );
  INV_X1 U446 ( .A(KEYINPUT93), .ZN(n383) );
  AND2_X1 U447 ( .A1(n646), .A2(G953), .ZN(n740) );
  NAND2_X1 U448 ( .A1(n385), .A2(G210), .ZN(n382) );
  INV_X1 U449 ( .A(KEYINPUT89), .ZN(n406) );
  XNOR2_X1 U450 ( .A(n439), .B(n419), .ZN(n420) );
  XNOR2_X1 U451 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n419) );
  NAND2_X1 U452 ( .A1(G234), .A2(G237), .ZN(n429) );
  XNOR2_X1 U453 ( .A(G146), .B(G137), .ZN(n490) );
  XOR2_X1 U454 ( .A(KEYINPUT77), .B(KEYINPUT5), .Z(n491) );
  NOR2_X1 U455 ( .A1(G953), .A2(G237), .ZN(n492) );
  OR2_X1 U456 ( .A1(n576), .A2(n569), .ZN(n526) );
  NAND2_X1 U457 ( .A1(n595), .A2(n435), .ZN(n438) );
  XNOR2_X1 U458 ( .A(KEYINPUT16), .B(G122), .ZN(n415) );
  XOR2_X1 U459 ( .A(G122), .B(G107), .Z(n456) );
  XNOR2_X1 U460 ( .A(KEYINPUT100), .B(KEYINPUT9), .ZN(n457) );
  XOR2_X1 U461 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n458) );
  INV_X1 U462 ( .A(KEYINPUT34), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n508), .B(n507), .ZN(n736) );
  NAND2_X1 U464 ( .A1(n477), .A2(n370), .ZN(n560) );
  AND2_X2 U465 ( .A1(n364), .A2(n544), .ZN(n666) );
  XNOR2_X1 U466 ( .A(n401), .B(KEYINPUT87), .ZN(n400) );
  INV_X1 U467 ( .A(n740), .ZN(n380) );
  NAND2_X1 U468 ( .A1(n376), .A2(n566), .ZN(n369) );
  NOR2_X1 U469 ( .A1(n551), .A2(n514), .ZN(n370) );
  XOR2_X1 U470 ( .A(n644), .B(n645), .Z(n371) );
  XOR2_X1 U471 ( .A(n720), .B(KEYINPUT115), .Z(n372) );
  XOR2_X1 U472 ( .A(n605), .B(KEYINPUT79), .Z(n374) );
  XOR2_X1 U473 ( .A(KEYINPUT70), .B(KEYINPUT4), .Z(n375) );
  XOR2_X1 U474 ( .A(n384), .B(n406), .Z(n376) );
  NOR2_X1 U475 ( .A1(n717), .A2(n372), .ZN(n377) );
  XNOR2_X1 U476 ( .A(KEYINPUT117), .B(KEYINPUT56), .ZN(n378) );
  XNOR2_X1 U477 ( .A(n379), .B(n378), .ZN(G51) );
  NAND2_X1 U478 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U479 ( .A(n382), .B(n371), .ZN(n381) );
  NOR2_X1 U480 ( .A1(n678), .A2(n666), .ZN(n545) );
  BUF_X1 U481 ( .A(n407), .Z(n384) );
  XNOR2_X1 U482 ( .A(n407), .B(n406), .ZN(n561) );
  NOR2_X2 U483 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U484 ( .A(n392), .B(n567), .ZN(n746) );
  NAND2_X1 U485 ( .A1(n386), .A2(n704), .ZN(n532) );
  INV_X1 U486 ( .A(n607), .ZN(n386) );
  NAND2_X1 U487 ( .A1(n388), .A2(n387), .ZN(n587) );
  INV_X1 U488 ( .A(n770), .ZN(n387) );
  INV_X1 U489 ( .A(n585), .ZN(n388) );
  XNOR2_X2 U490 ( .A(n536), .B(n535), .ZN(n585) );
  XNOR2_X1 U491 ( .A(n549), .B(KEYINPUT102), .ZN(n558) );
  NAND2_X1 U492 ( .A1(n643), .A2(n635), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n390), .B(n389), .ZN(n643) );
  XNOR2_X1 U494 ( .A(n422), .B(n486), .ZN(n389) );
  XNOR2_X1 U495 ( .A(n488), .B(n415), .ZN(n741) );
  NAND2_X1 U496 ( .A1(n393), .A2(n395), .ZN(n394) );
  INV_X1 U497 ( .A(n529), .ZN(n393) );
  XNOR2_X2 U498 ( .A(n426), .B(n425), .ZN(n529) );
  NAND2_X1 U499 ( .A1(n569), .A2(KEYINPUT19), .ZN(n397) );
  NAND2_X1 U500 ( .A1(n529), .A2(KEYINPUT19), .ZN(n398) );
  INV_X1 U501 ( .A(n363), .ZN(n663) );
  NAND2_X1 U502 ( .A1(n360), .A2(n477), .ZN(n401) );
  NAND2_X1 U503 ( .A1(n709), .A2(n554), .ZN(n405) );
  NAND2_X1 U504 ( .A1(n408), .A2(n377), .ZN(n721) );
  NAND2_X1 U505 ( .A1(n373), .A2(n409), .ZN(n408) );
  INV_X1 U506 ( .A(n684), .ZN(n409) );
  BUF_X1 U507 ( .A(n385), .Z(n734) );
  BUF_X1 U508 ( .A(n741), .Z(n743) );
  AND2_X1 U509 ( .A1(G214), .A2(n492), .ZN(n410) );
  INV_X1 U510 ( .A(n546), .ZN(n547) );
  NAND2_X1 U511 ( .A1(n548), .A2(n547), .ZN(n549) );
  INV_X1 U512 ( .A(KEYINPUT88), .ZN(n563) );
  XNOR2_X1 U513 ( .A(n439), .B(G140), .ZN(n440) );
  XNOR2_X1 U514 ( .A(KEYINPUT74), .B(KEYINPUT24), .ZN(n499) );
  XNOR2_X1 U515 ( .A(n443), .B(n410), .ZN(n444) );
  XNOR2_X1 U516 ( .A(n500), .B(n499), .ZN(n504) );
  XNOR2_X1 U517 ( .A(n756), .B(n444), .ZN(n450) );
  AND2_X1 U518 ( .A1(n625), .A2(n624), .ZN(n759) );
  NOR2_X1 U519 ( .A1(n539), .A2(n538), .ZN(n697) );
  XNOR2_X1 U520 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U521 ( .A(n541), .B(KEYINPUT31), .ZN(n678) );
  XNOR2_X1 U522 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X2 U523 ( .A(G101), .B(KEYINPUT73), .ZN(n411) );
  XNOR2_X1 U524 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U525 ( .A(n414), .B(n413), .ZN(n488) );
  XNOR2_X1 U526 ( .A(n416), .B(G107), .ZN(n742) );
  XNOR2_X1 U527 ( .A(n742), .B(KEYINPUT75), .ZN(n486) );
  NAND2_X1 U528 ( .A1(n765), .A2(G224), .ZN(n417) );
  XNOR2_X1 U529 ( .A(n417), .B(KEYINPUT91), .ZN(n421) );
  INV_X1 U530 ( .A(n480), .ZN(n422) );
  NOR2_X1 U531 ( .A1(G237), .A2(G902), .ZN(n423) );
  XNOR2_X1 U532 ( .A(n423), .B(KEYINPUT76), .ZN(n427) );
  INV_X1 U533 ( .A(G210), .ZN(n424) );
  OR2_X1 U534 ( .A1(n427), .A2(n424), .ZN(n425) );
  INV_X1 U535 ( .A(n427), .ZN(n428) );
  AND2_X1 U536 ( .A1(n428), .A2(G214), .ZN(n569) );
  XNOR2_X1 U537 ( .A(n429), .B(KEYINPUT14), .ZN(n432) );
  NAND2_X1 U538 ( .A1(G952), .A2(n432), .ZN(n430) );
  XNOR2_X1 U539 ( .A(KEYINPUT92), .B(n430), .ZN(n715) );
  INV_X1 U540 ( .A(n715), .ZN(n431) );
  NAND2_X1 U541 ( .A1(n431), .A2(n765), .ZN(n522) );
  NAND2_X1 U542 ( .A1(G902), .A2(n432), .ZN(n518) );
  INV_X1 U543 ( .A(n518), .ZN(n433) );
  NOR2_X1 U544 ( .A1(G898), .A2(n765), .ZN(n744) );
  NAND2_X1 U545 ( .A1(n433), .A2(n744), .ZN(n434) );
  NAND2_X1 U546 ( .A1(n522), .A2(n434), .ZN(n435) );
  INV_X1 U547 ( .A(KEYINPUT68), .ZN(n436) );
  XOR2_X1 U548 ( .A(KEYINPUT95), .B(KEYINPUT12), .Z(n442) );
  XNOR2_X1 U549 ( .A(KEYINPUT11), .B(KEYINPUT94), .ZN(n441) );
  XNOR2_X1 U550 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U551 ( .A(n353), .B(n675), .ZN(n445) );
  XNOR2_X1 U552 ( .A(KEYINPUT96), .B(n445), .ZN(n446) );
  XNOR2_X1 U553 ( .A(n478), .B(n446), .ZN(n448) );
  XNOR2_X1 U554 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U555 ( .A(n450), .B(n449), .ZN(n658) );
  INV_X1 U556 ( .A(G902), .ZN(n467) );
  NAND2_X1 U557 ( .A1(n658), .A2(n467), .ZN(n454) );
  XOR2_X1 U558 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n452) );
  XNOR2_X1 U559 ( .A(KEYINPUT13), .B(G475), .ZN(n451) );
  XOR2_X1 U560 ( .A(n452), .B(n451), .Z(n453) );
  XNOR2_X1 U561 ( .A(n454), .B(n453), .ZN(n556) );
  XNOR2_X1 U562 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U563 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U564 ( .A(n460), .B(n459), .Z(n464) );
  NAND2_X1 U565 ( .A1(n765), .A2(G234), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n462), .B(n461), .ZN(n505) );
  NAND2_X1 U567 ( .A1(G217), .A2(n505), .ZN(n463) );
  XNOR2_X1 U568 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U569 ( .A(n466), .B(n465), .ZN(n732) );
  NAND2_X1 U570 ( .A1(n732), .A2(n467), .ZN(n470) );
  INV_X1 U571 ( .A(KEYINPUT101), .ZN(n468) );
  XNOR2_X1 U572 ( .A(n468), .B(G478), .ZN(n469) );
  XNOR2_X1 U573 ( .A(n470), .B(n469), .ZN(n555) );
  NAND2_X1 U574 ( .A1(G234), .A2(n635), .ZN(n471) );
  XNOR2_X1 U575 ( .A(KEYINPUT20), .B(n471), .ZN(n509) );
  NAND2_X1 U576 ( .A1(n509), .A2(G221), .ZN(n473) );
  INV_X1 U577 ( .A(KEYINPUT21), .ZN(n472) );
  XNOR2_X1 U578 ( .A(n473), .B(n472), .ZN(n574) );
  INV_X1 U579 ( .A(n574), .ZN(n689) );
  NOR2_X1 U580 ( .A1(n706), .A2(n689), .ZN(n474) );
  NAND2_X1 U581 ( .A1(n542), .A2(n474), .ZN(n476) );
  INV_X1 U582 ( .A(KEYINPUT22), .ZN(n475) );
  XNOR2_X1 U583 ( .A(n478), .B(G134), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n481), .B(G137), .ZN(n500) );
  NAND2_X1 U585 ( .A1(n765), .A2(G227), .ZN(n482) );
  XNOR2_X1 U586 ( .A(n482), .B(G140), .ZN(n484) );
  XNOR2_X1 U587 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U588 ( .A(n486), .B(n485), .ZN(n487) );
  BUF_X1 U589 ( .A(n488), .Z(n489) );
  XNOR2_X1 U590 ( .A(n491), .B(n490), .ZN(n494) );
  NAND2_X1 U591 ( .A1(n492), .A2(G210), .ZN(n493) );
  XNOR2_X1 U592 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U593 ( .A(n489), .B(n495), .ZN(n496) );
  XNOR2_X1 U594 ( .A(n497), .B(n496), .ZN(n647) );
  XNOR2_X2 U595 ( .A(n498), .B(G472), .ZN(n695) );
  XNOR2_X1 U596 ( .A(n695), .B(KEYINPUT103), .ZN(n576) );
  XNOR2_X1 U597 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U598 ( .A(n504), .B(n503), .Z(n508) );
  NAND2_X1 U599 ( .A1(G221), .A2(n505), .ZN(n506) );
  XNOR2_X1 U600 ( .A(n756), .B(n506), .ZN(n507) );
  NOR2_X1 U601 ( .A1(G902), .A2(n736), .ZN(n513) );
  NAND2_X1 U602 ( .A1(n509), .A2(G217), .ZN(n511) );
  INV_X1 U603 ( .A(KEYINPUT25), .ZN(n510) );
  XNOR2_X1 U604 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U605 ( .A(n513), .B(n512), .ZN(n515) );
  BUF_X1 U606 ( .A(n515), .Z(n690) );
  NAND2_X1 U607 ( .A1(n576), .A2(n690), .ZN(n514) );
  XNOR2_X1 U608 ( .A(n560), .B(G110), .ZN(G12) );
  XNOR2_X2 U609 ( .A(n516), .B(KEYINPUT69), .ZN(n687) );
  INV_X1 U610 ( .A(n580), .ZN(n517) );
  NAND2_X1 U611 ( .A1(n687), .A2(n517), .ZN(n543) );
  NOR2_X1 U612 ( .A1(G900), .A2(n518), .ZN(n519) );
  NAND2_X1 U613 ( .A1(G953), .A2(n519), .ZN(n520) );
  XNOR2_X1 U614 ( .A(KEYINPUT104), .B(n520), .ZN(n521) );
  NAND2_X1 U615 ( .A1(n522), .A2(n521), .ZN(n524) );
  INV_X1 U616 ( .A(KEYINPUT80), .ZN(n523) );
  XNOR2_X1 U617 ( .A(n524), .B(n523), .ZN(n572) );
  NOR2_X1 U618 ( .A1(n543), .A2(n572), .ZN(n528) );
  INV_X1 U619 ( .A(KEYINPUT30), .ZN(n525) );
  XNOR2_X1 U620 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U621 ( .A1(n528), .A2(n527), .ZN(n607) );
  BUF_X1 U622 ( .A(n529), .Z(n604) );
  INV_X1 U623 ( .A(KEYINPUT38), .ZN(n530) );
  XNOR2_X1 U624 ( .A(n604), .B(n530), .ZN(n568) );
  INV_X1 U625 ( .A(KEYINPUT39), .ZN(n531) );
  XNOR2_X1 U626 ( .A(n532), .B(n531), .ZN(n534) );
  INV_X1 U627 ( .A(n555), .ZN(n533) );
  OR2_X1 U628 ( .A1(n556), .A2(n533), .ZN(n665) );
  OR2_X1 U629 ( .A1(n534), .A2(n665), .ZN(n623) );
  XNOR2_X1 U630 ( .A(n623), .B(G134), .ZN(G36) );
  AND2_X1 U631 ( .A1(n556), .A2(n533), .ZN(n674) );
  INV_X1 U632 ( .A(n674), .ZN(n589) );
  OR2_X2 U633 ( .A1(n534), .A2(n589), .ZN(n536) );
  XNOR2_X1 U634 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n535) );
  XOR2_X1 U635 ( .A(G131), .B(n585), .Z(G33) );
  INV_X1 U636 ( .A(n690), .ZN(n573) );
  AND2_X1 U637 ( .A1(n589), .A2(n665), .ZN(n702) );
  NAND2_X1 U638 ( .A1(n687), .A2(n695), .ZN(n539) );
  NAND2_X1 U639 ( .A1(n540), .A2(n697), .ZN(n541) );
  NOR2_X1 U640 ( .A1(n543), .A2(n695), .ZN(n544) );
  NOR2_X1 U641 ( .A1(n702), .A2(n545), .ZN(n546) );
  INV_X1 U642 ( .A(n550), .ZN(n591) );
  AND2_X1 U643 ( .A1(n687), .A2(n591), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U645 ( .A(n553), .B(KEYINPUT33), .ZN(n709) );
  AND2_X1 U646 ( .A1(n556), .A2(n555), .ZN(n605) );
  AND2_X1 U647 ( .A1(n551), .A2(n690), .ZN(n559) );
  NAND2_X1 U648 ( .A1(n561), .A2(KEYINPUT44), .ZN(n562) );
  INV_X1 U649 ( .A(n653), .ZN(n565) );
  INV_X1 U650 ( .A(KEYINPUT44), .ZN(n564) );
  AND2_X1 U651 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U652 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n567) );
  INV_X1 U653 ( .A(KEYINPUT41), .ZN(n571) );
  INV_X1 U654 ( .A(n568), .ZN(n704) );
  INV_X1 U655 ( .A(n569), .ZN(n703) );
  NAND2_X1 U656 ( .A1(n704), .A2(n703), .ZN(n701) );
  OR2_X1 U657 ( .A1(n706), .A2(n701), .ZN(n570) );
  XNOR2_X1 U658 ( .A(n571), .B(n570), .ZN(n719) );
  NOR2_X1 U659 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U660 ( .A1(n575), .A2(n574), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n588), .A2(n576), .ZN(n577) );
  XNOR2_X1 U662 ( .A(KEYINPUT28), .B(n577), .ZN(n596) );
  INV_X1 U663 ( .A(n596), .ZN(n578) );
  NOR2_X1 U664 ( .A1(n719), .A2(n578), .ZN(n581) );
  INV_X1 U665 ( .A(KEYINPUT108), .ZN(n579) );
  XNOR2_X1 U666 ( .A(n580), .B(n579), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n581), .A2(n597), .ZN(n584) );
  INV_X1 U668 ( .A(KEYINPUT110), .ZN(n582) );
  XNOR2_X1 U669 ( .A(n582), .B(KEYINPUT42), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n584), .B(n583), .ZN(n770) );
  INV_X1 U671 ( .A(KEYINPUT46), .ZN(n586) );
  XNOR2_X1 U672 ( .A(n587), .B(n586), .ZN(n615) );
  NOR2_X1 U673 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U674 ( .A1(n590), .A2(n703), .ZN(n592) );
  NAND2_X1 U675 ( .A1(n592), .A2(n591), .ZN(n618) );
  NOR2_X1 U676 ( .A1(n618), .A2(n604), .ZN(n593) );
  XNOR2_X1 U677 ( .A(n593), .B(KEYINPUT36), .ZN(n594) );
  NAND2_X1 U678 ( .A1(n594), .A2(n551), .ZN(n682) );
  XNOR2_X1 U679 ( .A(n682), .B(KEYINPUT86), .ZN(n603) );
  AND2_X1 U680 ( .A1(n367), .A2(n596), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U682 ( .A(n599), .B(KEYINPUT47), .ZN(n601) );
  INV_X1 U683 ( .A(n599), .ZN(n672) );
  NAND2_X1 U684 ( .A1(n672), .A2(n702), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n605), .A2(n368), .ZN(n606) );
  OR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n609) );
  INV_X1 U689 ( .A(KEYINPUT107), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n609), .B(n608), .ZN(n771) );
  NAND2_X1 U691 ( .A1(n702), .A2(KEYINPUT47), .ZN(n610) );
  AND2_X1 U692 ( .A1(n771), .A2(n610), .ZN(n611) );
  XNOR2_X1 U693 ( .A(n611), .B(KEYINPUT81), .ZN(n612) );
  NOR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n617) );
  INV_X1 U696 ( .A(KEYINPUT48), .ZN(n616) );
  XNOR2_X1 U697 ( .A(n617), .B(n616), .ZN(n625) );
  NOR2_X1 U698 ( .A1(n618), .A2(n551), .ZN(n620) );
  XOR2_X1 U699 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n619) );
  XNOR2_X1 U700 ( .A(n620), .B(n619), .ZN(n621) );
  OR2_X1 U701 ( .A1(n621), .A2(n368), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n622), .B(KEYINPUT106), .ZN(n772) );
  AND2_X1 U703 ( .A1(n772), .A2(n623), .ZN(n624) );
  AND2_X2 U704 ( .A1(n746), .A2(n759), .ZN(n685) );
  NAND2_X1 U705 ( .A1(n685), .A2(KEYINPUT2), .ZN(n627) );
  INV_X1 U706 ( .A(KEYINPUT78), .ZN(n626) );
  XNOR2_X2 U707 ( .A(n627), .B(n626), .ZN(n684) );
  INV_X1 U708 ( .A(n635), .ZN(n630) );
  NAND2_X1 U709 ( .A1(KEYINPUT2), .A2(KEYINPUT85), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n628), .A2(KEYINPUT84), .ZN(n629) );
  NOR2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n637) );
  INV_X1 U712 ( .A(n637), .ZN(n631) );
  AND2_X1 U713 ( .A1(KEYINPUT84), .A2(n631), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n685), .A2(n632), .ZN(n639) );
  INV_X1 U715 ( .A(KEYINPUT2), .ZN(n633) );
  NOR2_X1 U716 ( .A1(n633), .A2(KEYINPUT85), .ZN(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  OR2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n641) );
  NOR2_X1 U720 ( .A1(n685), .A2(KEYINPUT84), .ZN(n640) );
  BUF_X1 U721 ( .A(n643), .Z(n644) );
  XNOR2_X1 U722 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n645) );
  INV_X1 U723 ( .A(G952), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n730), .A2(G472), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X2 U726 ( .A1(n650), .A2(n740), .ZN(n652) );
  XOR2_X1 U727 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(G57) );
  XOR2_X1 U729 ( .A(G122), .B(n359), .Z(G24) );
  BUF_X1 U730 ( .A(n654), .Z(n655) );
  XNOR2_X1 U731 ( .A(G119), .B(KEYINPUT126), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n655), .B(n656), .ZN(G21) );
  NAND2_X1 U733 ( .A1(n730), .A2(G475), .ZN(n660) );
  XOR2_X1 U734 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n657) );
  XNOR2_X1 U735 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X2 U736 ( .A1(n661), .A2(n740), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n662), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U738 ( .A(G101), .B(n663), .Z(G3) );
  NAND2_X1 U739 ( .A1(n666), .A2(n674), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n664), .B(G104), .ZN(G6) );
  XOR2_X1 U741 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n668) );
  INV_X1 U742 ( .A(n665), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n666), .A2(n677), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U745 ( .A(G107), .B(n669), .ZN(G9) );
  XOR2_X1 U746 ( .A(G128), .B(KEYINPUT29), .Z(n671) );
  NAND2_X1 U747 ( .A1(n672), .A2(n677), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n671), .B(n670), .ZN(G30) );
  NAND2_X1 U749 ( .A1(n672), .A2(n674), .ZN(n673) );
  XNOR2_X1 U750 ( .A(n673), .B(G146), .ZN(G48) );
  NAND2_X1 U751 ( .A1(n678), .A2(n674), .ZN(n676) );
  XNOR2_X1 U752 ( .A(n676), .B(n675), .ZN(G15) );
  XOR2_X1 U753 ( .A(G116), .B(KEYINPUT111), .Z(n680) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n680), .B(n679), .ZN(G18) );
  XOR2_X1 U756 ( .A(KEYINPUT37), .B(KEYINPUT112), .Z(n681) );
  XNOR2_X1 U757 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U758 ( .A(G125), .B(n683), .ZN(G27) );
  XNOR2_X1 U759 ( .A(KEYINPUT82), .B(KEYINPUT2), .ZN(n686) );
  NOR2_X1 U760 ( .A1(n551), .A2(n687), .ZN(n688) );
  XOR2_X1 U761 ( .A(KEYINPUT50), .B(n688), .Z(n694) );
  NAND2_X1 U762 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U763 ( .A(n691), .B(KEYINPUT113), .ZN(n692) );
  XNOR2_X1 U764 ( .A(KEYINPUT49), .B(n692), .ZN(n693) );
  NAND2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n696) );
  NOR2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n698) );
  NOR2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U768 ( .A(KEYINPUT51), .B(n699), .Z(n700) );
  NOR2_X1 U769 ( .A1(n719), .A2(n700), .ZN(n712) );
  NOR2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n710) );
  INV_X1 U774 ( .A(n709), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n710), .A2(n718), .ZN(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U777 ( .A(n713), .B(KEYINPUT52), .ZN(n714) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U779 ( .A(n716), .B(KEYINPUT114), .ZN(n717) );
  NOR2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U781 ( .A(KEYINPUT53), .B(KEYINPUT116), .ZN(n722) );
  XNOR2_X1 U782 ( .A(n723), .B(n722), .ZN(G75) );
  NAND2_X1 U783 ( .A1(n734), .A2(G469), .ZN(n728) );
  XOR2_X1 U784 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n724) );
  XNOR2_X1 U785 ( .A(n724), .B(KEYINPUT118), .ZN(n725) );
  XNOR2_X1 U786 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U787 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U788 ( .A1(n740), .A2(n729), .ZN(G54) );
  NAND2_X1 U789 ( .A1(n385), .A2(G478), .ZN(n731) );
  XOR2_X1 U790 ( .A(n732), .B(n731), .Z(n733) );
  NOR2_X1 U791 ( .A1(n740), .A2(n733), .ZN(G63) );
  NAND2_X1 U792 ( .A1(n734), .A2(G217), .ZN(n738) );
  INV_X1 U793 ( .A(KEYINPUT119), .ZN(n735) );
  NOR2_X1 U794 ( .A1(n740), .A2(n739), .ZN(G66) );
  XOR2_X1 U795 ( .A(n743), .B(n742), .Z(n745) );
  NOR2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n755) );
  BUF_X1 U797 ( .A(n746), .Z(n747) );
  NAND2_X1 U798 ( .A1(n747), .A2(n765), .ZN(n753) );
  XOR2_X1 U799 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n749) );
  NAND2_X1 U800 ( .A1(G224), .A2(G953), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U804 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U805 ( .A(n755), .B(n754), .ZN(G69) );
  XNOR2_X1 U806 ( .A(n757), .B(n756), .ZN(n761) );
  XNOR2_X1 U807 ( .A(n761), .B(KEYINPUT122), .ZN(n758) );
  XNOR2_X1 U808 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U809 ( .A1(G953), .A2(n760), .ZN(n768) );
  XNOR2_X1 U810 ( .A(n761), .B(G227), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n762), .A2(G900), .ZN(n763) );
  XNOR2_X1 U812 ( .A(KEYINPUT123), .B(n763), .ZN(n764) );
  NOR2_X1 U813 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U814 ( .A(n766), .B(KEYINPUT124), .ZN(n767) );
  NOR2_X1 U815 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U816 ( .A(KEYINPUT125), .B(n769), .ZN(G72) );
  XOR2_X1 U817 ( .A(G137), .B(n770), .Z(G39) );
  XNOR2_X1 U818 ( .A(n353), .B(n771), .ZN(G45) );
  XNOR2_X1 U819 ( .A(G140), .B(n772), .ZN(G42) );
endmodule

