//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n191), .A2(new_n192), .B1(new_n189), .B2(new_n190), .ZN(new_n193));
  INV_X1    g007(.A(G116), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT70), .B1(new_n194), .B2(G119), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(G119), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n193), .B(new_n200), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT66), .A2(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(G137), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n202), .A2(KEYINPUT11), .A3(G134), .A4(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT11), .B1(new_n205), .B2(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(G134), .B1(new_n202), .B2(new_n203), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(G134), .B2(new_n205), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT64), .A2(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT64), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n214), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT64), .A2(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT64), .A2(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(G143), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(G128), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G143), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n215), .A2(new_n216), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n221), .A2(KEYINPUT65), .A3(G143), .A4(new_n222), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT65), .B1(new_n226), .B2(G143), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n231), .B(new_n233), .C1(new_n218), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT67), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n223), .A2(new_n234), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n238), .A2(new_n239), .A3(new_n231), .A4(new_n233), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n213), .B1(new_n230), .B2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n238), .A2(KEYINPUT0), .A3(G128), .A4(new_n231), .ZN(new_n243));
  XOR2_X1   g057(.A(KEYINPUT0), .B(G128), .Z(new_n244));
  NAND2_X1  g058(.A1(new_n229), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n210), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n209), .B1(new_n204), .B2(new_n208), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n243), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT30), .B1(new_n242), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n229), .A2(new_n225), .B1(new_n237), .B2(new_n240), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n251), .B(new_n248), .C1(new_n252), .C2(new_n213), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n201), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n256), .B(KEYINPUT27), .Z(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n201), .B(new_n248), .C1(new_n252), .C2(new_n213), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n254), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n187), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n201), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n242), .B2(new_n249), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n268), .B2(new_n260), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI211_X1 g085(.A(KEYINPUT73), .B(new_n265), .C1(new_n268), .C2(new_n260), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n259), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n213), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n237), .A2(new_n240), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n232), .B1(new_n276), .B2(new_n214), .ZN(new_n277));
  INV_X1    g091(.A(new_n228), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n217), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n277), .A2(new_n224), .B1(new_n227), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n274), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n251), .B1(new_n281), .B2(new_n248), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n242), .A2(KEYINPUT30), .A3(new_n249), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n267), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n259), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n260), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n288));
  NAND2_X1  g102(.A1(new_n262), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n264), .A2(new_n273), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT74), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n290), .A2(new_n295), .A3(new_n291), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n290), .A2(KEYINPUT75), .A3(KEYINPUT32), .A4(new_n291), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n269), .B1(new_n265), .B2(new_n260), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n259), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n284), .A2(new_n260), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n259), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n304), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n271), .A2(new_n259), .A3(new_n272), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G472), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n297), .A2(new_n302), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT9), .B(G234), .ZN(new_n314));
  OAI21_X1  g128(.A(G221), .B1(new_n314), .B2(G902), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n230), .A2(new_n241), .ZN(new_n316));
  INV_X1    g130(.A(G104), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G107), .ZN(new_n318));
  INV_X1    g132(.A(G107), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G104), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n317), .A2(G107), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT77), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n325), .A3(KEYINPUT3), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n321), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G101), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n320), .A2(new_n318), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G101), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n316), .A2(KEYINPUT10), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n321), .ZN(new_n335));
  INV_X1    g149(.A(new_n326), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n325), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G101), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n329), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n243), .A2(new_n245), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n324), .A2(new_n326), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n328), .B1(new_n342), .B2(new_n335), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT78), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n346));
  NOR4_X1   g160(.A1(new_n327), .A2(new_n346), .A3(KEYINPUT4), .A4(new_n328), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n340), .B(new_n341), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n238), .A2(new_n231), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n232), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n352), .B2(new_n351), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n237), .A2(new_n240), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n349), .B1(new_n355), .B2(new_n332), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n334), .A2(new_n348), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n246), .A2(new_n247), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G110), .B(G140), .ZN(new_n360));
  INV_X1    g174(.A(G227), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G953), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n360), .B(new_n362), .Z(new_n363));
  NAND3_X1  g177(.A1(new_n334), .A2(new_n348), .A3(new_n356), .ZN(new_n364));
  INV_X1    g178(.A(new_n358), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n316), .A2(new_n333), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n355), .A2(new_n332), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n252), .A2(new_n332), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n354), .A2(new_n350), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n241), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n333), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n358), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT12), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n372), .A2(new_n378), .B1(new_n357), .B2(new_n358), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n367), .B(G469), .C1(new_n379), .C2(new_n363), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g195(.A1(G469), .A2(G902), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n370), .A2(new_n371), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n377), .A2(KEYINPUT12), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n359), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n363), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  INV_X1    g202(.A(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n363), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n359), .A2(new_n390), .A3(new_n366), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n387), .A2(new_n388), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n383), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n315), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(G214), .B1(G237), .B2(G902), .ZN(new_n396));
  OAI21_X1  g210(.A(G210), .B1(G237), .B2(G902), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n397), .B(KEYINPUT85), .Z(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n340), .B(new_n267), .C1(new_n345), .C2(new_n347), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n193), .A2(new_n198), .A3(new_n199), .A4(new_n195), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n195), .A2(new_n198), .A3(KEYINPUT5), .A4(new_n199), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n194), .A2(KEYINPUT5), .A3(G119), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n190), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n333), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G122), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n400), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G953), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G224), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT7), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(G125), .B1(new_n230), .B2(new_n241), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n243), .A2(G125), .A3(new_n245), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n402), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n404), .B1(new_n402), .B2(new_n417), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n401), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n333), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n408), .B(KEYINPUT8), .Z(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n406), .B2(new_n332), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n409), .A2(new_n416), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G125), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n415), .B1(new_n316), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT83), .A3(new_n412), .ZN(new_n428));
  INV_X1    g242(.A(new_n415), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n429), .B(new_n412), .C1(new_n252), .C2(G125), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  AOI211_X1 g247(.A(KEYINPUT84), .B(G902), .C1(new_n425), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n429), .B1(new_n252), .B2(G125), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n436), .A2(new_n413), .B1(new_n421), .B2(new_n423), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT83), .B1(new_n427), .B2(new_n412), .ZN(new_n438));
  NOR4_X1   g252(.A1(new_n414), .A2(new_n415), .A3(new_n431), .A4(new_n413), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n437), .B(new_n409), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n435), .B1(new_n440), .B2(new_n389), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n409), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n408), .B(KEYINPUT81), .Z(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n400), .B2(new_n407), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT6), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n445), .A2(KEYINPUT6), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n436), .B(new_n411), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n399), .B1(new_n442), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n440), .A2(new_n389), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n440), .A2(new_n435), .A3(new_n389), .ZN(new_n454));
  AND4_X1   g268(.A1(new_n399), .A2(new_n453), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n396), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G125), .B(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n228), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n226), .B2(new_n457), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT87), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n458), .B(new_n461), .C1(new_n226), .C2(new_n457), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n464));
  INV_X1    g278(.A(G237), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n410), .A3(G214), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n217), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(KEYINPUT18), .A2(G131), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n468), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n472), .A2(KEYINPUT86), .A3(KEYINPUT18), .A4(G131), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n470), .B(KEYINPUT88), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT89), .B1(new_n469), .B2(new_n475), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n463), .B(new_n474), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n457), .A2(KEYINPUT16), .ZN(new_n481));
  OR3_X1    g295(.A1(new_n426), .A2(KEYINPUT16), .A3(G140), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(G146), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(G146), .B1(new_n481), .B2(new_n482), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n472), .A2(KEYINPUT17), .A3(G131), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n469), .A2(new_n209), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n472), .A2(G131), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n486), .B(new_n487), .C1(new_n490), .C2(KEYINPUT17), .ZN(new_n491));
  XNOR2_X1  g305(.A(G113), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n317), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n480), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n457), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT19), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n490), .B(new_n483), .C1(new_n278), .C2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n480), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n494), .B1(new_n499), .B2(new_n493), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n480), .A2(new_n491), .A3(new_n493), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n493), .B1(new_n480), .B2(new_n498), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n502), .B(new_n503), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT91), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  INV_X1    g323(.A(new_n503), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT20), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n493), .B1(new_n480), .B2(new_n491), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n389), .B1(new_n505), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(KEYINPUT92), .B(new_n389), .C1(new_n505), .C2(new_n513), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(G475), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(G234), .A2(G237), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n521), .A2(G952), .A3(new_n410), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n521), .A2(G902), .A3(G953), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT21), .B(G898), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n217), .B2(G128), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n232), .A2(KEYINPUT93), .A3(G143), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G134), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n217), .A2(G128), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G122), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G116), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n194), .A2(G122), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n319), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n538), .A3(new_n319), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT13), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n533), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n531), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n547), .B2(KEYINPUT94), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(KEYINPUT94), .B2(new_n547), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n543), .B1(new_n549), .B2(G134), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n532), .B1(new_n531), .B2(new_n533), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n541), .B1(new_n534), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT14), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n537), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n538), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(KEYINPUT14), .B2(new_n538), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G107), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(KEYINPUT95), .A3(G107), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n553), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G217), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n314), .A2(new_n564), .A3(G953), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n551), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n565), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n550), .B2(new_n562), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI211_X1 g383(.A(KEYINPUT15), .B(new_n527), .C1(new_n569), .C2(new_n389), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n389), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n520), .A2(new_n526), .A3(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n395), .A2(new_n456), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT23), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n197), .B2(G128), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n232), .A2(KEYINPUT23), .A3(G119), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n578), .B(new_n579), .C1(G119), .C2(new_n232), .ZN(new_n580));
  XNOR2_X1  g394(.A(G119), .B(G128), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT24), .B(G110), .Z(new_n582));
  AOI22_X1  g396(.A1(new_n580), .A2(G110), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n484), .B2(new_n485), .ZN(new_n584));
  OAI22_X1  g398(.A1(new_n580), .A2(G110), .B1(new_n581), .B2(new_n582), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n483), .A3(new_n458), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT22), .B(G137), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n410), .A2(G221), .A3(G234), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n587), .B(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT25), .A3(new_n389), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n587), .A2(new_n590), .ZN(new_n593));
  INV_X1    g407(.A(new_n590), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n584), .B2(new_n586), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n389), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n592), .A2(new_n598), .A3(KEYINPUT76), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n564), .B1(G234), .B2(new_n389), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n598), .B2(KEYINPUT76), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n591), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n313), .A2(new_n576), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT96), .B(G101), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  NAND2_X1  g422(.A1(new_n290), .A2(new_n389), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n609), .A2(KEYINPUT97), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(KEYINPUT97), .ZN(new_n611));
  OAI21_X1  g425(.A(G472), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n293), .A2(new_n296), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n605), .B(new_n315), .C1(new_n393), .C2(new_n394), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n456), .A2(KEYINPUT98), .ZN(new_n618));
  INV_X1    g432(.A(new_n396), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n453), .A2(new_n450), .A3(new_n454), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n398), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n442), .A2(new_n399), .A3(new_n450), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n569), .A2(KEYINPUT33), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n566), .B2(new_n568), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n389), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G478), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n571), .A2(G478), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n519), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n626), .A2(new_n526), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n617), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT99), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  NAND2_X1  g454(.A1(new_n511), .A2(new_n507), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n511), .A2(KEYINPUT100), .A3(new_n507), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n518), .B1(new_n570), .B2(new_n573), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n626), .A2(new_n526), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n617), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT35), .B(G107), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NOR2_X1   g465(.A1(new_n594), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n587), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n603), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(new_n599), .B2(new_n601), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n576), .A2(new_n612), .A3(new_n613), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(new_n655), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n618), .B2(new_n625), .ZN(new_n660));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n523), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n522), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n645), .A2(new_n646), .A3(new_n665), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n666), .B(new_n315), .C1(new_n394), .C2(new_n393), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n660), .A2(new_n313), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  INV_X1    g484(.A(new_n395), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n664), .B(KEYINPUT39), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n621), .A2(new_n622), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n520), .A2(new_n574), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n680), .A2(new_n619), .A3(new_n655), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n674), .A2(new_n675), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n297), .A2(new_n302), .ZN(new_n683));
  INV_X1    g497(.A(G472), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n389), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n285), .B1(new_n268), .B2(new_n260), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n684), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n685), .B1(new_n286), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT102), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n682), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n217), .ZN(G45));
  NOR2_X1   g507(.A1(new_n634), .A2(new_n665), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n694), .B(new_n315), .C1(new_n394), .C2(new_n393), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n660), .A2(new_n313), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT103), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n660), .A2(new_n699), .A3(new_n313), .A4(new_n696), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  INV_X1    g516(.A(new_n315), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n391), .B(new_n389), .C1(new_n379), .C2(new_n390), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n392), .A3(KEYINPUT104), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n704), .A2(new_n707), .A3(G469), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n703), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n313), .A2(new_n605), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(new_n636), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT105), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NOR2_X1   g528(.A1(new_n710), .A2(new_n648), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT106), .B(G116), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G18));
  INV_X1    g531(.A(new_n709), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n575), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n660), .A2(new_n313), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  NOR2_X1   g535(.A1(new_n718), .A2(new_n525), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n609), .A2(G472), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n289), .B1(new_n303), .B2(new_n285), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n262), .A2(new_n263), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n291), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n605), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n626), .A2(new_n722), .A3(new_n679), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  AND4_X1   g544(.A1(new_n655), .A2(new_n723), .A3(new_n694), .A4(new_n726), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n626), .A2(new_n731), .A3(new_n709), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  INV_X1    g547(.A(new_n605), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n292), .A2(new_n735), .A3(new_n294), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(new_n312), .A3(new_n298), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n292), .A2(new_n294), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT109), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n734), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n386), .A2(new_n390), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n386), .A2(new_n743), .A3(new_n390), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n742), .A2(G469), .A3(new_n367), .A4(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n745), .A2(new_n382), .A3(new_n392), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n621), .A2(new_n622), .A3(new_n315), .A4(new_n396), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n694), .A4(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n313), .A2(new_n605), .A3(new_n694), .A4(new_n748), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n749), .B(KEYINPUT110), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT111), .B(G131), .Z(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G33));
  NAND4_X1  g575(.A1(new_n313), .A2(new_n605), .A3(new_n666), .A4(new_n748), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  NOR2_X1   g577(.A1(new_n676), .A2(new_n619), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n520), .A2(new_n631), .A3(new_n633), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT43), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n614), .A2(new_n655), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n672), .ZN(new_n771));
  INV_X1    g585(.A(new_n392), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n742), .A2(KEYINPUT45), .A3(new_n367), .A4(new_n744), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n741), .A2(new_n367), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n773), .B(G469), .C1(KEYINPUT45), .C2(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(new_n382), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n772), .B1(new_n776), .B2(KEYINPUT46), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n382), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n703), .B(new_n771), .C1(new_n777), .C2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n770), .B(new_n781), .C1(new_n769), .C2(new_n768), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  NAND2_X1  g597(.A1(new_n694), .A2(new_n734), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n313), .A2(new_n765), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n777), .A2(new_n780), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT47), .B1(new_n786), .B2(new_n315), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n788), .B(new_n703), .C1(new_n777), .C2(new_n780), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NOR2_X1   g605(.A1(new_n787), .A2(new_n789), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n706), .A2(new_n708), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n703), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n767), .A2(new_n728), .A3(new_n522), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n765), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n796), .A2(new_n396), .A3(new_n678), .A4(new_n718), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT50), .ZN(new_n800));
  INV_X1    g614(.A(new_n747), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n767), .A2(new_n522), .A3(new_n793), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n655), .A2(new_n803), .A3(new_n723), .A4(new_n726), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n605), .A2(new_n801), .A3(new_n522), .A4(new_n793), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n691), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n519), .B1(new_n631), .B2(new_n633), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n798), .A2(new_n800), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n798), .A2(KEYINPUT51), .A3(new_n800), .A4(new_n809), .ZN(new_n813));
  INV_X1    g627(.A(new_n626), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n796), .A2(new_n814), .A3(new_n718), .ZN(new_n815));
  INV_X1    g629(.A(G952), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n816), .A3(G953), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n634), .B2(new_n806), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n803), .A2(new_n819), .A3(new_n740), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n819), .B1(new_n803), .B2(new_n740), .ZN(new_n822));
  OR3_X1    g636(.A1(new_n821), .A2(KEYINPUT48), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT48), .B1(new_n821), .B2(new_n822), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n812), .A2(new_n813), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT116), .Z(new_n827));
  NAND2_X1  g641(.A1(new_n669), .A2(new_n732), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n700), .B2(new_n698), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n814), .A2(new_n680), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n746), .A2(new_n703), .A3(new_n655), .A4(new_n665), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n690), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n669), .A2(new_n732), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n701), .A2(KEYINPUT52), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n729), .B(new_n720), .C1(new_n636), .C2(new_n710), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n634), .B1(new_n519), .B2(new_n574), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n623), .A2(new_n526), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n615), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n612), .A3(new_n613), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n656), .A2(new_n606), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n655), .A2(new_n574), .A3(new_n518), .A4(new_n664), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n645), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n396), .A3(new_n621), .A4(new_n622), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n395), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n313), .A2(new_n848), .B1(new_n731), .B2(new_n748), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n762), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n838), .A2(new_n844), .A3(new_n850), .A4(new_n715), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n757), .A2(new_n851), .A3(new_n758), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT53), .B1(new_n837), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n835), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n701), .A2(new_n832), .A3(new_n834), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n829), .A2(KEYINPUT113), .A3(KEYINPUT52), .A4(new_n832), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n860), .B(new_n861), .C1(new_n852), .C2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n757), .A2(new_n851), .A3(new_n758), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(KEYINPUT112), .ZN(new_n865));
  OAI211_X1 g679(.A(KEYINPUT54), .B(new_n853), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n861), .B1(new_n837), .B2(new_n852), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  INV_X1    g682(.A(new_n715), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n729), .A2(new_n720), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n711), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT114), .B1(new_n838), .B2(new_n715), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n844), .A2(new_n850), .A3(new_n861), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n755), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n860), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n867), .A2(new_n868), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n866), .A2(new_n877), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n827), .A2(new_n878), .B1(G952), .B2(G953), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n793), .B(KEYINPUT49), .Z(new_n880));
  NAND4_X1  g694(.A1(new_n766), .A2(new_n605), .A3(new_n315), .A4(new_n396), .ZN(new_n881));
  OR4_X1    g695(.A1(new_n690), .A2(new_n880), .A3(new_n678), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(G75));
  XNOR2_X1  g697(.A(new_n449), .B(KEYINPUT55), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n448), .B(KEYINPUT117), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n389), .B1(new_n867), .B2(new_n876), .ZN(new_n888));
  AOI211_X1 g702(.A(KEYINPUT56), .B(new_n887), .C1(new_n888), .C2(new_n398), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n858), .A2(new_n835), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n864), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n860), .A2(new_n875), .ZN(new_n892));
  OAI211_X1 g706(.A(G902), .B(new_n398), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n885), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n389), .B(new_n399), .C1(new_n867), .C2(new_n876), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n887), .B1(new_n897), .B2(KEYINPUT56), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n893), .A2(new_n894), .A3(new_n886), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n899), .A3(new_n884), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n410), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n896), .A2(new_n900), .A3(new_n902), .ZN(G51));
  OAI21_X1  g717(.A(KEYINPUT54), .B1(new_n891), .B2(new_n892), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n877), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n382), .B(KEYINPUT57), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n387), .B(new_n391), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n775), .B(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n888), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n901), .B1(new_n908), .B2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n912), .A2(KEYINPUT119), .A3(new_n509), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT119), .B1(new_n912), .B2(new_n509), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n901), .B1(new_n912), .B2(new_n509), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G60));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n627), .A2(new_n629), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT59), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n878), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n918), .A2(new_n921), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n867), .A2(new_n868), .A3(new_n876), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n868), .B1(new_n867), .B2(new_n876), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n902), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n917), .B1(new_n922), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n901), .B1(new_n905), .B2(new_n923), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n920), .B1(new_n866), .B2(new_n877), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n929), .B(KEYINPUT120), .C1(new_n918), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n867), .B2(new_n876), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n653), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n936), .B(new_n902), .C1(new_n591), .C2(new_n935), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G66));
  NOR3_X1   g753(.A1(new_n838), .A2(new_n715), .A3(new_n844), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT121), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n941), .A2(KEYINPUT122), .A3(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT122), .B1(new_n941), .B2(G953), .ZN(new_n943));
  INV_X1    g757(.A(G224), .ZN(new_n944));
  OAI21_X1  g758(.A(G953), .B1(new_n524), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n887), .B1(G898), .B2(new_n410), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  NAND3_X1  g762(.A1(new_n781), .A2(new_n830), .A3(new_n740), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n790), .A2(new_n782), .A3(new_n762), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n701), .A2(new_n834), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n759), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n410), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n250), .A2(new_n253), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n497), .B(KEYINPUT123), .Z(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(G900), .B2(G953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n673), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n764), .A2(new_n839), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n313), .A3(new_n605), .A4(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n790), .A2(new_n782), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n951), .A2(new_n692), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n969), .B(new_n963), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n410), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n959), .B1(new_n971), .B2(new_n956), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n410), .B1(G227), .B2(G900), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n958), .B2(KEYINPUT125), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G72));
  XOR2_X1   g789(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(new_n685), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n968), .A2(new_n970), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n941), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n307), .A2(new_n285), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n853), .B1(new_n863), .B2(new_n865), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n308), .B(KEYINPUT127), .Z(new_n983));
  AOI211_X1 g797(.A(new_n977), .B(new_n982), .C1(new_n286), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n977), .B1(new_n952), .B2(new_n941), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n284), .A2(new_n259), .A3(new_n260), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n902), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n981), .A2(new_n984), .A3(new_n987), .ZN(G57));
endmodule


