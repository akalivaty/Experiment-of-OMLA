

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599;

  XNOR2_X1 U325 ( .A(n312), .B(n311), .ZN(n318) );
  NOR2_X1 U326 ( .A1(n514), .A2(n513), .ZN(n521) );
  XOR2_X1 U327 ( .A(G218GAT), .B(G162GAT), .Z(n293) );
  NOR2_X1 U328 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U329 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n415) );
  INV_X1 U330 ( .A(KEYINPUT27), .ZN(n471) );
  XNOR2_X1 U331 ( .A(n416), .B(n415), .ZN(n418) );
  XNOR2_X1 U332 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U333 ( .A(n471), .B(KEYINPUT100), .ZN(n472) );
  NOR2_X1 U334 ( .A1(n486), .A2(n485), .ZN(n487) );
  NOR2_X1 U335 ( .A1(n540), .A2(n429), .ZN(n579) );
  XNOR2_X1 U336 ( .A(n473), .B(n472), .ZN(n481) );
  XNOR2_X1 U337 ( .A(KEYINPUT105), .B(KEYINPUT36), .ZN(n358) );
  XNOR2_X1 U338 ( .A(n406), .B(n358), .ZN(n597) );
  NOR2_X1 U339 ( .A1(n557), .A2(n556), .ZN(n566) );
  XOR2_X1 U340 ( .A(KEYINPUT112), .B(n526), .Z(n532) );
  XNOR2_X1 U341 ( .A(n463), .B(n462), .ZN(n537) );
  XNOR2_X1 U342 ( .A(n465), .B(G190GAT), .ZN(n466) );
  XNOR2_X1 U343 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  XOR2_X1 U344 ( .A(G92GAT), .B(G106GAT), .Z(n294) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U346 ( .A(KEYINPUT82), .B(KEYINPUT79), .Z(n296) );
  XNOR2_X1 U347 ( .A(KEYINPUT78), .B(KEYINPUT65), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n305) );
  INV_X1 U350 ( .A(n305), .ZN(n303) );
  XOR2_X1 U351 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n300) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U354 ( .A(KEYINPUT9), .B(n301), .ZN(n304) );
  INV_X1 U355 ( .A(n304), .ZN(n302) );
  NAND2_X1 U356 ( .A1(n303), .A2(n302), .ZN(n307) );
  NAND2_X1 U357 ( .A1(n305), .A2(n304), .ZN(n306) );
  NAND2_X1 U358 ( .A1(n307), .A2(n306), .ZN(n312) );
  XOR2_X1 U359 ( .A(G134GAT), .B(KEYINPUT80), .Z(n334) );
  XOR2_X1 U360 ( .A(G190GAT), .B(KEYINPUT81), .Z(n419) );
  XOR2_X1 U361 ( .A(n334), .B(n419), .Z(n310) );
  XOR2_X1 U362 ( .A(G99GAT), .B(G85GAT), .Z(n308) );
  XNOR2_X1 U363 ( .A(KEYINPUT76), .B(n308), .ZN(n396) );
  INV_X1 U364 ( .A(n396), .ZN(n309) );
  XNOR2_X1 U365 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n313), .B(G29GAT), .ZN(n314) );
  XOR2_X1 U367 ( .A(n314), .B(KEYINPUT8), .Z(n316) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(G50GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n353) );
  INV_X1 U370 ( .A(n353), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n406) );
  INV_X1 U372 ( .A(n406), .ZN(n552) );
  XOR2_X1 U373 ( .A(KEYINPUT93), .B(G162GAT), .Z(n320) );
  XNOR2_X1 U374 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U376 ( .A(KEYINPUT3), .B(n321), .Z(n441) );
  XOR2_X1 U377 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n323) );
  XNOR2_X1 U378 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U380 ( .A(KEYINPUT98), .B(KEYINPUT4), .Z(n325) );
  XNOR2_X1 U381 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U383 ( .A(n327), .B(n326), .Z(n340) );
  XNOR2_X1 U384 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n328), .B(G127GAT), .ZN(n453) );
  XOR2_X1 U386 ( .A(n453), .B(KEYINPUT97), .Z(n330) );
  NAND2_X1 U387 ( .A1(G225GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n338) );
  XOR2_X1 U389 ( .A(G57GAT), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U390 ( .A(G141GAT), .B(G120GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U392 ( .A(n333), .B(G85GAT), .Z(n336) );
  XNOR2_X1 U393 ( .A(G29GAT), .B(n334), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n441), .B(n341), .ZN(n540) );
  XOR2_X1 U398 ( .A(KEYINPUT72), .B(KEYINPUT67), .Z(n343) );
  XNOR2_X1 U399 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n357) );
  XOR2_X1 U401 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n345) );
  XNOR2_X1 U402 ( .A(KEYINPUT68), .B(KEYINPUT71), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U404 ( .A(n346), .B(G197GAT), .Z(n348) );
  XOR2_X1 U405 ( .A(G15GAT), .B(G1GAT), .Z(n360) );
  XNOR2_X1 U406 ( .A(n360), .B(G113GAT), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U408 ( .A(G169GAT), .B(G8GAT), .Z(n423) );
  XOR2_X1 U409 ( .A(n423), .B(KEYINPUT29), .Z(n350) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U412 ( .A(n352), .B(n351), .Z(n355) );
  XOR2_X1 U413 ( .A(G141GAT), .B(G22GAT), .Z(n433) );
  XNOR2_X1 U414 ( .A(n353), .B(n433), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U416 ( .A(n357), .B(n356), .Z(n582) );
  XNOR2_X1 U417 ( .A(n582), .B(KEYINPUT73), .ZN(n569) );
  INV_X1 U418 ( .A(n569), .ZN(n545) );
  XNOR2_X1 U419 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n359), .B(KEYINPUT74), .ZN(n388) );
  XOR2_X1 U421 ( .A(n388), .B(n360), .Z(n362) );
  NAND2_X1 U422 ( .A1(G231GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n378) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n364) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(KEYINPUT15), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n376) );
  XOR2_X1 U427 ( .A(G71GAT), .B(G127GAT), .Z(n366) );
  XNOR2_X1 U428 ( .A(G22GAT), .B(G183GAT), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n374) );
  XOR2_X1 U430 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n368) );
  XNOR2_X1 U431 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U433 ( .A(G64GAT), .B(G78GAT), .Z(n370) );
  XNOR2_X1 U434 ( .A(G211GAT), .B(G155GAT), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U436 ( .A(n372), .B(n371), .Z(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U438 ( .A(n376), .B(n375), .Z(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n577) );
  NOR2_X1 U440 ( .A1(n597), .A2(n577), .ZN(n379) );
  XNOR2_X1 U441 ( .A(KEYINPUT45), .B(n379), .ZN(n399) );
  INV_X1 U442 ( .A(KEYINPUT32), .ZN(n380) );
  NAND2_X1 U443 ( .A1(KEYINPUT77), .A2(n380), .ZN(n383) );
  INV_X1 U444 ( .A(KEYINPUT77), .ZN(n381) );
  NAND2_X1 U445 ( .A1(n381), .A2(KEYINPUT32), .ZN(n382) );
  NAND2_X1 U446 ( .A1(n383), .A2(n382), .ZN(n385) );
  NAND2_X1 U447 ( .A1(G230GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U449 ( .A(KEYINPUT33), .B(n386), .Z(n390) );
  XNOR2_X1 U450 ( .A(G176GAT), .B(G92GAT), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n387), .B(G64GAT), .ZN(n412) );
  XNOR2_X1 U452 ( .A(n412), .B(n388), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n391), .B(KEYINPUT31), .ZN(n393) );
  XOR2_X1 U455 ( .A(G120GAT), .B(G71GAT), .Z(n450) );
  XOR2_X1 U456 ( .A(n450), .B(G204GAT), .Z(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U458 ( .A(G78GAT), .B(G148GAT), .Z(n395) );
  XNOR2_X1 U459 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n436) );
  XNOR2_X1 U461 ( .A(n436), .B(n396), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n398), .B(n397), .ZN(n587) );
  INV_X1 U463 ( .A(n587), .ZN(n402) );
  AND2_X1 U464 ( .A1(n399), .A2(n402), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n400), .B(KEYINPUT115), .ZN(n401) );
  NOR2_X1 U466 ( .A1(n545), .A2(n401), .ZN(n410) );
  XOR2_X1 U467 ( .A(n402), .B(KEYINPUT41), .Z(n574) );
  INV_X1 U468 ( .A(n574), .ZN(n403) );
  NAND2_X1 U469 ( .A1(n582), .A2(n403), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n404), .B(KEYINPUT46), .ZN(n405) );
  NAND2_X1 U471 ( .A1(n405), .A2(n577), .ZN(n407) );
  NOR2_X1 U472 ( .A1(n407), .A2(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(KEYINPUT47), .B(n408), .Z(n409) );
  NOR2_X1 U474 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n411), .B(KEYINPUT48), .ZN(n538) );
  XOR2_X1 U476 ( .A(G36GAT), .B(n412), .Z(n414) );
  NAND2_X1 U477 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n427) );
  XNOR2_X1 U479 ( .A(G211GAT), .B(G218GAT), .ZN(n416) );
  XOR2_X1 U480 ( .A(G197GAT), .B(G204GAT), .Z(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n442) );
  XOR2_X1 U482 ( .A(n419), .B(n442), .Z(n425) );
  XOR2_X1 U483 ( .A(KEYINPUT18), .B(KEYINPUT90), .Z(n421) );
  XNOR2_X1 U484 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U486 ( .A(KEYINPUT19), .B(n422), .Z(n461) );
  XNOR2_X1 U487 ( .A(n423), .B(n461), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U489 ( .A(n427), .B(n426), .Z(n473) );
  NOR2_X1 U490 ( .A1(n538), .A2(n473), .ZN(n428) );
  XOR2_X1 U491 ( .A(KEYINPUT54), .B(n428), .Z(n429) );
  XOR2_X1 U492 ( .A(KEYINPUT94), .B(KEYINPUT91), .Z(n431) );
  XNOR2_X1 U493 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U495 ( .A(n432), .B(KEYINPUT95), .Z(n435) );
  XNOR2_X1 U496 ( .A(G50GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U498 ( .A(KEYINPUT24), .B(n436), .Z(n438) );
  NAND2_X1 U499 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U501 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n482) );
  NAND2_X1 U504 ( .A1(n579), .A2(n482), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n446), .B(KEYINPUT120), .ZN(n464) );
  XOR2_X1 U507 ( .A(KEYINPUT20), .B(G99GAT), .Z(n448) );
  XNOR2_X1 U508 ( .A(G15GAT), .B(G190GAT), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U510 ( .A(n449), .B(G134GAT), .Z(n452) );
  XNOR2_X1 U511 ( .A(G43GAT), .B(n450), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(n457) );
  XOR2_X1 U513 ( .A(G169GAT), .B(n453), .Z(n455) );
  NAND2_X1 U514 ( .A1(G227GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U516 ( .A(n457), .B(n456), .Z(n463) );
  XOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT88), .Z(n459) );
  XNOR2_X1 U518 ( .A(KEYINPUT64), .B(KEYINPUT89), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n464), .A2(n537), .ZN(n568) );
  NOR2_X1 U522 ( .A1(n552), .A2(n568), .ZN(n467) );
  INV_X1 U523 ( .A(KEYINPUT58), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n569), .A2(n587), .ZN(n500) );
  INV_X1 U525 ( .A(n500), .ZN(n489) );
  INV_X1 U526 ( .A(n577), .ZN(n590) );
  NAND2_X1 U527 ( .A1(n590), .A2(n552), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT16), .ZN(n469) );
  XNOR2_X1 U529 ( .A(KEYINPUT87), .B(n469), .ZN(n488) );
  NOR2_X1 U530 ( .A1(n482), .A2(n537), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT26), .ZN(n580) );
  NAND2_X1 U532 ( .A1(n580), .A2(n481), .ZN(n557) );
  XNOR2_X1 U533 ( .A(n557), .B(KEYINPUT101), .ZN(n478) );
  INV_X1 U534 ( .A(n473), .ZN(n528) );
  NAND2_X1 U535 ( .A1(n528), .A2(n537), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n474), .A2(n482), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n475), .B(KEYINPUT102), .ZN(n476) );
  XNOR2_X1 U538 ( .A(KEYINPUT25), .B(n476), .ZN(n477) );
  XOR2_X1 U539 ( .A(KEYINPUT103), .B(n479), .Z(n480) );
  NOR2_X1 U540 ( .A1(n540), .A2(n480), .ZN(n486) );
  INV_X1 U541 ( .A(n481), .ZN(n483) );
  XOR2_X1 U542 ( .A(n482), .B(KEYINPUT28), .Z(n533) );
  NOR2_X1 U543 ( .A1(n483), .A2(n533), .ZN(n542) );
  NAND2_X1 U544 ( .A1(n542), .A2(n540), .ZN(n484) );
  NOR2_X1 U545 ( .A1(n537), .A2(n484), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT104), .B(n487), .Z(n498) );
  NAND2_X1 U547 ( .A1(n488), .A2(n498), .ZN(n513) );
  NOR2_X1 U548 ( .A1(n489), .A2(n513), .ZN(n495) );
  NAND2_X1 U549 ( .A1(n540), .A2(n495), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NAND2_X1 U552 ( .A1(n528), .A2(n495), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U555 ( .A1(n495), .A2(n537), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U557 ( .A1(n495), .A2(n533), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .Z(n503) );
  NOR2_X1 U560 ( .A1(n590), .A2(n597), .ZN(n497) );
  NAND2_X1 U561 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(KEYINPUT37), .B(n499), .ZN(n524) );
  NAND2_X1 U563 ( .A1(n500), .A2(n524), .ZN(n501) );
  XOR2_X1 U564 ( .A(KEYINPUT38), .B(n501), .Z(n508) );
  NAND2_X1 U565 ( .A1(n508), .A2(n540), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n508), .A2(n528), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n506) );
  NAND2_X1 U570 ( .A1(n537), .A2(n508), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U572 ( .A(G43GAT), .B(n507), .Z(G1330GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n510) );
  NAND2_X1 U574 ( .A1(n533), .A2(n508), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  NOR2_X1 U577 ( .A1(n582), .A2(n574), .ZN(n512) );
  XOR2_X1 U578 ( .A(KEYINPUT109), .B(n512), .Z(n525) );
  INV_X1 U579 ( .A(n525), .ZN(n514) );
  NAND2_X1 U580 ( .A1(n540), .A2(n521), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  NAND2_X1 U584 ( .A1(n528), .A2(n521), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n518), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U586 ( .A(G71GAT), .B(KEYINPUT111), .Z(n520) );
  NAND2_X1 U587 ( .A1(n521), .A2(n537), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U590 ( .A1(n521), .A2(n533), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U593 ( .A1(n532), .A2(n540), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n528), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U597 ( .A(G99GAT), .B(KEYINPUT113), .Z(n531) );
  NAND2_X1 U598 ( .A1(n537), .A2(n532), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1338GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U601 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U603 ( .A(n536), .B(G106GAT), .Z(G1339GAT) );
  INV_X1 U604 ( .A(n537), .ZN(n544) );
  INV_X1 U605 ( .A(n538), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n556) );
  INV_X1 U607 ( .A(n556), .ZN(n541) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n545), .A2(n553), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G113GAT), .B(n546), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U613 ( .A1(n553), .A2(n403), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n550) );
  NAND2_X1 U616 ( .A1(n553), .A2(n590), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(G127GAT), .B(n551), .Z(G1342GAT) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n406), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  XOR2_X1 U622 ( .A(G141GAT), .B(KEYINPUT117), .Z(n559) );
  NAND2_X1 U623 ( .A1(n566), .A2(n582), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1344GAT) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n561) );
  NAND2_X1 U627 ( .A1(n566), .A2(n403), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  XOR2_X1 U630 ( .A(G155GAT), .B(KEYINPUT119), .Z(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n590), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n406), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n573) );
  XNOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n574), .A2(n568), .ZN(n575) );
  XOR2_X1 U642 ( .A(n576), .B(n575), .Z(G1349GAT) );
  NOR2_X1 U643 ( .A1(n577), .A2(n568), .ZN(n578) );
  XOR2_X1 U644 ( .A(G183GAT), .B(n578), .Z(G1350GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT123), .ZN(n595) );
  NAND2_X1 U647 ( .A1(n595), .A2(n582), .ZN(n586) );
  XOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U652 ( .A(G204GAT), .B(KEYINPUT61), .Z(n589) );
  NAND2_X1 U653 ( .A1(n595), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1353GAT) );
  XOR2_X1 U655 ( .A(G211GAT), .B(KEYINPUT125), .Z(n592) );
  NAND2_X1 U656 ( .A1(n595), .A2(n590), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1354GAT) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n594) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n594), .B(n593), .ZN(n599) );
  INV_X1 U661 ( .A(n595), .ZN(n596) );
  NOR2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U663 ( .A(n599), .B(n598), .Z(G1355GAT) );
endmodule

