//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n208), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G155gat), .B(G162gat), .Z(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT2), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G141gat), .B(G148gat), .Z(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n218), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n214), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n213), .B1(new_n225), .B2(KEYINPUT29), .ZN(new_n226));
  AND2_X1   g025(.A1(G228gat), .A2(G233gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n222), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT3), .B1(new_n212), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n226), .B(new_n227), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n211), .A2(KEYINPUT83), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT29), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n210), .A2(KEYINPUT83), .A3(new_n211), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT3), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n226), .B1(new_n236), .B2(new_n229), .ZN(new_n237));
  INV_X1    g036(.A(new_n227), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n237), .A2(KEYINPUT84), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT84), .B1(new_n237), .B2(new_n238), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n232), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G22gat), .ZN(new_n242));
  INV_X1    g041(.A(G78gat), .ZN(new_n243));
  INV_X1    g042(.A(G22gat), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(new_n232), .C1(new_n239), .C2(new_n240), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n243), .B1(new_n242), .B2(new_n245), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT31), .B(G50gat), .ZN(new_n248));
  INV_X1    g047(.A(G106gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n246), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n242), .A2(new_n245), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G78gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(G64gat), .B(G92gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT27), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n264), .B2(G183gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT27), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(KEYINPUT69), .A2(KEYINPUT27), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(G183gat), .B1(KEYINPUT69), .B2(KEYINPUT27), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n263), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n277));
  AOI21_X1  g076(.A(G190gat), .B1(new_n277), .B2(KEYINPUT68), .ZN(new_n278));
  OR2_X1    g077(.A1(KEYINPUT69), .A2(KEYINPUT27), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(G183gat), .A3(new_n271), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT70), .A4(new_n268), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n275), .A2(new_n281), .A3(new_n284), .A4(new_n276), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n264), .A2(G183gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n277), .A2(new_n286), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n287), .A2(new_n276), .A3(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT64), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n291), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(KEYINPUT26), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n296), .A2(new_n300), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT25), .ZN(new_n305));
  NAND2_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n306));
  MUX2_X1   g105(.A(G183gat), .B(new_n306), .S(G190gat), .Z(new_n307));
  AOI21_X1  g106(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n308), .A2(KEYINPUT66), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(KEYINPUT66), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT67), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n308), .B(KEYINPUT66), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(new_n307), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n305), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n297), .B1(new_n295), .B2(new_n303), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT65), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n319), .B(new_n297), .C1(new_n295), .C2(new_n303), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n304), .A2(new_n323), .A3(new_n297), .ZN(new_n324));
  INV_X1    g123(.A(new_n308), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT25), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n302), .A2(KEYINPUT76), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n331));
  INV_X1    g130(.A(new_n301), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n288), .B1(new_n282), .B2(KEYINPUT71), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n285), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n327), .B1(new_n316), .B2(new_n321), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n330), .A2(new_n336), .A3(new_n230), .ZN(new_n337));
  NAND2_X1  g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT75), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n334), .A2(new_n335), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(new_n338), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n213), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n336), .A3(new_n339), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n338), .B1(new_n342), .B2(KEYINPUT29), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n212), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n343), .B1(new_n337), .B2(new_n340), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT77), .B(new_n350), .C1(new_n351), .C2(new_n212), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n262), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(G113gat), .B(G120gat), .Z(new_n354));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n228), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT72), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n359), .A2(KEYINPUT72), .A3(new_n360), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n229), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n364), .B1(new_n370), .B2(new_n363), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n361), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n359), .A2(KEYINPUT81), .A3(new_n360), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n224), .ZN(new_n377));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n371), .A2(new_n372), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n363), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n366), .A2(new_n229), .A3(KEYINPUT4), .A4(new_n367), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n382), .A2(new_n377), .A3(new_n383), .A4(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n375), .A2(new_n228), .A3(new_n376), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n362), .ZN(new_n387));
  INV_X1    g186(.A(new_n378), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n387), .A2(KEYINPUT82), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT82), .B1(new_n387), .B2(new_n388), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n385), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT0), .ZN(new_n393));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OR3_X1    g195(.A1(new_n381), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n381), .B2(new_n391), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT6), .B(new_n396), .C1(new_n381), .C2(new_n391), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT37), .B1(new_n347), .B2(new_n352), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(new_n261), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT37), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n348), .A2(new_n213), .A3(new_n349), .ZN(new_n406));
  AOI211_X1 g205(.A(new_n405), .B(new_n406), .C1(new_n212), .C2(new_n345), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT38), .ZN(new_n408));
  AOI211_X1 g207(.A(new_n353), .B(new_n402), .C1(new_n404), .C2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n404), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n212), .B1(new_n341), .B2(new_n344), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n351), .A2(KEYINPUT77), .A3(new_n212), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT78), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT78), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n347), .A2(new_n352), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n405), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT38), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n258), .B1(new_n409), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n353), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n421), .A2(new_n422), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n353), .A2(KEYINPUT80), .A3(KEYINPUT30), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n417), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n416), .B1(new_n347), .B2(new_n352), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n262), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT79), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n417), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT79), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n262), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n429), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n371), .A2(new_n377), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n388), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(KEYINPUT39), .C1(new_n388), .C2(new_n387), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(new_n395), .C1(KEYINPUT39), .C2(new_n439), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT40), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n442), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n399), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n420), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n342), .A2(new_n368), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n369), .B1(new_n334), .B2(new_n335), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT34), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI211_X1 g252(.A(KEYINPUT34), .B(new_n447), .C1(new_n448), .C2(new_n449), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(KEYINPUT73), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT73), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n452), .B2(new_n454), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n448), .A2(new_n447), .A3(new_n449), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460));
  XOR2_X1   g259(.A(G15gat), .B(G43gat), .Z(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n459), .B(KEYINPUT32), .C1(new_n460), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n459), .A2(KEYINPUT32), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n460), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n463), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n456), .A2(new_n458), .A3(new_n465), .A4(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n452), .A2(new_n454), .ZN(new_n470));
  INV_X1    g269(.A(new_n468), .ZN(new_n471));
  INV_X1    g270(.A(new_n465), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT73), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n257), .A2(KEYINPUT85), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n252), .B2(new_n256), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n347), .A2(new_n352), .ZN(new_n481));
  AND4_X1   g280(.A1(KEYINPUT80), .A2(new_n481), .A3(KEYINPUT30), .A4(new_n261), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n425), .B1(new_n353), .B2(new_n423), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n435), .B1(new_n434), .B2(new_n262), .ZN(new_n485));
  AOI211_X1 g284(.A(KEYINPUT79), .B(new_n261), .C1(new_n415), .C2(new_n417), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n402), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n476), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n446), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n257), .A2(new_n474), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT35), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n251), .B1(new_n246), .B2(new_n247), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n254), .A2(new_n255), .A3(new_n250), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT86), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT86), .B1(new_n469), .B2(new_n473), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n437), .A2(new_n498), .A3(new_n402), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(KEYINPUT88), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n502), .B2(KEYINPUT88), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G43gat), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(G50gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT89), .B(G50gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(G43gat), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n510), .A2(new_n504), .ZN(new_n511));
  INV_X1    g310(.A(G29gat), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n512), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT14), .B(G29gat), .ZN(new_n514));
  INV_X1    g313(.A(G36gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n506), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n506), .B2(new_n516), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(G1gat), .B2(new_n519), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(G8gat), .Z(new_n523));
  NOR2_X1   g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n518), .A2(KEYINPUT17), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n518), .A2(KEYINPUT17), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n528), .A2(new_n523), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n524), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(KEYINPUT18), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n518), .B(new_n523), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n531), .B(KEYINPUT13), .Z(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(KEYINPUT91), .A3(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G113gat), .B(G141gat), .Z(new_n537));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  XOR2_X1   g340(.A(new_n541), .B(KEYINPUT12), .Z(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n532), .A2(new_n535), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT18), .B1(new_n530), .B2(new_n531), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n536), .B(new_n543), .C1(new_n545), .C2(new_n546), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n501), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n554), .B2(new_n553), .ZN(new_n556));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT93), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n553), .B(KEYINPUT94), .ZN(new_n560));
  INV_X1    g359(.A(G71gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n243), .A3(KEYINPUT9), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n561), .B2(new_n243), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT95), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT96), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n570), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n523), .B1(new_n566), .B2(new_n567), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT7), .ZN(new_n584));
  INV_X1    g383(.A(G99gat), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT8), .B1(new_n585), .B2(new_n249), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n584), .B(new_n586), .C1(G85gat), .C2(G92gat), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n582), .B1(new_n518), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n518), .B2(KEYINPUT17), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n527), .B2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G190gat), .B(G218gat), .Z(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT97), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n593), .A2(new_n594), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n595), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n588), .A2(KEYINPUT98), .ZN(new_n607));
  OR3_X1    g406(.A1(new_n566), .A2(new_n589), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n589), .B1(new_n566), .B2(new_n607), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n559), .A2(new_n565), .A3(KEYINPUT10), .A4(new_n591), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT99), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT101), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(new_n618), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n615), .B1(new_n608), .B2(new_n610), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT100), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n622), .A2(new_n616), .A3(new_n626), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n581), .A2(new_n606), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n551), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n402), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g435(.A1(new_n551), .A2(new_n437), .ZN(new_n637));
  INV_X1    g436(.A(new_n632), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n639), .A2(G8gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT16), .B(G8gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT42), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(KEYINPUT42), .B2(new_n642), .ZN(G1325gat));
  NOR2_X1   g443(.A1(new_n496), .A2(new_n497), .ZN(new_n645));
  AOI21_X1  g444(.A(G15gat), .B1(new_n633), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT102), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n476), .A2(G15gat), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n633), .B2(new_n648), .ZN(G1326gat));
  INV_X1    g448(.A(new_n480), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n551), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n638), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT103), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT43), .B(G22gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  AND3_X1   g454(.A1(new_n491), .A2(new_n499), .A3(KEYINPUT104), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT104), .B1(new_n491), .B2(new_n499), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n489), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n658), .B2(new_n605), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660));
  AOI211_X1 g459(.A(new_n660), .B(new_n606), .C1(new_n489), .C2(new_n500), .ZN(new_n661));
  INV_X1    g460(.A(new_n550), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n581), .A2(new_n662), .A3(new_n630), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n659), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G29gat), .B1(new_n666), .B2(new_n402), .ZN(new_n667));
  INV_X1    g466(.A(new_n551), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n581), .A2(new_n606), .A3(new_n630), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n668), .A2(new_n512), .A3(new_n634), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n637), .A2(new_n515), .A3(new_n669), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT46), .Z(new_n674));
  OAI21_X1  g473(.A(G36gat), .B1(new_n666), .B2(new_n437), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(G1329gat));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n665), .A2(new_n476), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n669), .A2(new_n507), .A3(new_n645), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n679), .A2(G43gat), .B1(new_n668), .B2(new_n680), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n677), .B(new_n678), .C1(new_n681), .C2(KEYINPUT105), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT47), .B1(new_n681), .B2(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n680), .ZN(new_n684));
  INV_X1    g483(.A(new_n476), .ZN(new_n685));
  NOR4_X1   g484(.A1(new_n659), .A2(new_n661), .A3(new_n685), .A4(new_n664), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n686), .B2(new_n507), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT106), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n682), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(G1330gat));
  NAND3_X1  g490(.A1(new_n651), .A2(new_n509), .A3(new_n669), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n666), .A2(new_n257), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT48), .B(new_n692), .C1(new_n693), .C2(new_n509), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n509), .B1(new_n665), .B2(new_n480), .ZN(new_n695));
  INV_X1    g494(.A(new_n692), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(KEYINPUT48), .B2(new_n697), .ZN(G1331gat));
  INV_X1    g497(.A(new_n581), .ZN(new_n699));
  NOR4_X1   g498(.A1(new_n699), .A2(new_n550), .A3(new_n605), .A4(new_n631), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n658), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n634), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G57gat), .ZN(G1332gat));
  INV_X1    g502(.A(new_n437), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT49), .B(G64gat), .Z(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n705), .B2(new_n707), .ZN(G1333gat));
  NAND3_X1  g507(.A1(new_n701), .A2(G71gat), .A3(new_n476), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT107), .ZN(new_n710));
  INV_X1    g509(.A(new_n701), .ZN(new_n711));
  INV_X1    g510(.A(new_n645), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n561), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n701), .A2(new_n480), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g516(.A1(new_n659), .A2(new_n661), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n581), .A2(new_n550), .A3(new_n631), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721), .B2(new_n402), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n500), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n491), .A2(new_n499), .A3(KEYINPUT104), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n606), .B1(new_n726), .B2(new_n489), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n581), .A2(new_n550), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT51), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n658), .A2(KEYINPUT51), .A3(new_n605), .A4(new_n728), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n630), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n402), .A2(G85gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n722), .B1(new_n732), .B2(new_n733), .ZN(G1336gat));
  AOI22_X1  g533(.A1(new_n724), .A2(new_n725), .B1(new_n446), .B2(new_n488), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n660), .B1(new_n735), .B2(new_n606), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n501), .A2(KEYINPUT44), .A3(new_n605), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n736), .A2(new_n704), .A3(new_n737), .A4(new_n719), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G92gat), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n437), .A2(new_n631), .A3(G92gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n729), .B2(new_n731), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744));
  INV_X1    g543(.A(new_n740), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n658), .A2(new_n605), .A3(new_n728), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n748), .B2(new_n730), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n739), .B1(KEYINPUT108), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n744), .B(KEYINPUT52), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n741), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n756), .A3(new_n739), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n744), .B1(new_n757), .B2(KEYINPUT52), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n743), .B1(new_n753), .B2(new_n758), .ZN(G1337gat));
  NAND2_X1  g558(.A1(new_n720), .A2(new_n476), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n585), .B1(new_n760), .B2(KEYINPUT110), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(KEYINPUT110), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n645), .A2(new_n585), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n732), .B2(new_n763), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n718), .A2(new_n480), .A3(new_n719), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n765), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT111), .B1(new_n765), .B2(G106gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n729), .A2(new_n731), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n258), .A2(new_n249), .A3(new_n630), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT112), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n766), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n249), .B1(new_n720), .B2(new_n258), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n768), .B2(new_n769), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(G1339gat));
  NOR2_X1   g575(.A1(new_n632), .A2(new_n550), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n617), .A2(new_n778), .A3(new_n619), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n614), .B2(new_n615), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n611), .A2(G230gat), .A3(G233gat), .A4(new_n613), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n626), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(new_n629), .ZN(new_n784));
  INV_X1    g583(.A(new_n541), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n530), .A2(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n547), .A2(new_n542), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n779), .A2(new_n782), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n784), .A2(new_n605), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n788), .A2(new_n789), .B1(new_n548), .B2(new_n549), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n792), .A2(new_n784), .B1(new_n630), .B2(new_n787), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n793), .B2(new_n605), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n581), .B1(new_n794), .B2(KEYINPUT113), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n777), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n480), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT114), .B1(new_n797), .B2(new_n480), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n437), .A2(new_n634), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n712), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n550), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G113gat), .ZN(new_n804));
  NOR4_X1   g603(.A1(new_n797), .A2(new_n402), .A3(new_n704), .A4(new_n490), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n662), .A2(G113gat), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT115), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(new_n810), .A3(new_n630), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n800), .A2(new_n630), .A3(new_n802), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n812), .A2(new_n813), .A3(G120gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n812), .B2(G120gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n805), .A2(new_n817), .A3(new_n581), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n581), .A3(new_n802), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n817), .ZN(G1342gat));
  INV_X1    g620(.A(G134gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n822), .A3(new_n605), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT56), .Z(new_n824));
  NAND3_X1  g623(.A1(new_n800), .A2(new_n605), .A3(new_n802), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n825), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT117), .B1(new_n825), .B2(G134gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(G1343gat));
  NAND2_X1  g627(.A1(new_n795), .A2(new_n796), .ZN(new_n829));
  INV_X1    g628(.A(new_n777), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n634), .ZN(new_n832));
  NOR4_X1   g631(.A1(new_n832), .A2(new_n704), .A3(new_n257), .A4(new_n476), .ZN(new_n833));
  INV_X1    g632(.A(G141gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n550), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n836), .A3(new_n258), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n605), .B1(new_n793), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n784), .A2(new_n792), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n630), .A2(new_n787), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT118), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n581), .B1(new_n843), .B2(new_n791), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n480), .B1(new_n844), .B2(new_n777), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n801), .A2(new_n476), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n837), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G141gat), .B1(new_n848), .B2(new_n662), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n835), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g650(.A(G148gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n833), .A2(new_n852), .A3(new_n630), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(KEYINPUT59), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n848), .B2(new_n631), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n844), .B2(new_n777), .ZN(new_n860));
  INV_X1    g659(.A(new_n791), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n839), .B2(new_n842), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT120), .B(new_n830), .C1(new_n862), .C2(new_n581), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n650), .A2(KEYINPUT57), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT57), .B1(new_n797), .B2(new_n257), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n865), .A2(new_n630), .A3(new_n847), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n858), .B1(new_n867), .B2(G148gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n853), .B1(new_n857), .B2(new_n868), .ZN(G1345gat));
  NAND3_X1  g668(.A1(new_n833), .A2(new_n216), .A3(new_n581), .ZN(new_n870));
  OAI21_X1  g669(.A(G155gat), .B1(new_n848), .B2(new_n699), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1346gat));
  NAND3_X1  g671(.A1(new_n833), .A2(new_n217), .A3(new_n605), .ZN(new_n873));
  OAI21_X1  g672(.A(G162gat), .B1(new_n848), .B2(new_n606), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT121), .ZN(G1347gat));
  NOR4_X1   g675(.A1(new_n797), .A2(new_n634), .A3(new_n437), .A4(new_n490), .ZN(new_n877));
  AOI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n550), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n437), .A2(new_n634), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n645), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT122), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n798), .B2(new_n799), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n550), .A2(G169gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(G1348gat));
  NAND3_X1  g683(.A1(new_n882), .A2(G176gat), .A3(new_n630), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(KEYINPUT123), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(KEYINPUT123), .ZN(new_n887));
  AOI21_X1  g686(.A(G176gat), .B1(new_n877), .B2(new_n630), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G1349gat));
  AOI21_X1  g688(.A(new_n267), .B1(new_n882), .B2(new_n581), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n877), .A2(new_n277), .A3(new_n286), .A4(new_n581), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT124), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n890), .A2(KEYINPUT60), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT60), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1350gat));
  AOI21_X1  g694(.A(new_n269), .B1(new_n882), .B2(new_n605), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT61), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n877), .A2(new_n269), .A3(new_n605), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT125), .Z(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(KEYINPUT61), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(G1351gat));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n685), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT126), .Z(new_n903));
  NAND3_X1  g702(.A1(new_n865), .A2(new_n866), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(G197gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(new_n662), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n685), .A2(new_n704), .A3(new_n258), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n634), .B(new_n907), .C1(new_n829), .C2(new_n830), .ZN(new_n908));
  AOI21_X1  g707(.A(G197gat), .B1(new_n908), .B2(new_n550), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n906), .A2(new_n909), .ZN(G1352gat));
  INV_X1    g709(.A(G204gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n911), .A3(new_n630), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT62), .Z(new_n913));
  OAI21_X1  g712(.A(G204gat), .B1(new_n904), .B2(new_n631), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1353gat));
  NAND3_X1  g714(.A1(new_n908), .A2(new_n203), .A3(new_n581), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n865), .A2(new_n866), .A3(new_n581), .A4(new_n903), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n917), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT63), .B1(new_n917), .B2(G211gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n916), .B(new_n922), .C1(new_n918), .C2(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1354gat));
  OAI21_X1  g723(.A(G218gat), .B1(new_n904), .B2(new_n606), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n204), .A3(new_n605), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1355gat));
endmodule


