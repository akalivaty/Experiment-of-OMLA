//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982;
  OAI21_X1  g000(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(KEYINPUT83), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(KEYINPUT83), .B2(new_n207), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(new_n205), .B2(new_n206), .ZN(new_n210));
  AND2_X1   g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT15), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT84), .B(G43gat), .Z(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  AOI211_X1 g016(.A(KEYINPUT15), .B(new_n211), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT85), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n207), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n204), .A2(new_n205), .A3(new_n206), .A4(KEYINPUT85), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n203), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n213), .B1(new_n205), .B2(new_n206), .ZN(new_n223));
  OR3_X1    g022(.A1(new_n218), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n215), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n226), .A2(G1gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228));
  AOI21_X1  g027(.A(G8gat), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n230), .B2(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n229), .B(new_n232), .ZN(new_n233));
  OR3_X1    g032(.A1(new_n225), .A2(KEYINPUT88), .A3(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT88), .B1(new_n225), .B2(new_n233), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n224), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT17), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n233), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT89), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G197gat), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT11), .B(G169gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n249), .B(KEYINPUT12), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n233), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n242), .B(KEYINPUT13), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(new_n244), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n236), .A2(new_n241), .A3(KEYINPUT18), .A4(new_n242), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n254), .A2(new_n255), .B1(new_n243), .B2(new_n244), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n261), .B(new_n258), .C1(new_n245), .C2(new_n251), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g062(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n265));
  AND2_X1   g064(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n268), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n264), .A2(new_n270), .A3(new_n265), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT27), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G183gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n277), .B2(new_n267), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT26), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(KEYINPUT26), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(new_n279), .A3(KEYINPUT26), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n269), .A2(new_n278), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  AND2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n292), .B1(KEYINPUT23), .B2(new_n282), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT65), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n282), .A2(new_n296), .A3(KEYINPUT23), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT24), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(G190gat), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n300), .A2(new_n302), .B1(new_n273), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n291), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n264), .A2(new_n274), .A3(new_n276), .A4(new_n265), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n300), .A2(new_n302), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n296), .B1(new_n282), .B2(KEYINPUT23), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n294), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n291), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT23), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n288), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT66), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n309), .A2(new_n312), .A3(new_n314), .A4(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n305), .A2(new_n306), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n306), .B1(new_n305), .B2(new_n318), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n290), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G127gat), .B(G134gat), .Z(new_n322));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(KEYINPUT1), .B2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G113gat), .B(G120gat), .Z(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  XNOR2_X1  g125(.A(G127gat), .B(G134gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  AND4_X1   g129(.A1(new_n312), .A2(new_n309), .A3(new_n314), .A4(new_n317), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n316), .B1(new_n310), .B2(new_n311), .ZN(new_n332));
  INV_X1    g131(.A(new_n304), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT25), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT69), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n305), .A2(new_n318), .A3(new_n306), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n324), .A2(new_n328), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n290), .ZN(new_n339));
  NAND2_X1  g138(.A1(G227gat), .A2(G233gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n340), .B(KEYINPUT64), .Z(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n330), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT34), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT34), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n330), .A2(new_n339), .A3(new_n345), .A4(new_n342), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(G15gat), .B(G43gat), .Z(new_n348));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n338), .B1(new_n337), .B2(new_n290), .ZN(new_n352));
  INV_X1    g151(.A(new_n290), .ZN(new_n353));
  AOI211_X1 g152(.A(new_n329), .B(new_n353), .C1(new_n335), .C2(new_n336), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n341), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT33), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n342), .B1(new_n330), .B2(new_n339), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n350), .B1(new_n359), .B2(KEYINPUT33), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n344), .A3(new_n346), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(KEYINPUT32), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(new_n217), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT2), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT73), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n372), .A3(KEYINPUT2), .ZN(new_n373));
  AND2_X1   g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n378), .B2(new_n379), .ZN(new_n383));
  INV_X1    g182(.A(G155gat), .ZN(new_n384));
  INV_X1    g183(.A(G162gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(KEYINPUT74), .A3(new_n369), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n383), .A2(new_n387), .A3(new_n370), .A4(new_n376), .ZN(new_n388));
  XOR2_X1   g187(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(G211gat), .A2(G218gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(G211gat), .A2(G218gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(G197gat), .A2(G204gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(G197gat), .A2(G204gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G211gat), .B(G218gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(G197gat), .B(G204gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n399), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n392), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n389), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n405), .B2(new_n391), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n387), .A2(new_n370), .A3(new_n376), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n410), .A2(new_n383), .B1(new_n377), .B2(new_n380), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT79), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n373), .ZN(new_n413));
  XNOR2_X1  g212(.A(G141gat), .B(G148gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n372), .B1(new_n369), .B2(KEYINPUT2), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n380), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n388), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT29), .B1(new_n400), .B2(new_n404), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n418), .B(new_n419), .C1(new_n408), .C2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n407), .A2(new_n412), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n392), .B2(new_n406), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n414), .A2(new_n415), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n417), .B1(new_n427), .B2(new_n373), .ZN(new_n428));
  AND4_X1   g227(.A1(new_n370), .A2(new_n383), .A3(new_n387), .A4(new_n376), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n388), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n430), .B(new_n431), .C1(KEYINPUT3), .C2(new_n420), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n368), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(G22gat), .B1(new_n434), .B2(KEYINPUT80), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n422), .A2(new_n423), .B1(new_n432), .B2(new_n425), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n436), .A2(new_n368), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n438));
  INV_X1    g237(.A(G22gat), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n438), .B(new_n439), .C1(new_n436), .C2(new_n368), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n435), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n435), .B2(new_n440), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n363), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n358), .A2(new_n361), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n364), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G8gat), .B(G36gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(G64gat), .B(G92gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT71), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n353), .B1(new_n335), .B2(new_n336), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(KEYINPUT29), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n269), .A2(new_n278), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n456), .A2(new_n289), .B1(new_n305), .B2(new_n318), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(new_n451), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n405), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n451), .B1(new_n457), .B2(KEYINPUT29), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(new_n405), .C1(new_n454), .C2(new_n453), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n450), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT72), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n452), .B1(new_n321), .B2(new_n391), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n406), .B1(new_n466), .B2(new_n458), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT72), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n450), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n462), .A3(new_n449), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT30), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT30), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n467), .A2(new_n473), .A3(new_n462), .A4(new_n449), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n465), .A2(new_n470), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT4), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n418), .B2(new_n329), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n381), .A4(new_n388), .ZN(new_n478));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n430), .A2(KEYINPUT3), .A3(new_n431), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n338), .B1(new_n411), .B2(new_n389), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n479), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n388), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT75), .B1(new_n381), .B2(new_n388), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n486), .A2(new_n487), .A3(new_n338), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n418), .A2(new_n329), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(KEYINPUT5), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n485), .A2(KEYINPUT5), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT77), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT77), .B1(new_n477), .B2(new_n478), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n483), .B(new_n492), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G1gat), .B(G29gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT0), .ZN(new_n499));
  XNOR2_X1  g298(.A(G57gat), .B(G85gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n499), .B(new_n500), .Z(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g301(.A(new_n501), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n497), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n491), .A2(new_n496), .A3(new_n504), .A4(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n475), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT35), .B1(new_n446), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n358), .A2(new_n361), .A3(new_n444), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n444), .B1(new_n358), .B2(new_n361), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n465), .A2(new_n470), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n472), .A2(new_n474), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n514), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n513), .A2(new_n516), .A3(new_n517), .A4(new_n443), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n511), .B2(new_n512), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n364), .A2(KEYINPUT36), .A3(new_n445), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n506), .A2(new_n507), .A3(new_n471), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT37), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n290), .B1(new_n331), .B2(new_n334), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n391), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n321), .A2(new_n452), .B1(new_n528), .B2(new_n451), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n529), .B2(new_n406), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n405), .B1(new_n466), .B2(new_n458), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n449), .B1(new_n467), .B2(new_n462), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n449), .A2(new_n526), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n525), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n534), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n464), .A2(new_n536), .B1(new_n468), .B2(KEYINPUT37), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n524), .B(new_n535), .C1(new_n537), .C2(new_n525), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT40), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n477), .A2(new_n478), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT77), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n493), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n479), .B1(new_n543), .B2(new_n483), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT39), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n501), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n430), .A2(new_n329), .A3(new_n431), .ZN(new_n548));
  INV_X1    g347(.A(new_n489), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(new_n479), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT39), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(KEYINPUT81), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT81), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n553), .B1(new_n550), .B2(KEYINPUT39), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n544), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n539), .B1(new_n547), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n503), .B1(new_n544), .B2(new_n545), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n544), .A2(new_n554), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT40), .B(new_n557), .C1(new_n558), .C2(new_n552), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n497), .A2(new_n503), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n538), .B(new_n443), .C1(new_n475), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n443), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n509), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n523), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n263), .B1(new_n519), .B2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G57gat), .B(G64gat), .Z(new_n567));
  INV_X1    g366(.A(KEYINPUT9), .ZN(new_n568));
  INV_X1    g367(.A(G71gat), .ZN(new_n569));
  INV_X1    g368(.A(G78gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n567), .B1(KEYINPUT90), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n571), .A2(KEYINPUT90), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G71gat), .B(G78gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G127gat), .B(G155gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT91), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n580), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G183gat), .B(G211gat), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n233), .B1(new_n576), .B2(new_n577), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT93), .B(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT8), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT94), .ZN(new_n605));
  XOR2_X1   g404(.A(G99gat), .B(G106gat), .Z(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  OR3_X1    g406(.A1(new_n607), .A2(new_n600), .A3(KEYINPUT7), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT7), .B1(new_n607), .B2(new_n600), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT95), .A2(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n606), .A2(KEYINPUT95), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n605), .B(new_n610), .C1(KEYINPUT95), .C2(new_n606), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT96), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n617), .A3(new_n614), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n238), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n615), .A2(new_n237), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(KEYINPUT97), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n598), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  AOI211_X1 g425(.A(new_n624), .B(new_n597), .C1(new_n619), .C2(new_n621), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT92), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(KEYINPUT97), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n626), .B2(new_n627), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n596), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(G230gat), .ZN(new_n639));
  INV_X1    g438(.A(G233gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n576), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n615), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n613), .A2(new_n576), .A3(new_n614), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n642), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n641), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n643), .A2(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n641), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n649), .A2(new_n651), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n638), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n566), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n508), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n663), .A2(new_n475), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G8gat), .B1(new_n663), .B2(new_n475), .ZN(new_n672));
  NOR2_X1   g471(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n673));
  MUX2_X1   g472(.A(KEYINPUT100), .B(new_n673), .S(new_n670), .Z(new_n674));
  AOI22_X1  g473(.A1(new_n671), .A2(new_n672), .B1(new_n669), .B2(new_n674), .ZN(G1325gat));
  AOI21_X1  g474(.A(G15gat), .B1(new_n664), .B2(new_n513), .ZN(new_n676));
  INV_X1    g475(.A(new_n523), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT101), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(new_n664), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n443), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NOR3_X1   g482(.A1(new_n596), .A2(new_n637), .A3(new_n661), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n566), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(G29gat), .A3(new_n508), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n596), .A2(new_n263), .A3(new_n661), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n519), .A2(new_n565), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(new_n636), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n633), .A2(KEYINPUT104), .A3(new_n635), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT104), .B1(new_n633), .B2(new_n635), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n692), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n565), .B2(new_n519), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n691), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT105), .B(new_n691), .C1(new_n694), .C2(new_n699), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n704), .A2(new_n665), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n690), .B1(new_n705), .B2(new_n205), .ZN(G1328gat));
  NOR3_X1   g505(.A1(new_n687), .A2(G36gat), .A3(new_n475), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT46), .ZN(new_n708));
  INV_X1    g507(.A(new_n475), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT106), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G36gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n710), .A2(KEYINPUT106), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n708), .B1(new_n712), .B2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(new_n216), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n700), .B2(new_n523), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n686), .A2(new_n216), .A3(new_n513), .A4(new_n566), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(KEYINPUT47), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n677), .A3(new_n703), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(new_n715), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(KEYINPUT108), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI211_X1 g522(.A(KEYINPUT108), .B(new_n216), .C1(new_n704), .C2(new_n677), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n718), .B1(new_n723), .B2(new_n724), .ZN(G1330gat));
  OAI21_X1  g524(.A(G50gat), .B1(new_n700), .B2(new_n443), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n217), .B(new_n563), .C1(new_n687), .C2(KEYINPUT110), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n687), .A2(KEYINPUT110), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT48), .B(new_n726), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n702), .A2(new_n563), .A3(new_n703), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n730), .A2(new_n731), .A3(G50gat), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n730), .B2(G50gat), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n727), .A2(new_n728), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n729), .B1(new_n735), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g535(.A1(new_n260), .A2(new_n262), .ZN(new_n737));
  INV_X1    g536(.A(new_n661), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n638), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n693), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n665), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n709), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT49), .B(G64gat), .Z(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(G1333gat));
  AOI21_X1  g545(.A(new_n569), .B1(new_n740), .B2(new_n677), .ZN(new_n747));
  INV_X1    g546(.A(new_n513), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(G71gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n740), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n563), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT112), .B(G78gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n694), .A2(new_n699), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n595), .A2(new_n263), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n756), .A2(new_n738), .A3(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(new_n665), .ZN(new_n759));
  AOI211_X1 g558(.A(new_n637), .B(new_n757), .C1(new_n519), .C2(new_n565), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(KEYINPUT51), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(KEYINPUT51), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n661), .A2(new_n665), .A3(new_n599), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n759), .A2(new_n599), .B1(new_n763), .B2(new_n764), .ZN(G1336gat));
  NAND2_X1  g564(.A1(new_n661), .A2(new_n600), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n763), .A2(new_n475), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n600), .B1(new_n758), .B2(new_n709), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1337gat));
  AND2_X1   g570(.A1(new_n758), .A2(new_n677), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(G99gat), .A3(new_n774), .ZN(new_n775));
  OR4_X1    g574(.A1(G99gat), .A2(new_n763), .A3(new_n748), .A4(new_n738), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1338gat));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n563), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G106gat), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n738), .A2(G106gat), .A3(new_n443), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT114), .Z(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n761), .B2(new_n762), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT53), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  INV_X1    g587(.A(new_n780), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n779), .B(new_n788), .C1(new_n763), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1339gat));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n636), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n695), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n646), .A2(new_n647), .A3(new_n641), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n649), .A2(KEYINPUT54), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n659), .B1(new_n648), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n660), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  INV_X1    g601(.A(new_n795), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n803), .A2(new_n648), .A3(new_n797), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n648), .A2(new_n797), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n657), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n802), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n796), .A2(new_n798), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(KEYINPUT116), .A3(new_n802), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n801), .A2(new_n809), .A3(new_n737), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n254), .A2(new_n255), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n242), .B1(new_n236), .B2(new_n241), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n249), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n261), .A2(new_n251), .A3(new_n258), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n661), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n794), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n696), .A2(new_n697), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n816), .A2(new_n815), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n801), .A2(new_n809), .A3(new_n821), .A4(new_n811), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n595), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n638), .A2(new_n737), .A3(new_n661), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n563), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n475), .A2(new_n665), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n748), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(G113gat), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n830), .A2(new_n831), .A3(new_n263), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n508), .B1(new_n824), .B2(new_n826), .ZN(new_n833));
  INV_X1    g632(.A(new_n446), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n833), .A2(new_n475), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n737), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n832), .B1(new_n836), .B2(new_n831), .ZN(G1340gat));
  INV_X1    g636(.A(G120gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n838), .A3(new_n661), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n827), .A2(new_n661), .A3(new_n829), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n840), .A2(KEYINPUT117), .A3(G120gat), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT117), .B1(new_n840), .B2(G120gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n835), .A2(new_n844), .A3(new_n596), .ZN(new_n845));
  OAI21_X1  g644(.A(G127gat), .B1(new_n830), .B2(new_n595), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  INV_X1    g646(.A(G134gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n637), .A2(new_n709), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n848), .A3(new_n834), .A4(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n830), .B2(new_n637), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NOR2_X1   g653(.A1(new_n677), .A2(new_n828), .ZN(new_n855));
  INV_X1    g654(.A(G141gat), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n263), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n824), .A2(new_n826), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n858), .B2(new_n563), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n443), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT55), .B1(new_n810), .B2(KEYINPUT118), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(KEYINPUT118), .B2(new_n810), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n737), .A3(new_n801), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n636), .B1(new_n865), .B2(new_n818), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n595), .B1(new_n866), .B2(new_n823), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n862), .B1(new_n867), .B2(new_n826), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n855), .B(new_n857), .C1(new_n859), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n677), .A2(new_n443), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n833), .A2(new_n737), .A3(new_n475), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n856), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT58), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n873), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1344gat));
  AND2_X1   g678(.A1(new_n833), .A2(new_n870), .ZN(new_n880));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n475), .A4(new_n661), .ZN(new_n882));
  XNOR2_X1  g681(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n800), .B1(new_n808), .B2(new_n807), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n636), .A3(new_n821), .A4(new_n811), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n263), .A2(new_n800), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n817), .B1(new_n886), .B2(new_n864), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(new_n636), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n825), .B1(new_n888), .B2(new_n595), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n860), .B1(new_n889), .B2(new_n443), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n858), .A2(new_n861), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n661), .A3(new_n855), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n883), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n881), .A2(KEYINPUT59), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n855), .B1(new_n859), .B2(new_n868), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n661), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n882), .B1(new_n894), .B2(new_n898), .ZN(G1345gat));
  NAND2_X1  g698(.A1(new_n596), .A2(G155gat), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT121), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n475), .A3(new_n596), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n897), .A2(new_n901), .B1(new_n902), .B2(new_n384), .ZN(G1346gat));
  NAND3_X1  g702(.A1(new_n880), .A2(new_n385), .A3(new_n849), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT122), .B1(new_n896), .B2(new_n820), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G162gat), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n896), .A2(KEYINPUT122), .A3(new_n820), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n475), .A2(new_n665), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n748), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n827), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n284), .A3(new_n263), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n665), .B1(new_n824), .B2(new_n826), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n446), .A2(new_n475), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n737), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n913), .B1(new_n284), .B2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n912), .B2(new_n738), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n661), .A2(new_n285), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1349gat));
  OAI211_X1 g723(.A(new_n917), .B(new_n596), .C1(new_n267), .C2(new_n266), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n274), .A2(new_n276), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n912), .B2(new_n595), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n925), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1350gat));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n264), .A3(new_n265), .A4(new_n794), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n303), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n912), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n636), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n933), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  INV_X1    g741(.A(G197gat), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n677), .A2(new_n910), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n890), .B2(new_n891), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n943), .B1(new_n946), .B2(new_n737), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n870), .A2(new_n709), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT125), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n914), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n950), .A2(G197gat), .A3(new_n263), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT126), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n885), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n595), .B1(new_n866), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n826), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT57), .B1(new_n955), .B2(new_n563), .ZN(new_n956));
  INV_X1    g755(.A(new_n891), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n737), .B(new_n944), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G197gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n960));
  INV_X1    g759(.A(new_n951), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n952), .A2(new_n962), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n661), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G204gat), .ZN(new_n965));
  INV_X1    g764(.A(new_n950), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n738), .A2(G204gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n965), .B(new_n969), .C1(new_n972), .C2(new_n973), .ZN(G1353gat));
  OR3_X1    g773(.A1(new_n950), .A2(G211gat), .A3(new_n595), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n892), .A2(new_n596), .A3(new_n944), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  INV_X1    g778(.A(G218gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n966), .A2(new_n980), .A3(new_n794), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n946), .A2(new_n636), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n980), .ZN(G1355gat));
endmodule


