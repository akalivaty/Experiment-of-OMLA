//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n189), .A3(new_n190), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n191), .A2(new_n192), .B1(KEYINPUT2), .B2(G113), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT66), .B1(new_n193), .B2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n193), .A2(new_n199), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT30), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT0), .A3(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(G137), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT11), .A3(G134), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n221), .A3(new_n224), .A4(new_n219), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n223), .A2(KEYINPUT67), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n223), .B2(new_n225), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n215), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n220), .A2(G134), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n217), .A2(G137), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n225), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT64), .A2(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT64), .A2(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n212), .A3(G128), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n205), .A3(new_n236), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n239), .A2(G128), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n240), .B2(new_n212), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n232), .B1(new_n225), .B2(new_n231), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n234), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n203), .B1(new_n228), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n223), .A2(new_n225), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n215), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n237), .A2(new_n212), .A3(G128), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n212), .B1(new_n239), .B2(G128), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n225), .B(new_n231), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(KEYINPUT30), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n202), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(G101), .ZN(new_n255));
  INV_X1    g069(.A(G210), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n256), .A2(G237), .A3(G953), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n255), .B(new_n257), .Z(new_n258));
  XOR2_X1   g072(.A(new_n200), .B(new_n201), .Z(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n228), .A3(new_n244), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT31), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n253), .A2(KEYINPUT31), .A3(new_n258), .A4(new_n260), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n246), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n223), .A2(KEYINPUT67), .A3(new_n225), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n214), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n248), .A2(new_n249), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n270), .A2(new_n233), .A3(new_n242), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n265), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n228), .A2(new_n244), .A3(KEYINPUT71), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n259), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n277));
  NAND2_X1  g091(.A1(new_n228), .A2(new_n244), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n202), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n251), .A2(new_n202), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n258), .B(KEYINPUT69), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n263), .A2(new_n264), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n187), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n253), .A2(new_n260), .ZN(new_n289));
  INV_X1    g103(.A(new_n258), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n291), .B(new_n292), .C1(new_n282), .C2(new_n284), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n278), .A2(new_n202), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n260), .A3(KEYINPUT72), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n278), .A2(new_n297), .A3(new_n202), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(KEYINPUT28), .A3(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(KEYINPUT29), .A3(new_n258), .A4(new_n276), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G472), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n263), .A2(new_n264), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n282), .A2(new_n284), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n287), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n306), .B2(KEYINPUT32), .ZN(new_n307));
  NOR4_X1   g121(.A1(new_n285), .A2(KEYINPUT73), .A3(new_n187), .A4(new_n287), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n288), .B(new_n302), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G217), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(G234), .B2(new_n294), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n194), .A2(G128), .ZN(new_n313));
  INV_X1    g127(.A(G128), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT24), .B(G110), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(KEYINPUT23), .A3(G119), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n313), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n322), .B2(G110), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(G146), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n323), .A2(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n204), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n325), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n329), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n204), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n322), .A2(G110), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n336), .B(new_n337), .C1(new_n316), .C2(new_n317), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT22), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(G137), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n333), .A2(new_n338), .A3(new_n343), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n294), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT25), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n312), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n312), .B2(new_n348), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n309), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G214), .B1(G237), .B2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(G234), .A2(G237), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(G952), .A3(new_n340), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT21), .B(G898), .Z(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(G902), .A3(G953), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(G107), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT78), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G107), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n370), .A2(new_n372), .A3(KEYINPUT78), .A4(G104), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n368), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n376), .B(KEYINPUT3), .C1(new_n367), .C2(G107), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(G104), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n376), .B1(new_n379), .B2(KEYINPUT3), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G101), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n367), .B2(G107), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT77), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n377), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n370), .A2(new_n372), .A3(G104), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n373), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n385), .A2(new_n389), .A3(new_n390), .A4(new_n368), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(G101), .C1(new_n375), .C2(new_n381), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n202), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n396));
  OAI21_X1  g210(.A(G113), .B1(new_n396), .B2(new_n195), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n199), .B2(new_n396), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n193), .A2(new_n199), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n368), .A2(new_n379), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n391), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n401), .B1(new_n391), .B2(new_n403), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n395), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n408));
  XOR2_X1   g222(.A(G110), .B(G122), .Z(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT84), .ZN(new_n411));
  INV_X1    g225(.A(new_n409), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n395), .B2(new_n406), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n408), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n413), .A2(new_n408), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n395), .A2(new_n406), .A3(new_n412), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n411), .A2(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n214), .A2(G125), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n241), .B2(G125), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n340), .A2(G224), .ZN(new_n422));
  XOR2_X1   g236(.A(new_n421), .B(new_n422), .Z(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n407), .A2(new_n409), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n426));
  AND4_X1   g240(.A1(new_n414), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n414), .B1(new_n413), .B2(new_n408), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n423), .B(new_n426), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT85), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G210), .B1(G237), .B2(G902), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n391), .A2(new_n403), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n397), .B1(KEYINPUT5), .B2(new_n199), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n399), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n409), .B(KEYINPUT8), .Z(new_n437));
  NAND2_X1  g251(.A1(new_n400), .A2(new_n433), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n417), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n422), .A2(KEYINPUT7), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n421), .B(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n294), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT86), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n431), .A2(new_n432), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n432), .B1(new_n431), .B2(new_n444), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n357), .B(new_n366), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT89), .ZN(new_n448));
  NOR2_X1   g262(.A1(KEYINPUT87), .A2(G143), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G237), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n340), .A3(G214), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT87), .A2(G143), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(G214), .A3(new_n451), .A4(new_n340), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n448), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n456), .A2(new_n224), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n336), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n456), .A2(new_n224), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n457), .A2(KEYINPUT18), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(KEYINPUT18), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n326), .B(new_n204), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n461), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G113), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n367), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G475), .ZN(new_n475));
  INV_X1    g289(.A(new_n473), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n458), .A2(new_n461), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n326), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT19), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n330), .B1(new_n480), .B2(G146), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n470), .B(new_n476), .C1(new_n477), .C2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n474), .A2(new_n475), .A3(new_n294), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n476), .A2(KEYINPUT90), .ZN(new_n486));
  AOI21_X1  g300(.A(G902), .B1(new_n471), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n486), .B2(new_n471), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n483), .A2(new_n484), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT91), .B(G122), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n492), .A2(new_n196), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n372), .B1(new_n493), .B2(KEYINPUT14), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n196), .A2(G122), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n492), .A2(new_n196), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G128), .B(G143), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(new_n217), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n493), .B(new_n495), .C1(KEYINPUT14), .C2(new_n372), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n372), .A3(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(G107), .B1(new_n497), .B2(new_n496), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n499), .A2(KEYINPUT13), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n314), .A2(KEYINPUT13), .A3(G143), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n217), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n506), .A2(new_n508), .B1(new_n217), .B2(new_n499), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n505), .A2(KEYINPUT92), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT92), .B1(new_n505), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n502), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT9), .B(G234), .Z(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(G217), .A3(new_n340), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n514), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n502), .B(new_n516), .C1(new_n510), .C2(new_n511), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT93), .A3(new_n294), .ZN(new_n519));
  INV_X1    g333(.A(G478), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n519), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n491), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G221), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n513), .B2(new_n294), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(KEYINPUT76), .Z(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G140), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n340), .A2(G227), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n527), .B(new_n528), .Z(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n226), .A2(new_n227), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n392), .A2(new_n215), .A3(new_n394), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n314), .B1(new_n535), .B2(KEYINPUT79), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n212), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n248), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n534), .B1(new_n539), .B2(new_n433), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT10), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n270), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n404), .B2(new_n405), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(KEYINPUT82), .B(new_n543), .C1(new_n404), .C2(new_n405), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n532), .B(new_n541), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n533), .A2(new_n540), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n531), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n530), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n433), .A2(KEYINPUT81), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n391), .A2(new_n401), .A3(new_n403), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT82), .B1(new_n555), .B2(new_n543), .ZN(new_n556));
  INV_X1    g370(.A(new_n547), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n550), .B(new_n531), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n433), .A2(new_n270), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n539), .A2(new_n433), .ZN(new_n561));
  OAI211_X1 g375(.A(KEYINPUT12), .B(new_n246), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n561), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n531), .B1(new_n563), .B2(new_n559), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n564), .B2(KEYINPUT12), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n565), .A3(new_n529), .ZN(new_n566));
  AOI211_X1 g380(.A(G469), .B(G902), .C1(new_n552), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n558), .A2(new_n565), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n530), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n532), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n558), .A3(new_n529), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n572), .A3(G469), .ZN(new_n573));
  NAND2_X1  g387(.A1(G469), .A2(G902), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n526), .B1(new_n567), .B2(new_n575), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n447), .A2(new_n523), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n356), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G101), .ZN(G3));
  INV_X1    g393(.A(new_n353), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n304), .A2(new_n305), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n294), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G472), .ZN(new_n583));
  INV_X1    g397(.A(new_n306), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR4_X1   g399(.A1(new_n447), .A2(new_n580), .A3(new_n576), .A4(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n515), .A2(new_n587), .A3(new_n517), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n587), .B1(new_n515), .B2(new_n517), .ZN(new_n590));
  OAI211_X1 g404(.A(G478), .B(new_n294), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n518), .A2(KEYINPUT33), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n588), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n595), .A2(KEYINPUT94), .A3(G478), .A4(new_n294), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n518), .A2(new_n294), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n520), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n593), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n586), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT34), .B(G104), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT95), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n603), .B(new_n605), .ZN(G6));
  NOR2_X1   g420(.A1(new_n522), .A2(new_n600), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n586), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT35), .B(G107), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  INV_X1    g424(.A(new_n352), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n343), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n339), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n294), .A3(new_n312), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n611), .A2(KEYINPUT97), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n618));
  INV_X1    g432(.A(new_n616), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n352), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n577), .A2(new_n584), .A3(new_n583), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT98), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT37), .B(G110), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  NAND2_X1  g439(.A1(new_n302), .A2(new_n288), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n581), .A2(KEYINPUT32), .A3(new_n286), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT73), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n306), .A2(new_n303), .A3(KEYINPUT32), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n576), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n357), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n419), .B1(new_n418), .B2(new_n423), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n429), .A2(KEYINPUT85), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n444), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n432), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n431), .A2(new_n432), .A3(new_n444), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n633), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n607), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n360), .B1(new_n364), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n632), .A2(new_n640), .A3(new_n621), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT99), .B(G128), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G30));
  NAND2_X1  g461(.A1(new_n638), .A2(new_n639), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT38), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n296), .A2(new_n298), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT100), .B1(new_n650), .B2(new_n283), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n261), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n650), .A2(new_n283), .A3(KEYINPUT100), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n294), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n631), .A2(new_n288), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n611), .A2(new_n616), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n657), .A2(new_n491), .A3(new_n522), .A4(new_n633), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n649), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n526), .ZN(new_n660));
  INV_X1    g474(.A(new_n575), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n552), .A2(new_n566), .ZN(new_n662));
  INV_X1    g476(.A(G469), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n294), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n643), .B(KEYINPUT39), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT40), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT101), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n206), .ZN(G45));
  INV_X1    g485(.A(new_n643), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n599), .A2(new_n600), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n632), .A2(new_n640), .A3(new_n621), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n357), .B(new_n621), .C1(new_n445), .C2(new_n446), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n632), .A4(new_n674), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  AOI21_X1  g496(.A(new_n529), .B1(new_n571), .B2(new_n558), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n558), .A2(new_n565), .A3(new_n529), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n294), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  INV_X1    g500(.A(new_n525), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n664), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n686), .A2(new_n664), .A3(new_n690), .A4(new_n687), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(new_n447), .A3(new_n354), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n602), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT41), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G113), .ZN(G15));
  NAND2_X1  g510(.A1(new_n693), .A2(new_n607), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  NOR2_X1   g512(.A1(new_n692), .A2(new_n677), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n523), .B(new_n365), .C1(new_n627), .C2(new_n631), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  AND4_X1   g516(.A1(new_n357), .A2(new_n648), .A3(new_n689), .A4(new_n691), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n519), .B(new_n521), .Z(new_n704));
  AND3_X1   g518(.A1(new_n704), .A2(KEYINPUT105), .A3(new_n600), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT105), .B1(new_n704), .B2(new_n600), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n366), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT104), .B(G472), .Z(new_n711));
  NAND2_X1  g525(.A1(new_n582), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n304), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n283), .B1(new_n299), .B2(new_n276), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n286), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n580), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n703), .A2(new_n709), .A3(new_n710), .A4(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n640), .A2(new_n691), .A3(new_n689), .A4(new_n717), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT106), .B1(new_n719), .B2(new_n708), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT107), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NAND3_X1  g537(.A1(new_n712), .A2(new_n657), .A3(new_n715), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n673), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n640), .A3(new_n691), .A4(new_n689), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  INV_X1    g541(.A(new_n628), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n353), .B1(new_n626), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n445), .A2(new_n446), .A3(new_n633), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n525), .B1(new_n661), .B2(new_n664), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n731), .A2(new_n674), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n638), .A3(new_n357), .A4(new_n639), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n354), .A3(new_n673), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n734), .B1(new_n736), .B2(KEYINPUT42), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n354), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n644), .A2(KEYINPUT108), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n644), .A2(KEYINPUT108), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NAND2_X1  g557(.A1(new_n599), .A2(new_n491), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n585), .A3(new_n657), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n732), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n569), .A2(new_n572), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(G469), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n574), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n756), .B(G469), .C1(new_n753), .C2(G902), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n664), .A3(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n758), .A2(new_n687), .A3(new_n666), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n748), .A2(KEYINPUT109), .A3(new_n732), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n751), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  AOI21_X1  g576(.A(KEYINPUT47), .B1(new_n758), .B2(new_n687), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n758), .A2(KEYINPUT47), .A3(new_n687), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n673), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n638), .A2(new_n357), .A3(new_n639), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n309), .A3(new_n353), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(KEYINPUT110), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n601), .A2(new_n641), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n356), .A2(new_n577), .B1(new_n586), .B2(new_n776), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n693), .A2(new_n776), .B1(new_n699), .B2(new_n700), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n721), .A3(new_n622), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n309), .A2(new_n665), .ZN(new_n780));
  INV_X1    g594(.A(new_n621), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n780), .A2(new_n767), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT111), .B1(new_n523), .B2(new_n643), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n491), .A2(new_n522), .A3(new_n785), .A4(new_n672), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n632), .A2(new_n732), .A3(new_n787), .A4(new_n621), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n724), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n732), .A2(new_n674), .A3(new_n792), .A4(new_n733), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n737), .A3(new_n742), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n779), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n645), .A2(new_n726), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n656), .A2(new_n672), .A3(new_n733), .ZN(new_n798));
  INV_X1    g612(.A(new_n657), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n640), .A3(new_n799), .A4(new_n707), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n681), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n796), .B1(new_n680), .B2(new_n676), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .A3(new_n800), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n795), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n783), .B1(new_n782), .B2(new_n787), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n789), .A2(KEYINPUT112), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n793), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n737), .A2(new_n742), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n721), .A2(new_n778), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n586), .A2(new_n776), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n578), .A2(new_n622), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n813), .A2(KEYINPUT53), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(new_n804), .B2(new_n800), .ZN(new_n818));
  AND4_X1   g632(.A1(KEYINPUT52), .A2(new_n681), .A3(new_n797), .A4(new_n800), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n779), .A2(new_n794), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT113), .B1(new_n824), .B2(new_n806), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n775), .B(new_n808), .C1(new_n822), .C2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n692), .A2(new_n359), .A3(new_n767), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n827), .A2(new_n746), .ZN(new_n828));
  INV_X1    g642(.A(new_n729), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  INV_X1    g645(.A(new_n656), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n827), .A2(new_n353), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n602), .ZN(new_n836));
  INV_X1    g650(.A(G952), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n716), .A2(new_n580), .A3(new_n359), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n691), .A2(new_n746), .A3(new_n689), .A4(new_n838), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n837), .B(G953), .C1(new_n839), .C2(new_n640), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n831), .A2(new_n836), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n817), .A2(new_n820), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT54), .B1(new_n844), .B2(new_n807), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n826), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n599), .A2(new_n600), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n834), .A2(new_n835), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n649), .A2(new_n357), .ZN(new_n849));
  NAND2_X1  g663(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n849), .A2(new_n839), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n849), .B2(new_n839), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n851), .A2(new_n852), .B1(KEYINPUT114), .B2(KEYINPUT50), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n686), .A2(new_n664), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n660), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n764), .A2(new_n765), .A3(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(new_n732), .A3(new_n746), .A4(new_n838), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n828), .A2(new_n792), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n848), .A2(new_n853), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT51), .Z(new_n860));
  OAI22_X1  g674(.A1(new_n846), .A2(new_n860), .B1(G952), .B2(G953), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n854), .B(KEYINPUT49), .Z(new_n862));
  NOR4_X1   g676(.A1(new_n862), .A2(new_n633), .A3(new_n660), .A4(new_n744), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n649), .A2(new_n580), .A3(new_n656), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(KEYINPUT117), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(G75));
  XOR2_X1   g684(.A(new_n418), .B(new_n423), .Z(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT55), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n821), .B1(new_n817), .B2(new_n820), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n824), .A2(KEYINPUT113), .A3(new_n806), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n807), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n878), .A2(new_n256), .A3(new_n294), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n875), .B1(new_n879), .B2(KEYINPUT56), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n837), .A2(G953), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT119), .Z(new_n882));
  OAI21_X1  g696(.A(new_n808), .B1(new_n822), .B2(new_n825), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(G210), .A3(G902), .ZN(new_n884));
  INV_X1    g698(.A(new_n875), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n874), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n880), .A2(new_n889), .A3(new_n886), .A4(new_n882), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(G51));
  INV_X1    g705(.A(new_n882), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n883), .A2(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(KEYINPUT121), .A3(new_n826), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n878), .A2(KEYINPUT121), .A3(new_n775), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n574), .B(KEYINPUT57), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n662), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n878), .A2(new_n294), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(G469), .A3(new_n753), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n892), .B1(new_n898), .B2(new_n900), .ZN(G54));
  NAND3_X1  g715(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n474), .A2(new_n482), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n892), .B1(new_n904), .B2(new_n905), .ZN(G60));
  NAND2_X1  g720(.A1(new_n826), .A2(new_n845), .ZN(new_n907));
  NAND2_X1  g721(.A1(G478), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT59), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n595), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n892), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n894), .A2(new_n595), .A3(new_n895), .A4(new_n909), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(G63));
  XNOR2_X1  g727(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n310), .A2(new_n294), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n883), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n345), .A2(new_n346), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n892), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n883), .A2(new_n615), .A3(new_n916), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n883), .A2(KEYINPUT123), .A3(new_n615), .A4(new_n916), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n919), .A2(new_n922), .A3(KEYINPUT61), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(G66));
  INV_X1    g742(.A(G224), .ZN(new_n929));
  OAI21_X1  g743(.A(G953), .B1(new_n362), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n779), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(G953), .ZN(new_n932));
  INV_X1    g746(.A(new_n418), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(G898), .B2(new_n340), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n932), .B(new_n934), .ZN(G69));
  AOI21_X1  g749(.A(new_n340), .B1(G227), .B2(G900), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n804), .B1(new_n668), .B2(new_n659), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n773), .A2(new_n761), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n941));
  INV_X1    g755(.A(new_n356), .ZN(new_n942));
  INV_X1    g756(.A(new_n776), .ZN(new_n943));
  NOR4_X1   g757(.A1(new_n942), .A2(new_n667), .A3(new_n767), .A4(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n773), .A2(new_n941), .A3(new_n761), .A4(new_n938), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT125), .B1(new_n947), .B2(new_n944), .ZN(new_n948));
  AOI21_X1  g762(.A(G953), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n245), .A2(new_n252), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT124), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(new_n480), .Z(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n759), .A2(new_n640), .A3(new_n707), .A4(new_n829), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n804), .A2(new_n737), .A3(new_n742), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n773), .A2(new_n761), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n340), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n340), .A2(G900), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n958), .A2(new_n963), .A3(new_n960), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n952), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n936), .B1(new_n954), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n963), .B1(new_n958), .B2(new_n960), .ZN(new_n967));
  AOI211_X1 g781(.A(KEYINPUT126), .B(new_n959), .C1(new_n957), .C2(new_n340), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n953), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n936), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n969), .B(new_n970), .C1(new_n949), .C2(new_n953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n966), .A2(new_n971), .ZN(G72));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n957), .B2(new_n779), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n289), .B(KEYINPUT127), .Z(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n290), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n291), .A2(new_n261), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n974), .B(new_n978), .C1(new_n844), .C2(new_n807), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n882), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n946), .A2(new_n948), .A3(new_n931), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n976), .B1(new_n981), .B2(new_n974), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n982), .B2(new_n258), .ZN(G57));
endmodule


