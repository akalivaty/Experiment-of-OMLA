//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT96), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT96), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n205), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(new_n202), .A3(new_n203), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G43gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G50gat), .ZN(new_n213));
  INV_X1    g012(.A(G50gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G43gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT15), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n207), .A2(new_n211), .A3(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(KEYINPUT94), .A2(G43gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT95), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT94), .A2(G43gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n214), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT15), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n214), .A3(new_n220), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT95), .A3(new_n213), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n217), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n210), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT93), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n227), .A2(new_n228), .B1(G29gat), .B2(G36gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n209), .A2(KEYINPUT93), .A3(new_n210), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n216), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(KEYINPUT97), .B(KEYINPUT17), .C1(new_n226), .C2(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n207), .A2(new_n211), .A3(new_n216), .ZN(new_n233));
  INV_X1    g032(.A(new_n225), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n221), .A2(new_n222), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n231), .ZN(new_n237));
  OR2_X1    g036(.A1(KEYINPUT97), .A2(KEYINPUT17), .ZN(new_n238));
  NAND2_X1  g037(.A1(KEYINPUT97), .A2(KEYINPUT17), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT7), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT7), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(G85gat), .A3(G92gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247));
  INV_X1    g046(.A(G85gat), .ZN(new_n248));
  INV_X1    g047(.A(G92gat), .ZN(new_n249));
  AOI22_X1  g048(.A1(KEYINPUT8), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G99gat), .B(G106gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n246), .A2(new_n250), .A3(new_n252), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n226), .A2(new_n231), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n257), .B(new_n258), .C1(new_n256), .C2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G190gat), .B(G218gat), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n262), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT103), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT102), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT103), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(new_n267), .A3(new_n262), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G134gat), .B(G162gat), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n265), .A2(new_n268), .A3(new_n266), .A4(new_n272), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278));
  INV_X1    g077(.A(G1gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT16), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G1gat), .B2(new_n278), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n282), .A2(G8gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(G8gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT99), .ZN(new_n286));
  INV_X1    g085(.A(G57gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G64gat), .ZN(new_n288));
  INV_X1    g087(.A(G64gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G57gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G71gat), .ZN(new_n292));
  INV_X1    g091(.A(G78gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G71gat), .A2(G78gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT9), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n291), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n296), .B1(new_n298), .B2(new_n291), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n286), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n291), .A2(new_n298), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n294), .A2(new_n295), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n291), .A2(new_n296), .A3(new_n298), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT99), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n285), .B1(KEYINPUT21), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n310), .B(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n307), .A2(KEYINPUT21), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G155gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(G231gat), .A2(G233gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G183gat), .B(G211gat), .Z(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  XNOR2_X1  g118(.A(new_n314), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n313), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n277), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G78gat), .B(G106gat), .Z(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT31), .B(G50gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G228gat), .A2(G233gat), .ZN(new_n328));
  XOR2_X1   g127(.A(G211gat), .B(G218gat), .Z(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(G218gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT22), .B1(new_n330), .B2(G211gat), .ZN(new_n331));
  XOR2_X1   g130(.A(G197gat), .B(G204gat), .Z(new_n332));
  OAI21_X1  g131(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  INV_X1    g133(.A(G218gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT76), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G218gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n338), .A3(G211gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n329), .ZN(new_n342));
  INV_X1    g141(.A(new_n332), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n333), .A2(new_n334), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n343), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT77), .A3(new_n329), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n345), .A2(KEYINPUT87), .A3(new_n346), .A4(new_n348), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355));
  INV_X1    g154(.A(G141gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(G148gat), .ZN(new_n357));
  INV_X1    g156(.A(G148gat), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT80), .B1(new_n358), .B2(G141gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(G141gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT81), .ZN(new_n362));
  XNOR2_X1  g161(.A(G155gat), .B(G162gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT2), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n357), .C1(new_n359), .C2(new_n360), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n362), .A2(new_n363), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n356), .A2(G148gat), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT79), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n356), .A2(G148gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n358), .A2(G141gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n365), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n363), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT82), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n368), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n354), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n367), .A2(new_n363), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n361), .A2(KEYINPUT81), .B1(KEYINPUT2), .B2(new_n364), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n385), .A2(new_n386), .B1(new_n376), .B2(new_n375), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n387), .B2(new_n352), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n345), .A2(new_n348), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n328), .B1(new_n383), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n333), .A2(new_n344), .ZN(new_n393));
  INV_X1    g192(.A(new_n384), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n387), .B1(new_n395), .B2(new_n352), .ZN(new_n396));
  INV_X1    g195(.A(new_n328), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n390), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(G22gat), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  INV_X1    g199(.A(G22gat), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n390), .B1(new_n354), .B2(new_n382), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n400), .B(new_n401), .C1(new_n402), .C2(new_n328), .ZN(new_n403));
  AOI211_X1 g202(.A(KEYINPUT88), .B(new_n327), .C1(new_n399), .C2(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n399), .A2(KEYINPUT88), .A3(new_n403), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT88), .B1(new_n399), .B2(new_n403), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n407), .B2(new_n327), .ZN(new_n408));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(new_n289), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT66), .B(G169gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT23), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G176gat), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT25), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417));
  INV_X1    g216(.A(G169gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n413), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT65), .ZN(new_n421));
  INV_X1    g220(.A(G183gat), .ZN(new_n422));
  INV_X1    g221(.A(G190gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(G183gat), .A2(G190gat), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT24), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n428), .A2(KEYINPUT64), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT64), .B1(new_n428), .B2(new_n429), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n426), .B(new_n427), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n420), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n419), .A2(KEYINPUT26), .ZN(new_n434));
  NOR2_X1   g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT26), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n417), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT27), .B(G183gat), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT28), .A3(new_n423), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT28), .B1(new_n440), .B2(new_n423), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n439), .B(new_n428), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n445), .B(new_n427), .C1(G183gat), .C2(G190gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n419), .A2(new_n413), .B1(new_n447), .B2(new_n417), .ZN(new_n448));
  NAND3_X1  g247(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n435), .A2(KEYINPUT23), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n446), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT25), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n444), .A3(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(G226gat), .A2(G233gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n453), .B2(new_n394), .ZN(new_n457));
  OR3_X1    g256(.A1(new_n456), .A2(new_n457), .A3(new_n389), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n423), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT28), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n438), .B1(new_n461), .B2(new_n441), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n462), .A2(new_n428), .B1(KEYINPUT25), .B2(new_n451), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n463), .B2(new_n433), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n455), .B1(new_n464), .B2(new_n454), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n389), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n411), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n389), .B1(new_n456), .B2(new_n457), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(KEYINPUT37), .C1(new_n389), .C2(new_n465), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n467), .A2(new_n411), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n458), .A2(KEYINPUT37), .A3(new_n466), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n470), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G120gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G113gat), .ZN(new_n480));
  INV_X1    g279(.A(G113gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G120gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT68), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G127gat), .B(G134gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT1), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n479), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G127gat), .ZN(new_n489));
  INV_X1    g288(.A(G134gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G127gat), .A2(G134gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(G113gat), .B(G120gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(KEYINPUT1), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT69), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n488), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n488), .B2(new_n494), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(KEYINPUT4), .A3(new_n387), .ZN(new_n499));
  NAND2_X1  g298(.A1(G225gat), .A2(G233gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n488), .A2(new_n494), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n368), .A2(new_n502), .A3(new_n377), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n502), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n352), .B1(new_n379), .B2(new_n381), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n368), .A2(new_n380), .A3(new_n377), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n380), .B1(new_n368), .B2(new_n377), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n508), .B(KEYINPUT3), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n387), .A2(new_n352), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n499), .B(new_n505), .C1(new_n509), .C2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n502), .B1(new_n379), .B2(new_n381), .ZN(new_n516));
  INV_X1    g315(.A(new_n503), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n501), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT3), .B1(new_n510), .B2(new_n511), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT83), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n522), .A2(new_n506), .A3(new_n512), .A4(new_n513), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n387), .B(new_n504), .C1(new_n497), .C2(new_n496), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(KEYINPUT85), .A3(new_n525), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n519), .A2(new_n501), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n523), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n520), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT86), .ZN(new_n534));
  XNOR2_X1  g333(.A(G1gat), .B(G29gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT0), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G57gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G85gat), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT6), .A4(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(KEYINPUT6), .A3(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT86), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n538), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n543));
  INV_X1    g342(.A(new_n538), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n520), .A2(new_n544), .A3(new_n532), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n478), .A2(new_n539), .A3(new_n541), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n500), .B1(new_n523), .B2(new_n530), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT39), .ZN(new_n549));
  AOI211_X1 g348(.A(KEYINPUT89), .B(new_n538), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT85), .B1(new_n524), .B2(new_n525), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n524), .A2(KEYINPUT85), .A3(new_n525), .ZN(new_n553));
  OAI22_X1  g352(.A1(new_n509), .A2(new_n514), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n549), .A3(new_n501), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n551), .B1(new_n555), .B2(new_n544), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n548), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n516), .A2(new_n517), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n549), .B1(new_n559), .B2(new_n500), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n560), .A2(KEYINPUT90), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(KEYINPUT90), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT91), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT40), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n542), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n555), .A2(new_n544), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT89), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n555), .A2(new_n551), .A3(new_n544), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n565), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT30), .B1(new_n467), .B2(new_n411), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n474), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n408), .B(new_n547), .C1(new_n566), .C2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577));
  XNOR2_X1  g376(.A(G15gat), .B(G43gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT72), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(new_n292), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G99gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n453), .A2(new_n498), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n496), .A2(new_n497), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n463), .A2(new_n583), .A3(new_n433), .ZN(new_n584));
  NAND2_X1  g383(.A1(G227gat), .A2(G233gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT33), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n581), .B1(new_n589), .B2(KEYINPUT70), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT70), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n591), .A3(new_n588), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(KEYINPUT32), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT71), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT71), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(new_n595), .A3(KEYINPUT32), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n590), .A2(new_n592), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n587), .B(KEYINPUT32), .C1(new_n581), .C2(new_n588), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n586), .B1(new_n582), .B2(new_n584), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(new_n585), .B2(KEYINPUT74), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n597), .A3(new_n598), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n577), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n597), .A2(new_n603), .A3(new_n598), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n603), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n599), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n597), .A2(KEYINPUT75), .A3(new_n603), .A4(new_n598), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n609), .B1(new_n577), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n408), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n541), .A2(new_n546), .A3(new_n539), .ZN(new_n619));
  INV_X1    g418(.A(new_n574), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n617), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n576), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n408), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n619), .A2(KEYINPUT35), .A3(new_n620), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n408), .A2(new_n619), .A3(new_n620), .A4(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT35), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n625), .A2(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n323), .B1(new_n623), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n285), .B1(new_n232), .B2(new_n240), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n284), .A2(new_n283), .B1(new_n236), .B2(new_n237), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT18), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT18), .ZN(new_n637));
  INV_X1    g436(.A(new_n635), .ZN(new_n638));
  NOR4_X1   g437(.A1(new_n632), .A2(new_n637), .A3(new_n633), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n642));
  XNOR2_X1  g441(.A(G113gat), .B(G141gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G169gat), .B(G197gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  INV_X1    g446(.A(new_n285), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n259), .ZN(new_n649));
  INV_X1    g448(.A(new_n633), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n635), .B(KEYINPUT13), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n640), .A2(new_n641), .A3(new_n647), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n241), .A2(new_n648), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n650), .A3(new_n635), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n637), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n634), .A2(KEYINPUT18), .A3(new_n635), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n647), .A4(new_n654), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT98), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n640), .A2(new_n654), .ZN(new_n662));
  INV_X1    g461(.A(new_n647), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n655), .A2(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n301), .A2(new_n256), .A3(new_n306), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n299), .A2(new_n300), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n253), .A2(KEYINPUT104), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n251), .A2(KEYINPUT104), .A3(new_n253), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n666), .A2(new_n255), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n256), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n307), .A2(KEYINPUT10), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n665), .A2(new_n669), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n665), .A2(new_n669), .A3(KEYINPUT105), .A4(new_n676), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n672), .B1(new_n681), .B2(new_n671), .ZN(new_n682));
  XNOR2_X1  g481(.A(G120gat), .B(G148gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n415), .ZN(new_n684));
  INV_X1    g483(.A(G204gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n664), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n631), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n619), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(new_n279), .ZN(G1324gat));
  NOR2_X1   g492(.A1(new_n691), .A2(new_n620), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT16), .ZN(new_n695));
  INV_X1    g494(.A(G8gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n694), .A2(new_n696), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(KEYINPUT42), .B2(new_n699), .ZN(G1325gat));
  INV_X1    g501(.A(new_n691), .ZN(new_n703));
  AOI21_X1  g502(.A(G15gat), .B1(new_n703), .B2(new_n627), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n617), .A2(G15gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT106), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n703), .B2(new_n706), .ZN(G1326gat));
  NAND3_X1  g506(.A1(new_n631), .A2(new_n690), .A3(new_n618), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n401), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(G22gat), .A3(new_n712), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1327gat));
  AOI211_X1 g517(.A(new_n322), .B(new_n277), .C1(new_n623), .C2(new_n630), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n719), .A2(new_n690), .ZN(new_n720));
  INV_X1    g519(.A(new_n619), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n202), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT45), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n689), .B(KEYINPUT108), .ZN(new_n724));
  INV_X1    g523(.A(new_n664), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n725), .A3(new_n321), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT109), .ZN(new_n727));
  NAND2_X1  g526(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n623), .A2(new_n630), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n276), .ZN(new_n733));
  AOI211_X1 g532(.A(new_n277), .B(new_n729), .C1(new_n623), .C2(new_n630), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G29gat), .B1(new_n735), .B2(new_n619), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n723), .A2(new_n736), .ZN(G1328gat));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n690), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n738), .A2(G36gat), .A3(new_n620), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n735), .B2(new_n620), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(G1329gat));
  NAND2_X1  g543(.A1(new_n218), .A2(new_n220), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n720), .A2(new_n745), .A3(new_n627), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n617), .B(new_n727), .C1(new_n733), .C2(new_n734), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n748), .B2(new_n745), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1330gat));
  OAI211_X1 g550(.A(new_n618), .B(new_n727), .C1(new_n733), .C2(new_n734), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n752), .A2(new_n753), .A3(G50gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n752), .B2(G50gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n738), .A2(G50gat), .A3(new_n408), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n752), .A2(G50gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n720), .A2(new_n214), .A3(new_n618), .ZN(new_n759));
  AND4_X1   g558(.A1(KEYINPUT112), .A2(new_n758), .A3(KEYINPUT48), .A4(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n752), .B2(G50gat), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT112), .B1(new_n762), .B2(new_n759), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n757), .A2(KEYINPUT48), .B1(new_n760), .B2(new_n763), .ZN(G1331gat));
  NOR2_X1   g563(.A1(new_n724), .A2(new_n725), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n631), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n619), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(new_n287), .ZN(G1332gat));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n620), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n766), .A2(KEYINPUT113), .A3(new_n616), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT113), .B1(new_n766), .B2(new_n616), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n292), .ZN(new_n778));
  INV_X1    g577(.A(new_n766), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n292), .B1(new_n779), .B2(new_n617), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n774), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  AOI211_X1 g581(.A(KEYINPUT50), .B(new_n780), .C1(new_n777), .C2(new_n292), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(G1334gat));
  NOR2_X1   g583(.A1(new_n766), .A2(new_n408), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(new_n293), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n322), .A2(new_n725), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n689), .B(new_n787), .C1(new_n733), .C2(new_n734), .ZN(new_n788));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788), .B2(new_n619), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n719), .A2(KEYINPUT51), .A3(new_n664), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n719), .B2(new_n664), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(new_n248), .A3(new_n721), .ZN(new_n793));
  INV_X1    g592(.A(new_n689), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  INV_X1    g594(.A(new_n724), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n620), .A2(G92gat), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n796), .B(new_n797), .C1(new_n790), .C2(new_n791), .ZN(new_n798));
  OAI21_X1  g597(.A(G92gat), .B1(new_n788), .B2(new_n620), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1337gat));
  INV_X1    g603(.A(new_n617), .ZN(new_n805));
  OAI21_X1  g604(.A(G99gat), .B1(new_n788), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(G99gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n807), .A3(new_n627), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n808), .B2(new_n794), .ZN(G1338gat));
  NOR2_X1   g608(.A1(new_n408), .A2(G106gat), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n796), .B(new_n810), .C1(new_n790), .C2(new_n791), .ZN(new_n811));
  OAI21_X1  g610(.A(G106gat), .B1(new_n788), .B2(new_n408), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1339gat));
  NOR3_X1   g616(.A1(new_n323), .A2(new_n689), .A3(new_n725), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n681), .A2(new_n671), .B1(KEYINPUT114), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n681), .B2(new_n671), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT55), .B(new_n686), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n824), .A2(new_n825), .A3(new_n687), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n824), .B2(new_n687), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n655), .A2(new_n661), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT116), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n634), .A2(new_n635), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n646), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n820), .B(new_n821), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n686), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n828), .A2(new_n276), .A3(new_n834), .A4(new_n838), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n829), .A2(new_n689), .A3(new_n833), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT55), .B1(new_n835), .B2(new_n686), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n664), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n828), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n843), .B2(new_n276), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n818), .B1(new_n844), .B2(new_n321), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n619), .A3(new_n574), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n625), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n481), .A3(new_n725), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n618), .A2(new_n616), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n664), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n851), .ZN(G1340gat));
  NAND3_X1  g651(.A1(new_n847), .A2(new_n479), .A3(new_n689), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n850), .B2(new_n724), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(G1341gat));
  NOR3_X1   g656(.A1(new_n850), .A2(new_n489), .A3(new_n321), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n860));
  AOI21_X1  g659(.A(G127gat), .B1(new_n847), .B2(new_n322), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G1342gat));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n490), .A3(new_n276), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n850), .B2(new_n277), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n619), .A2(new_n574), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n805), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n845), .B2(new_n408), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n824), .A2(new_n687), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n841), .A3(new_n664), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n876), .B2(new_n840), .ZN(new_n877));
  INV_X1    g676(.A(new_n840), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n838), .A2(new_n725), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n878), .B(KEYINPUT120), .C1(new_n879), .C2(new_n875), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n277), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n322), .B1(new_n881), .B2(new_n839), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT57), .B(new_n618), .C1(new_n882), .C2(new_n818), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n664), .B(new_n870), .C1(new_n873), .C2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n868), .B1(new_n884), .B2(new_n356), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n617), .A2(new_n408), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n664), .A2(G141gat), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n846), .A2(new_n888), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n884), .B2(new_n356), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n885), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI221_X1 g693(.A(new_n891), .B1(new_n868), .B2(KEYINPUT58), .C1(new_n884), .C2(new_n356), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(G1344gat));
  AND3_X1   g695(.A1(new_n846), .A2(new_n888), .A3(new_n889), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n358), .A3(new_n689), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n870), .B1(new_n873), .B2(new_n883), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n689), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(G148gat), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n794), .B(new_n870), .C1(new_n873), .C2(new_n883), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(G148gat), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT123), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n618), .B1(new_n882), .B2(new_n818), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n844), .A2(new_n321), .ZN(new_n912));
  INV_X1    g711(.A(new_n818), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n618), .A3(new_n871), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n617), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n689), .A3(new_n869), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n908), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n898), .B1(new_n907), .B2(new_n918), .ZN(G1345gat));
  AOI21_X1  g718(.A(G155gat), .B1(new_n897), .B2(new_n322), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n322), .A2(G155gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n899), .B2(new_n921), .ZN(G1346gat));
  AOI21_X1  g721(.A(G162gat), .B1(new_n897), .B2(new_n276), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n276), .A2(G162gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n899), .B2(new_n924), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n845), .A2(new_n721), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n574), .A3(new_n849), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n664), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n619), .A2(new_n914), .A3(new_n574), .A4(new_n625), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n664), .A2(new_n412), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1348gat));
  AOI21_X1  g731(.A(G176gat), .B1(new_n929), .B2(new_n689), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n927), .A2(new_n415), .A3(new_n724), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(G1349gat));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n926), .A2(new_n440), .A3(new_n574), .A4(new_n625), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n321), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n929), .A2(KEYINPUT125), .A3(new_n440), .A4(new_n322), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G183gat), .B1(new_n927), .B2(new_n321), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT60), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n940), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n423), .A3(new_n276), .ZN(new_n947));
  OAI21_X1  g746(.A(G190gat), .B1(new_n927), .B2(new_n277), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  NOR4_X1   g750(.A1(new_n845), .A2(new_n721), .A3(new_n620), .A4(new_n887), .ZN(new_n952));
  XNOR2_X1  g751(.A(KEYINPUT126), .B(G197gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n725), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n721), .A2(new_n620), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n916), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n956), .A2(new_n725), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n957), .B2(new_n953), .ZN(G1352gat));
  NAND3_X1  g757(.A1(new_n916), .A2(new_n796), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n916), .A2(new_n961), .A3(new_n796), .A4(new_n955), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(G204gat), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n952), .A2(new_n685), .A3(new_n689), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1353gat));
  INV_X1    g765(.A(G211gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n967), .A3(new_n322), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n916), .A2(new_n322), .A3(new_n955), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  AOI21_X1  g771(.A(G218gat), .B1(new_n952), .B2(new_n276), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n276), .A2(new_n330), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n956), .B2(new_n974), .ZN(G1355gat));
endmodule


