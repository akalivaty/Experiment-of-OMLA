//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT26), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n207), .A2(KEYINPUT27), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT27), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n217), .B1(new_n214), .B2(new_n216), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n208), .A2(KEYINPUT28), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT27), .B(G183gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT28), .B1(new_n222), .B2(new_n208), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n213), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n210), .B1(KEYINPUT23), .B2(new_n211), .ZN(new_n225));
  OR2_X1    g024(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT64), .B1(new_n205), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n211), .A2(new_n229), .A3(KEYINPUT23), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n225), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n207), .B2(new_n208), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n236));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n229), .B1(new_n211), .B2(KEYINPUT23), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n205), .A2(KEYINPUT64), .A3(new_n227), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n231), .B(new_n235), .C1(new_n241), .C2(KEYINPUT65), .ZN(new_n242));
  NAND4_X1  g041(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n234), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n233), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n239), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n225), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT25), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n224), .A2(new_n242), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G127gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(G134gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G127gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT68), .ZN(new_n255));
  INV_X1    g054(.A(G113gat), .ZN(new_n256));
  INV_X1    g055(.A(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g058(.A1(G113gat), .A2(G120gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  OR3_X1    g060(.A1(new_n253), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n260), .ZN(new_n264));
  NOR2_X1   g063(.A1(G113gat), .A2(G120gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n267));
  NOR2_X1   g066(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n250), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n224), .A2(new_n242), .A3(new_n272), .A4(new_n249), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n274), .A2(KEYINPUT70), .A3(new_n276), .A4(new_n277), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n202), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT72), .ZN(new_n284));
  XOR2_X1   g083(.A(G71gat), .B(G99gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n276), .B1(new_n274), .B2(new_n277), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n287), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n280), .B2(new_n281), .ZN(new_n298));
  NOR4_X1   g097(.A1(new_n298), .A2(new_n282), .A3(KEYINPUT73), .A4(new_n286), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n281), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n286), .B1(new_n301), .B2(KEYINPUT32), .ZN(new_n302));
  INV_X1    g101(.A(new_n298), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n296), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT75), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n296), .B(new_n307), .C1(new_n299), .C2(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n310), .A3(new_n314), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n315), .A2(new_n321), .A3(new_n317), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n325), .B(KEYINPUT77), .Z(new_n326));
  NAND2_X1  g125(.A1(new_n250), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n326), .B1(new_n250), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n324), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n222), .A2(new_n217), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n215), .A2(G183gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n207), .A2(KEYINPUT27), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT67), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n333), .A2(new_n334), .A3(G190gat), .ZN(new_n337));
  OAI22_X1  g136(.A1(new_n336), .A2(new_n220), .B1(KEYINPUT28), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n338), .A2(new_n213), .B1(KEYINPUT25), .B2(new_n248), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n339), .B2(new_n242), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n323), .B(new_n327), .C1(new_n340), .C2(new_n326), .ZN(new_n341));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n331), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT30), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n331), .B2(new_n341), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI211_X1 g148(.A(KEYINPUT30), .B(new_n345), .C1(new_n331), .C2(new_n341), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n320), .A2(new_n329), .A3(new_n322), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G148gat), .ZN(new_n358));
  INV_X1    g157(.A(G148gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G141gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n358), .A2(new_n360), .B1(KEYINPUT2), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n361), .ZN(new_n363));
  NOR2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT78), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G155gat), .ZN(new_n366));
  INV_X1    g165(.A(G162gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n361), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n362), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n361), .ZN(new_n372));
  XNOR2_X1  g171(.A(G141gat), .B(G148gat), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(G155gat), .B2(G162gat), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n372), .B(KEYINPUT78), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n371), .A2(new_n376), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n355), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n380), .A2(new_n329), .B1(new_n322), .B2(new_n320), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G228gat), .ZN(new_n383));
  INV_X1    g182(.A(G233gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n378), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n318), .A2(new_n319), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n329), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n379), .B1(new_n388), .B2(new_n355), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n381), .A2(new_n389), .B1(new_n383), .B2(new_n384), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G22gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT31), .B(G50gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G22gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n386), .A2(new_n397), .A3(new_n390), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(KEYINPUT82), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n386), .A2(new_n401), .A3(new_n397), .A4(new_n390), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n402), .A3(new_n392), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n403), .A2(new_n404), .A3(new_n395), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n404), .B1(new_n403), .B2(new_n395), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n353), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n377), .B2(new_n272), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n379), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n272), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n263), .A2(new_n271), .A3(KEYINPUT79), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n371), .A2(KEYINPUT3), .A3(new_n376), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n380), .A2(new_n416), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n371), .A2(KEYINPUT3), .A3(new_n376), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT3), .B1(new_n371), .B2(new_n376), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n263), .A2(KEYINPUT79), .A3(new_n271), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT79), .B1(new_n263), .B2(new_n271), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT80), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n413), .B(new_n414), .C1(new_n421), .C2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n416), .A2(new_n377), .A3(new_n417), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n273), .A2(new_n379), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n414), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n420), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n424), .A2(KEYINPUT80), .A3(new_n427), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n412), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT5), .A3(new_n414), .ZN(new_n441));
  XNOR2_X1  g240(.A(G1gat), .B(G29gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT0), .ZN(new_n443));
  XNOR2_X1  g242(.A(G57gat), .B(G85gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n437), .A2(KEYINPUT6), .A3(new_n441), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n429), .A2(new_n430), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n435), .B1(new_n440), .B2(new_n414), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n446), .A3(new_n441), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT86), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n452), .A2(new_n454), .A3(new_n457), .A4(new_n453), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n449), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n290), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n299), .B2(new_n304), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n295), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n309), .A2(new_n408), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n447), .B(KEYINPUT81), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n351), .B1(new_n465), .B2(new_n455), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n463), .A2(new_n466), .A3(new_n305), .A4(new_n407), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n407), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n466), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n458), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n331), .A2(new_n341), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n331), .B2(new_n341), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n345), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n477), .A2(KEYINPUT38), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n348), .B1(new_n477), .B2(KEYINPUT38), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n473), .A2(new_n465), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n347), .A2(new_n348), .ZN(new_n481));
  INV_X1    g280(.A(new_n350), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n481), .A2(new_n454), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT84), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n413), .B1(new_n421), .B2(new_n428), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(new_n434), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n440), .A2(KEYINPUT84), .A3(new_n414), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n445), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n485), .A3(new_n434), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT84), .B1(new_n440), .B2(new_n414), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT39), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT85), .B1(new_n494), .B2(new_n446), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n487), .A2(new_n488), .ZN(new_n496));
  INV_X1    g295(.A(new_n433), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n484), .B1(new_n497), .B2(new_n414), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n491), .A2(new_n495), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n483), .B1(new_n499), .B2(KEYINPUT40), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n491), .A2(new_n495), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n496), .A2(new_n498), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n501), .A2(KEYINPUT40), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n480), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n472), .B1(new_n504), .B2(new_n407), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n309), .A2(new_n506), .A3(new_n463), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n463), .A2(new_n305), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT36), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n469), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(new_n366), .ZN(new_n513));
  XNOR2_X1  g312(.A(G183gat), .B(G211gat), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n513), .B(new_n514), .Z(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G57gat), .B(G64gat), .Z(new_n517));
  AND2_X1   g316(.A1(G71gat), .A2(G78gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(KEYINPUT9), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n521));
  INV_X1    g320(.A(G71gat), .ZN(new_n522));
  INV_X1    g321(.A(G78gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n518), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI211_X1 g327(.A(KEYINPUT93), .B(new_n518), .C1(new_n524), .C2(new_n525), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n519), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n522), .A2(new_n523), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n517), .A2(KEYINPUT9), .A3(new_n527), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g333(.A1(G231gat), .A2(G233gat), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n251), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n533), .A2(KEYINPUT21), .ZN(new_n540));
  XOR2_X1   g339(.A(G15gat), .B(G22gat), .Z(new_n541));
  INV_X1    g340(.A(G1gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT16), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(G1gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n543), .A2(new_n546), .A3(new_n552), .A4(new_n547), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n540), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(G127gat), .B1(new_n536), .B2(new_n537), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n539), .B2(new_n556), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n516), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n556), .ZN(new_n561));
  INV_X1    g360(.A(new_n555), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n557), .A3(new_n515), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT94), .ZN(new_n567));
  AND2_X1   g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(KEYINPUT41), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT95), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT95), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT7), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n574), .A2(new_n576), .A3(G85gat), .A4(G92gat), .ZN(new_n577));
  OR2_X1    g376(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n578));
  INV_X1    g377(.A(G92gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT8), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(KEYINPUT95), .A3(new_n573), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n577), .A2(new_n581), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(G29gat), .A2(G36gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT14), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G29gat), .A2(G36gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT88), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT15), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(KEYINPUT15), .A3(new_n594), .ZN(new_n598));
  XNOR2_X1  g397(.A(G43gat), .B(G50gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n598), .A2(new_n599), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n588), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n600), .A2(new_n602), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n586), .A2(new_n587), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n586), .A2(new_n587), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n607), .A2(new_n610), .B1(KEYINPUT41), .B2(new_n568), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n572), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n570), .B1(new_n612), .B2(KEYINPUT97), .ZN(new_n613));
  INV_X1    g412(.A(new_n605), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n610), .B1(new_n614), .B2(new_n603), .ZN(new_n615));
  INV_X1    g414(.A(new_n611), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n571), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n606), .A2(new_n572), .A3(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT97), .A4(new_n570), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n565), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT98), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n565), .A2(new_n625), .A3(new_n622), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n551), .A2(new_n553), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT90), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n554), .A2(KEYINPUT90), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n630), .B(new_n631), .C1(new_n604), .C2(new_n605), .ZN(new_n632));
  NAND2_X1  g431(.A1(G229gat), .A2(G233gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT91), .Z(new_n634));
  NAND2_X1  g433(.A1(new_n628), .A2(new_n607), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT18), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n600), .A2(new_n602), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n554), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n640), .A2(new_n635), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n634), .B(KEYINPUT13), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n632), .A2(KEYINPUT18), .A3(new_n634), .A4(new_n635), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G197gat), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT11), .B(G169gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n638), .A2(new_n643), .A3(new_n650), .A4(new_n644), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G230gat), .A2(G233gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n610), .B2(new_n533), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n586), .A2(new_n587), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n609), .B1(KEYINPUT100), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n659), .A2(KEYINPUT100), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n533), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n588), .A2(KEYINPUT99), .A3(new_n530), .A4(new_n532), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n658), .A2(new_n662), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n610), .A2(new_n533), .A3(KEYINPUT10), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n656), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(KEYINPUT101), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n658), .A2(new_n662), .A3(new_n664), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n656), .ZN(new_n673));
  XOR2_X1   g472(.A(G120gat), .B(G148gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT102), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n671), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n656), .B1(new_n665), .B2(new_n666), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n673), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n627), .A2(new_n654), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n511), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n465), .A2(new_n455), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(new_n542), .ZN(G1324gat));
  INV_X1    g489(.A(new_n687), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT16), .B(G8gat), .Z(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n351), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n693), .A2(new_n694), .A3(KEYINPUT42), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT42), .B1(new_n693), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n351), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n697), .A2(KEYINPUT104), .A3(G8gat), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT104), .B1(new_n697), .B2(G8gat), .ZN(new_n699));
  OAI22_X1  g498(.A1(new_n695), .A2(new_n696), .B1(new_n698), .B2(new_n699), .ZN(G1325gat));
  AOI21_X1  g499(.A(new_n506), .B1(new_n463), .B2(new_n305), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n306), .A2(new_n308), .B1(new_n462), .B2(new_n295), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n506), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n687), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n702), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n687), .B2(new_n706), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n687), .A2(new_n407), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(new_n622), .ZN(new_n711));
  INV_X1    g510(.A(new_n654), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(new_n565), .A3(new_n684), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n511), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G29gat), .A3(new_n688), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT45), .Z(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n353), .A2(new_n407), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n459), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n702), .A2(new_n719), .B1(new_n467), .B2(KEYINPUT35), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n481), .A2(new_n454), .A3(new_n482), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n490), .B1(new_n489), .B2(new_n445), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n494), .A2(KEYINPUT85), .A3(new_n446), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n502), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT40), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n499), .A2(KEYINPUT40), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n478), .A2(new_n479), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n726), .A2(new_n727), .B1(new_n459), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n471), .B1(new_n729), .B2(new_n470), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n720), .B1(new_n730), .B2(new_n703), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n717), .B1(new_n731), .B2(new_n622), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n511), .A2(KEYINPUT44), .A3(new_n711), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n688), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n735), .A3(new_n713), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G29gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n716), .A2(new_n737), .ZN(G1328gat));
  NAND4_X1  g537(.A1(new_n732), .A2(new_n351), .A3(new_n713), .A4(new_n733), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G36gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n351), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(G36gat), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n511), .A2(new_n711), .A3(new_n713), .A4(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT105), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n740), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(G43gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n703), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n732), .A2(new_n713), .A3(new_n733), .A4(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n751), .B1(new_n714), .B2(new_n705), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1330gat));
  AOI21_X1  g558(.A(new_n407), .B1(new_n714), .B2(KEYINPUT107), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n726), .A2(new_n727), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n470), .B1(new_n761), .B2(new_n480), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n703), .B1(new_n762), .B2(new_n472), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n622), .B1(new_n763), .B2(new_n469), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(new_n765), .A3(new_n713), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(G50gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n470), .A2(G50gat), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AND4_X1   g570(.A1(new_n713), .A2(new_n732), .A3(new_n733), .A4(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n769), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(G50gat), .B1(new_n760), .B2(new_n766), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT48), .B1(new_n776), .B2(new_n772), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1331gat));
  AND3_X1   g577(.A1(new_n627), .A2(new_n712), .A3(new_n684), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n511), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n735), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G57gat), .ZN(G1332gat));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n784));
  INV_X1    g583(.A(G64gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n511), .A2(KEYINPUT108), .A3(new_n779), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT108), .B1(new_n511), .B2(new_n779), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n780), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n511), .A2(KEYINPUT108), .A3(new_n779), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n791), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n786), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n790), .A2(new_n787), .A3(new_n791), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n784), .A4(new_n785), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1333gat));
  XOR2_X1   g601(.A(new_n702), .B(KEYINPUT110), .Z(new_n803));
  NAND3_X1  g602(.A1(new_n781), .A2(new_n522), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n788), .A2(new_n789), .A3(new_n703), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n522), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n804), .B(new_n807), .C1(new_n805), .C2(new_n522), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1334gat));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n470), .ZN(new_n812));
  XNOR2_X1  g611(.A(KEYINPUT112), .B(G78gat), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n812), .B(new_n813), .ZN(G1335gat));
  NOR2_X1   g613(.A1(new_n565), .A2(new_n654), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n764), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  AND4_X1   g617(.A1(KEYINPUT51), .A2(new_n511), .A3(new_n711), .A4(new_n815), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT113), .B1(new_n816), .B2(new_n819), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n578), .A2(new_n580), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n688), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n821), .A2(new_n822), .A3(new_n684), .A4(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n685), .A2(new_n565), .A3(new_n654), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n734), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n827), .B2(new_n688), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1336gat));
  NAND4_X1  g628(.A1(new_n732), .A2(new_n351), .A3(new_n733), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G92gat), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n685), .A2(new_n741), .A3(G92gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n816), .B2(new_n819), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1337gat));
  NOR2_X1   g637(.A1(new_n705), .A2(G99gat), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n822), .A3(new_n684), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G99gat), .B1(new_n827), .B2(new_n703), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1338gat));
  NAND4_X1  g641(.A1(new_n732), .A2(new_n470), .A3(new_n733), .A4(new_n826), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(G106gat), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n407), .A2(new_n685), .A3(G106gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n816), .B2(new_n819), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n844), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1339gat));
  INV_X1    g650(.A(new_n565), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n665), .A2(new_n656), .A3(new_n666), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n669), .B2(new_n670), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n678), .B1(new_n680), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n853), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n665), .A2(KEYINPUT101), .A3(new_n666), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT101), .B1(new_n665), .B2(new_n666), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n861), .A2(new_n862), .A3(new_n656), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT55), .B(new_n858), .C1(new_n863), .C2(new_n855), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n654), .A2(new_n860), .A3(new_n679), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n640), .A2(new_n635), .A3(new_n642), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT114), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n640), .A2(new_n868), .A3(new_n635), .A4(new_n642), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n634), .B1(new_n632), .B2(new_n635), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n649), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n684), .A2(new_n653), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n711), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  AND4_X1   g673(.A1(new_n653), .A2(new_n620), .A3(new_n872), .A4(new_n621), .ZN(new_n875));
  AND4_X1   g674(.A1(new_n679), .A2(new_n875), .A3(new_n860), .A4(new_n864), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n852), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n624), .A2(new_n712), .A3(new_n626), .A4(new_n685), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n470), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n735), .A2(new_n741), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n705), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n879), .B2(new_n882), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n883), .A2(new_n884), .A3(new_n712), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n881), .B1(new_n877), .B2(new_n878), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n463), .A2(new_n305), .A3(new_n407), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n654), .A2(new_n256), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT116), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n885), .A2(new_n256), .B1(new_n889), .B2(new_n891), .ZN(G1340gat));
  NOR3_X1   g691(.A1(new_n883), .A2(new_n884), .A3(new_n685), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n684), .A2(new_n257), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n893), .A2(new_n257), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT117), .ZN(G1341gat));
  NOR3_X1   g695(.A1(new_n883), .A2(new_n884), .A3(new_n852), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n565), .A2(new_n251), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n897), .A2(new_n251), .B1(new_n889), .B2(new_n898), .ZN(G1342gat));
  NAND2_X1  g698(.A1(new_n711), .A2(new_n253), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n889), .A2(new_n900), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g700(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n901), .B(new_n902), .Z(new_n903));
  NOR3_X1   g702(.A1(new_n883), .A2(new_n884), .A3(new_n622), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n253), .B2(new_n904), .ZN(G1343gat));
  NAND3_X1  g704(.A1(new_n703), .A2(new_n735), .A3(new_n741), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n856), .B2(new_n859), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT119), .B(new_n858), .C1(new_n863), .C2(new_n855), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n908), .A2(new_n853), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n654), .A2(new_n679), .A3(new_n864), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n873), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n876), .B1(new_n912), .B2(new_n622), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT120), .B1(new_n913), .B2(new_n565), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n908), .A2(new_n853), .A3(new_n909), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n916), .A2(new_n654), .A3(new_n679), .A4(new_n864), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n711), .B1(new_n917), .B2(new_n873), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n915), .B(new_n852), .C1(new_n918), .C2(new_n876), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n914), .A2(new_n878), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n470), .A2(KEYINPUT57), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n407), .B1(new_n877), .B2(new_n878), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT57), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n906), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n357), .B1(new_n926), .B2(new_n654), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n510), .A2(KEYINPUT121), .A3(new_n407), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT121), .B1(new_n510), .B2(new_n407), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n928), .A2(new_n886), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n654), .A2(new_n357), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT122), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT58), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  AOI211_X1 g735(.A(new_n712), .B(new_n906), .C1(new_n923), .C2(new_n925), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n936), .B(new_n933), .C1(new_n937), .C2(new_n357), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(G1344gat));
  NAND3_X1  g738(.A1(new_n930), .A2(new_n359), .A3(new_n684), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT59), .B(new_n359), .C1(new_n926), .C2(new_n684), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n470), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n878), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n852), .B1(new_n918), .B2(new_n876), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n924), .A2(new_n943), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n906), .A2(new_n685), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n942), .B1(new_n952), .B2(G148gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n940), .B1(new_n941), .B2(new_n953), .ZN(G1345gat));
  AND2_X1   g753(.A1(new_n930), .A2(new_n565), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(G155gat), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n852), .A2(new_n366), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n957), .A2(new_n958), .B1(new_n926), .B2(new_n959), .ZN(G1346gat));
  AOI21_X1  g759(.A(G162gat), .B1(new_n930), .B2(new_n711), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n622), .A2(new_n367), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n926), .B2(new_n962), .ZN(G1347gat));
  NAND4_X1  g762(.A1(new_n803), .A2(new_n879), .A3(new_n688), .A4(new_n351), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(new_n203), .A3(new_n712), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n877), .A2(new_n878), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n688), .A2(new_n351), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n887), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(G169gat), .B1(new_n970), .B2(new_n654), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n965), .A2(new_n971), .ZN(G1348gat));
  OAI21_X1  g771(.A(G176gat), .B1(new_n964), .B2(new_n685), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n970), .A2(new_n204), .A3(new_n684), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1349gat));
  OAI21_X1  g774(.A(G183gat), .B1(new_n964), .B2(new_n852), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n565), .A2(new_n335), .A3(new_n332), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n969), .B2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT60), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n979), .A2(KEYINPUT125), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n978), .B(new_n980), .ZN(G1350gat));
  NAND3_X1  g780(.A1(new_n970), .A2(new_n208), .A3(new_n711), .ZN(new_n982));
  OAI21_X1  g781(.A(G190gat), .B1(new_n964), .B2(new_n622), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  OR3_X1    g785(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT126), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n510), .A2(new_n967), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(KEYINPUT127), .B1(new_n510), .B2(new_n967), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(KEYINPUT126), .B1(new_n948), .B2(new_n949), .ZN(new_n993));
  INV_X1    g792(.A(G197gat), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n712), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n987), .A2(new_n992), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n988), .A2(new_n924), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n994), .B1(new_n997), .B2(new_n712), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n996), .A2(new_n998), .ZN(G1352gat));
  NAND3_X1  g798(.A1(new_n987), .A2(new_n992), .A3(new_n993), .ZN(new_n1000));
  OAI21_X1  g799(.A(G204gat), .B1(new_n1000), .B2(new_n685), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n997), .A2(G204gat), .A3(new_n685), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1003), .ZN(G1353gat));
  NAND3_X1  g803(.A1(new_n950), .A2(new_n565), .A3(new_n992), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n565), .A2(new_n312), .ZN(new_n1008));
  OAI22_X1  g807(.A1(new_n1006), .A2(new_n1007), .B1(new_n997), .B2(new_n1008), .ZN(G1354gat));
  NOR2_X1   g808(.A1(new_n622), .A2(new_n313), .ZN(new_n1010));
  NAND4_X1  g809(.A1(new_n987), .A2(new_n992), .A3(new_n993), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n313), .B1(new_n997), .B2(new_n622), .ZN(new_n1012));
  AND2_X1   g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1355gat));
endmodule


