//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  AOI21_X1  g001(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT18), .A3(G131), .ZN(new_n192));
  XNOR2_X1  g006(.A(G125), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT18), .A2(G131), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n189), .A2(new_n190), .A3(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n190), .ZN(new_n199));
  OAI21_X1  g013(.A(G131), .B1(new_n199), .B2(new_n188), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n189), .A2(new_n201), .A3(new_n190), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT75), .B1(new_n193), .B2(KEYINPUT16), .ZN(new_n208));
  OAI211_X1 g022(.A(G146), .B(new_n207), .C1(new_n208), .C2(new_n205), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n193), .A2(KEYINPUT19), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n193), .A2(KEYINPUT19), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n194), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n203), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n209), .A2(new_n214), .A3(new_n212), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n198), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G113), .B(G122), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n200), .A2(new_n202), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G140), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G125), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n204), .A2(G140), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT16), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n205), .B1(new_n227), .B2(new_n206), .ZN(new_n228));
  INV_X1    g042(.A(new_n207), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n194), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n191), .A2(KEYINPUT17), .A3(G131), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n223), .A2(new_n230), .A3(new_n209), .A4(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n220), .A3(new_n198), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT90), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n232), .A2(new_n235), .A3(new_n220), .A4(new_n198), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n217), .A2(new_n221), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(G475), .A2(G902), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT20), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n236), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n214), .B1(new_n209), .B2(new_n212), .ZN(new_n242));
  INV_X1    g056(.A(new_n203), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n216), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n198), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n221), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT20), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n238), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n232), .A2(new_n198), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n221), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n241), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G902), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT91), .B(G475), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n240), .A2(new_n249), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G478), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT15), .ZN(new_n258));
  INV_X1    g072(.A(G122), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G116), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G122), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT92), .ZN(new_n264));
  XNOR2_X1  g078(.A(G116), .B(G122), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT92), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G107), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n264), .A2(new_n267), .A3(G107), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT93), .ZN(new_n273));
  INV_X1    g087(.A(G143), .ZN(new_n274));
  OAI22_X1  g088(.A1(new_n273), .A2(KEYINPUT13), .B1(new_n274), .B2(G128), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT13), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(KEYINPUT93), .ZN(new_n277));
  OAI21_X1  g091(.A(G134), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(G128), .B(G143), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n279), .B(G134), .C1(new_n275), .C2(new_n277), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n272), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n261), .A2(KEYINPUT14), .A3(G122), .ZN(new_n285));
  OAI211_X1 g099(.A(G107), .B(new_n285), .C1(new_n263), .C2(KEYINPUT14), .ZN(new_n286));
  INV_X1    g100(.A(G134), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n279), .A2(G134), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G107), .B1(new_n264), .B2(new_n267), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT9), .B(G234), .ZN(new_n293));
  INV_X1    g107(.A(G217), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(new_n294), .A3(G953), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n284), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n270), .A2(new_n271), .B1(new_n282), .B2(new_n281), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n290), .A2(new_n291), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n258), .B1(new_n301), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n258), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n297), .A2(new_n300), .A3(new_n253), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(KEYINPUT94), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(G234), .A2(G237), .ZN(new_n310));
  INV_X1    g124(.A(G953), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n310), .A2(G952), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT21), .B(G898), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT95), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n310), .A2(G902), .A3(G953), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n256), .A2(new_n309), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G122), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n269), .A3(G104), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n219), .A2(G107), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G101), .ZN(new_n327));
  INV_X1    g141(.A(G101), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n322), .A2(new_n324), .A3(new_n328), .A4(new_n325), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(KEYINPUT4), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G116), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n261), .A2(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT2), .B(G113), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT69), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n335), .ZN(new_n337));
  INV_X1    g151(.A(G113), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT2), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G113), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G116), .B(G119), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n326), .A2(new_n347), .A3(G101), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n330), .A2(new_n336), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n325), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n219), .A2(G107), .ZN(new_n351));
  OAI21_X1  g165(.A(G101), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(new_n329), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n261), .A2(G119), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT5), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n338), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n354), .A2(new_n357), .B1(new_n343), .B2(new_n342), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n321), .B1(new_n349), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT6), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n349), .A2(new_n359), .A3(new_n321), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT84), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT84), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n349), .A2(new_n365), .A3(new_n359), .A4(new_n321), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n361), .B1(new_n367), .B2(new_n360), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n274), .A2(G146), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT64), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n194), .B2(G143), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n274), .A2(KEYINPUT64), .A3(G146), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G128), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n194), .A2(G143), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(KEYINPUT1), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT65), .B1(new_n194), .B2(G143), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT65), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n274), .A3(G146), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n369), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT1), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G128), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n379), .A2(new_n385), .A3(new_n204), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(KEYINPUT0), .A2(G128), .ZN(new_n388));
  NOR2_X1   g202(.A1(KEYINPUT0), .A2(G128), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n374), .A2(new_n390), .B1(new_n383), .B2(new_n388), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n204), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n311), .A2(G224), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n368), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G210), .B1(G237), .B2(G902), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(KEYINPUT7), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n387), .B2(new_n392), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n386), .B(new_n400), .C1(new_n204), .C2(new_n391), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n366), .B2(new_n364), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n354), .A2(new_n357), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n344), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n352), .A2(new_n329), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n407), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n353), .A2(new_n358), .A3(KEYINPUT86), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n321), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(KEYINPUT87), .A3(new_n413), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(G902), .B1(new_n403), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n396), .A2(new_n397), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n397), .B1(new_n396), .B2(new_n419), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G214), .B1(G237), .B2(G902), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT88), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n427), .B(new_n424), .C1(new_n421), .C2(new_n422), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n320), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(KEYINPUT68), .A2(G137), .ZN(new_n432));
  NOR2_X1   g246(.A1(KEYINPUT68), .A2(G137), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT11), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(new_n287), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n434), .A2(new_n436), .B1(new_n287), .B2(G137), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT67), .ZN(new_n438));
  INV_X1    g252(.A(G137), .ZN(new_n439));
  AOI22_X1  g253(.A1(KEYINPUT66), .A2(new_n435), .B1(new_n439), .B2(G134), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT66), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT11), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n438), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(G134), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(KEYINPUT66), .ZN(new_n445));
  AND4_X1   g259(.A1(new_n438), .A2(new_n442), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n437), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G131), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n437), .B(new_n201), .C1(new_n443), .C2(new_n446), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT80), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n381), .B1(new_n274), .B2(G146), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n194), .A2(KEYINPUT65), .A3(G143), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n376), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n384), .A2(G128), .ZN(new_n455));
  OAI22_X1  g269(.A1(new_n454), .A2(new_n455), .B1(new_n373), .B2(new_n377), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n451), .B1(new_n456), .B2(new_n353), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n379), .A2(new_n385), .A3(KEYINPUT80), .A4(new_n407), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI211_X1 g273(.A(new_n455), .B(new_n369), .C1(new_n380), .C2(new_n382), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n378), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT79), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n378), .A3(KEYINPUT79), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n407), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n450), .B1(new_n459), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n462), .B1(new_n383), .B2(new_n377), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n469), .A3(new_n385), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n353), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n457), .A3(new_n458), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT12), .A3(new_n450), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(KEYINPUT81), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G140), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n311), .A2(G227), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n456), .A2(new_n353), .A3(KEYINPUT10), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n330), .A2(new_n348), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n374), .A2(new_n390), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n383), .A2(new_n388), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n479), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT10), .B1(new_n470), .B2(new_n353), .ZN(new_n485));
  OR3_X1    g299(.A1(new_n484), .A2(new_n485), .A3(new_n450), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT81), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n466), .A2(new_n487), .A3(new_n467), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n474), .A2(new_n478), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n450), .B1(new_n484), .B2(new_n485), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n490), .B1(new_n492), .B2(new_n477), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G469), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n488), .A2(new_n486), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n496), .A2(new_n490), .A3(new_n478), .A4(new_n474), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n253), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(G469), .A2(G902), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT82), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n473), .A2(KEYINPUT81), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT12), .B1(new_n472), .B2(new_n450), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n488), .A2(new_n486), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n474), .A2(KEYINPUT82), .A3(new_n486), .A4(new_n488), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n477), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n492), .A2(new_n477), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(G469), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n431), .B1(new_n500), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n429), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n294), .B1(G234), .B2(new_n253), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT74), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n311), .A2(G221), .A3(G234), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n230), .A2(new_n209), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n375), .A2(G119), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT23), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n375), .A2(KEYINPUT23), .A3(G119), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n331), .A2(G128), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G110), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n520), .A2(new_n524), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT24), .B(G110), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G110), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n522), .A2(new_n523), .A3(new_n532), .A4(new_n524), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n528), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n533), .A2(new_n534), .B1(new_n194), .B2(new_n193), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n519), .A2(new_n531), .B1(new_n209), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n518), .B1(new_n536), .B2(KEYINPUT76), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n519), .A2(new_n531), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n209), .A2(new_n535), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(KEYINPUT76), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT76), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n530), .B1(new_n230), .B2(new_n209), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n209), .A2(new_n535), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n537), .B1(new_n545), .B2(new_n518), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT25), .B1(new_n546), .B2(new_n253), .ZN(new_n547));
  INV_X1    g361(.A(new_n518), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n540), .B2(new_n544), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n550));
  NOR4_X1   g364(.A1(new_n549), .A2(new_n537), .A3(new_n550), .A4(G902), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n515), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT77), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT77), .B(new_n515), .C1(new_n547), .C2(new_n551), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n514), .A2(G902), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n556), .B(KEYINPUT78), .Z(new_n557));
  NAND2_X1  g371(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n346), .A2(new_n336), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n483), .B1(new_n448), .B2(new_n449), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n444), .B1(new_n434), .B2(G134), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G131), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n449), .A2(new_n566), .A3(new_n456), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n564), .A2(new_n567), .A3(KEYINPUT30), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n569));
  INV_X1    g383(.A(new_n449), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n441), .A2(KEYINPUT11), .B1(new_n287), .B2(G137), .ZN(new_n571));
  INV_X1    g385(.A(new_n442), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT67), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n440), .A2(new_n438), .A3(new_n442), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n201), .B1(new_n575), .B2(new_n437), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n391), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n449), .A2(new_n566), .A3(new_n456), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n563), .B1(new_n568), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n346), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT70), .B1(new_n346), .B2(new_n336), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n577), .A2(new_n583), .A3(new_n578), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n585));
  NAND2_X1  g399(.A1(new_n187), .A2(G210), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT26), .B(G101), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(new_n584), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT31), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n584), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT30), .B1(new_n564), .B2(new_n567), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n577), .A2(new_n569), .A3(new_n578), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n594), .B1(new_n597), .B2(new_n563), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(KEYINPUT31), .A3(new_n590), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n563), .B1(new_n564), .B2(new_n567), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n584), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT28), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT28), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n584), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT72), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n584), .A2(KEYINPUT72), .A3(new_n604), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n603), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n589), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n561), .B1(new_n600), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n608), .ZN(new_n612));
  OAI22_X1  g426(.A1(new_n564), .A2(new_n567), .B1(new_n581), .B2(new_n582), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n604), .B1(new_n613), .B2(new_n584), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT72), .B1(new_n584), .B2(new_n604), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT29), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n589), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT73), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n598), .B2(new_n590), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n562), .B1(new_n595), .B2(new_n596), .ZN(new_n622));
  OAI211_X1 g436(.A(KEYINPUT73), .B(new_n589), .C1(new_n622), .C2(new_n594), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n603), .A2(new_n607), .A3(new_n608), .A4(new_n590), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n617), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n619), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AOI22_X1  g441(.A1(KEYINPUT32), .A2(new_n611), .B1(new_n627), .B2(G472), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT32), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n593), .A2(new_n599), .B1(new_n609), .B2(new_n589), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n561), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n559), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n513), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n328), .ZN(G3));
  NAND2_X1  g449(.A1(new_n396), .A2(new_n419), .ZN(new_n636));
  INV_X1    g450(.A(new_n397), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n420), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n396), .A2(new_n419), .A3(KEYINPUT96), .A4(new_n397), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(new_n424), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n234), .A2(new_n236), .B1(new_n221), .B2(new_n250), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n255), .B1(new_n644), .B2(G902), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n248), .B1(new_n247), .B2(new_n238), .ZN(new_n646));
  AOI211_X1 g460(.A(KEYINPUT20), .B(new_n239), .C1(new_n241), .C2(new_n246), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n257), .B1(new_n301), .B2(G902), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n297), .A2(new_n300), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n284), .A2(new_n292), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n652), .B1(new_n653), .B2(KEYINPUT98), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n296), .B2(KEYINPUT99), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n654), .A2(new_n296), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n651), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n253), .A2(G478), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n649), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n648), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n643), .A2(new_n317), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n630), .B2(G902), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT31), .B1(new_n598), .B2(new_n590), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n622), .A2(new_n592), .A3(new_n594), .A4(new_n589), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n604), .B1(new_n601), .B2(new_n584), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n612), .A2(new_n667), .A3(new_n615), .ZN(new_n668));
  OAI22_X1  g482(.A1(new_n665), .A2(new_n666), .B1(new_n668), .B2(new_n590), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n560), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n559), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n663), .A2(new_n672), .A3(new_n512), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT34), .B(G104), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n646), .B2(new_n647), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n240), .A2(new_n249), .A3(KEYINPUT100), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n307), .A2(new_n645), .A3(new_n308), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n318), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n643), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n672), .A3(new_n512), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G107), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G9));
  NOR2_X1   g500(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n536), .B(new_n687), .Z(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n557), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n554), .A2(new_n555), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n513), .A2(new_n671), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT37), .B(G110), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  INV_X1    g508(.A(G900), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n312), .B1(new_n316), .B2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n678), .A2(new_n680), .A3(new_n677), .A4(new_n697), .ZN(new_n698));
  AND4_X1   g512(.A1(new_n640), .A2(new_n698), .A3(new_n642), .A4(new_n690), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n627), .A2(G472), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n669), .A2(KEYINPUT32), .A3(new_n560), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n631), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n699), .A2(new_n702), .A3(new_n512), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  XOR2_X1   g518(.A(new_n696), .B(KEYINPUT39), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n512), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n690), .A2(new_n425), .A3(new_n256), .A4(new_n309), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n423), .B(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n598), .A2(new_n589), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n613), .A2(new_n584), .A3(new_n589), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n253), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n631), .A2(new_n701), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n709), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n707), .A2(new_n708), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  AND3_X1   g533(.A1(new_n648), .A2(new_n661), .A3(new_n697), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n640), .A2(new_n690), .A3(new_n720), .A4(new_n642), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n702), .A3(new_n512), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  NAND3_X1  g537(.A1(new_n494), .A2(new_n253), .A3(new_n497), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n430), .A3(new_n498), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n633), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n663), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT103), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n728), .B(new_n730), .ZN(G15));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n682), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  AND2_X1   g547(.A1(new_n690), .A2(new_n319), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n725), .A2(new_n430), .A3(new_n498), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n640), .A2(new_n642), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n735), .A3(new_n702), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  INV_X1    g552(.A(G472), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n669), .B2(new_n253), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n607), .A2(new_n608), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n589), .B1(new_n741), .B2(new_n614), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n561), .B1(new_n600), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n559), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n256), .A2(new_n309), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n640), .A2(new_n745), .A3(new_n642), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n735), .A3(new_n746), .A4(new_n318), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NOR2_X1   g562(.A1(new_n726), .A2(new_n643), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n740), .A2(new_n743), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n751), .B2(new_n690), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n600), .A2(new_n742), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n560), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n750), .A2(new_n690), .A3(new_n664), .A4(new_n754), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n720), .B(new_n749), .C1(new_n752), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n631), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n670), .A2(KEYINPUT108), .A3(new_n629), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n701), .A3(new_n760), .A4(new_n700), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n638), .A2(new_n430), .A3(new_n424), .A4(new_n420), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n508), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n506), .A2(KEYINPUT106), .A3(new_n507), .A4(new_n477), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n509), .B(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(G469), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n499), .B(KEYINPUT105), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n498), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n762), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n559), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n761), .A2(new_n772), .A3(new_n773), .A4(new_n720), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT42), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  INV_X1    g590(.A(new_n720), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT42), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n632), .A2(new_n772), .A3(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n775), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G131), .ZN(G33));
  NAND3_X1  g597(.A1(new_n632), .A2(new_n698), .A3(new_n772), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  AOI21_X1  g599(.A(KEYINPUT43), .B1(new_n256), .B2(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n256), .A2(new_n661), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n671), .A3(new_n690), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n508), .B2(new_n510), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n495), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n764), .A2(KEYINPUT45), .A3(new_n765), .A4(new_n767), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n770), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n498), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n431), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n423), .A2(new_n424), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n789), .B2(new_n790), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n794), .A2(new_n705), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  OAI221_X1 g624(.A(new_n430), .B1(KEYINPUT112), .B2(new_n810), .C1(new_n802), .C2(new_n803), .ZN(new_n811));
  XNOR2_X1  g625(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n805), .B2(new_n812), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n702), .A2(new_n773), .A3(new_n777), .A4(new_n806), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n813), .A2(KEYINPUT113), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT113), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NAND2_X1  g633(.A1(new_n725), .A2(new_n498), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT114), .Z(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT49), .Z(new_n822));
  OR4_X1    g636(.A1(new_n559), .A2(new_n431), .A3(new_n425), .A4(new_n787), .ZN(new_n823));
  OR4_X1    g637(.A1(new_n711), .A2(new_n822), .A3(new_n716), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n821), .A2(new_n431), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT119), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n802), .A2(new_n803), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n812), .B1(new_n828), .B2(new_n430), .ZN(new_n829));
  INV_X1    g643(.A(new_n811), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n788), .A2(new_n312), .A3(new_n744), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n806), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n832), .A2(new_n424), .A3(new_n711), .A4(new_n726), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT50), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n752), .A2(new_n755), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n726), .A2(new_n806), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n838), .A2(new_n788), .A3(new_n312), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n773), .A2(new_n312), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n840), .A2(new_n716), .A3(new_n726), .A4(new_n806), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n648), .A2(new_n661), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n837), .A2(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT51), .B1(new_n834), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n761), .A2(new_n773), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n839), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT48), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT48), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n839), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n749), .ZN(new_n853));
  OAI211_X1 g667(.A(G952), .B(new_n311), .C1(new_n832), .C2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n662), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n855), .B2(new_n841), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n852), .A2(new_n856), .A3(KEYINPUT120), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n833), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n813), .B2(new_n826), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n836), .A2(KEYINPUT51), .A3(new_n843), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n825), .B1(new_n846), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n864), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n813), .A2(new_n826), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n868), .B2(new_n862), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n862), .B1(new_n813), .B2(new_n827), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(new_n844), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n872), .A3(KEYINPUT121), .A4(new_n861), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n747), .A2(new_n737), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n632), .B(new_n735), .C1(new_n663), .C2(new_n682), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n256), .A2(new_n305), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n662), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n317), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n426), .A2(new_n428), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n672), .A3(new_n881), .A4(new_n512), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n671), .A2(new_n691), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n512), .B(new_n429), .C1(new_n632), .C2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n875), .A2(new_n876), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n720), .B(new_n772), .C1(new_n752), .C2(new_n755), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n305), .A2(new_n696), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n645), .A2(new_n690), .A3(new_n679), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n762), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n500), .A2(new_n511), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n888), .A2(new_n889), .A3(new_n702), .A4(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n784), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n886), .A2(new_n784), .A3(KEYINPUT115), .A4(new_n891), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n885), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n896), .A2(new_n782), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n702), .B(new_n512), .C1(new_n699), .C2(new_n721), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n690), .A2(new_n431), .A3(new_n696), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n768), .A2(new_n771), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n716), .A4(new_n746), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n756), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n899), .A2(new_n756), .A3(KEYINPUT52), .A4(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT53), .A4(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n909));
  NOR2_X1   g723(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n756), .A2(new_n899), .A3(new_n902), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n903), .B2(new_n909), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n782), .A3(new_n896), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT117), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n896), .A2(new_n782), .A3(new_n907), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n908), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT54), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n915), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n775), .A2(KEYINPUT53), .A3(new_n779), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n913), .A2(new_n896), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(KEYINPUT118), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n919), .A2(new_n928), .A3(KEYINPUT54), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n874), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(G952), .A2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n824), .B1(new_n930), .B2(new_n931), .ZN(G75));
  AND2_X1   g746(.A1(new_n921), .A2(new_n924), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n253), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(G210), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n368), .B(new_n395), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT55), .Z(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n311), .A2(G952), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(G51));
  NOR3_X1   g757(.A1(new_n933), .A2(new_n253), .A3(new_n798), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n494), .A2(new_n497), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n921), .A2(new_n924), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT54), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n925), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n769), .B(KEYINPUT57), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n944), .B1(new_n950), .B2(KEYINPUT123), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  INV_X1    g766(.A(new_n949), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n947), .B2(new_n925), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(new_n954), .B2(new_n945), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n942), .B1(new_n951), .B2(new_n955), .ZN(G54));
  AND2_X1   g770(.A1(KEYINPUT58), .A2(G475), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n934), .A2(new_n247), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n247), .B1(new_n934), .B2(new_n957), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n942), .ZN(G60));
  INV_X1    g774(.A(new_n942), .ZN(new_n961));
  INV_X1    g775(.A(new_n948), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n659), .B(KEYINPUT124), .Z(new_n963));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT59), .Z(new_n965));
  OR2_X1    g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n961), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n965), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n927), .A2(new_n929), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n967), .B1(new_n969), .B2(new_n963), .ZN(G63));
  XOR2_X1   g784(.A(new_n546), .B(KEYINPUT125), .Z(new_n971));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT60), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n933), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n946), .A2(new_n688), .A3(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n974), .A2(new_n961), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g792(.A(G224), .ZN(new_n979));
  OAI21_X1  g793(.A(G953), .B1(new_n315), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n885), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(G953), .ZN(new_n982));
  INV_X1    g796(.A(new_n368), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(G898), .B2(new_n311), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  NOR2_X1   g799(.A1(new_n210), .A2(new_n211), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n597), .B(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(G900), .B2(G953), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n899), .A2(new_n756), .A3(new_n784), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n808), .A2(new_n782), .A3(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n805), .A2(new_n705), .A3(new_n746), .A4(new_n847), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n818), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n988), .B1(new_n992), .B2(G953), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n718), .A2(new_n756), .A3(new_n899), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  OR4_X1    g810(.A1(new_n633), .A2(new_n706), .A3(new_n806), .A4(new_n879), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n996), .A2(new_n808), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n816), .B2(new_n817), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n987), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n311), .B1(G227), .B2(G900), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT126), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n993), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n993), .B2(new_n1000), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(G72));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT127), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n992), .B2(new_n885), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1009), .A2(new_n589), .A3(new_n598), .ZN(new_n1010));
  INV_X1    g824(.A(new_n998), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n818), .A2(new_n1011), .A3(new_n981), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n1008), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n942), .B1(new_n1013), .B2(new_n712), .ZN(new_n1014));
  INV_X1    g828(.A(new_n591), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n919), .B(new_n1007), .C1(new_n1015), .C2(new_n624), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1010), .A2(new_n1014), .A3(new_n1016), .ZN(G57));
endmodule


