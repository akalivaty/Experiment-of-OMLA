//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n446, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  XOR2_X1   g035(.A(G325), .B(KEYINPUT67), .Z(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  OR2_X1    g047(.A1(new_n467), .A2(new_n468), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n463), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n469), .A2(new_n463), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n463), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n473), .A2(new_n463), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n479), .B1(new_n480), .B2(new_n481), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n482), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n470), .A2(KEYINPUT4), .A3(G138), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n478), .A2(G126), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT71), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(new_n500), .A3(KEYINPUT5), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n509), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND2_X1  g090(.A1(new_n503), .A2(new_n505), .ZN(new_n516));
  INV_X1    g091(.A(new_n501), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n516), .A2(new_n517), .A3(new_n511), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n519));
  AND3_X1   g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n518), .A2(G89), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(KEYINPUT72), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n527), .A2(new_n531), .A3(G51), .A4(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(KEYINPUT73), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n524), .B2(new_n532), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n523), .B1(new_n534), .B2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND4_X1  g113(.A1(new_n527), .A2(new_n531), .A3(G52), .A4(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n506), .A2(new_n511), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n506), .A2(G64), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n508), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  AND3_X1   g121(.A1(new_n516), .A2(G56), .A3(new_n517), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n527), .A2(new_n531), .A3(G43), .A4(G543), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n516), .A2(G81), .A3(new_n517), .A4(new_n511), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n553), .A3(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  AND2_X1   g133(.A1(KEYINPUT75), .A2(G65), .ZN(new_n559));
  NOR2_X1   g134(.A1(KEYINPUT75), .A2(G65), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n504), .B1(KEYINPUT5), .B2(new_n500), .ZN(new_n562));
  NOR3_X1   g137(.A1(new_n502), .A2(KEYINPUT71), .A3(G543), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n561), .B(new_n517), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n518), .B2(G91), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n527), .A2(new_n531), .A3(G53), .A4(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n500), .B1(new_n511), .B2(new_n528), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n570), .A2(new_n571), .A3(G53), .A4(new_n527), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n567), .A2(KEYINPUT76), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT76), .B1(new_n567), .B2(new_n573), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  NAND2_X1  g152(.A1(new_n518), .A2(G87), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n527), .A2(new_n531), .A3(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n506), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n583), .A2(new_n508), .B1(new_n584), .B2(new_n512), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n579), .A2(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n540), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n508), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n579), .A2(KEYINPUT78), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n579), .A2(KEYINPUT78), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n598), .A2(G54), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n518), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n540), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n508), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n600), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  AOI21_X1  g191(.A(new_n549), .B1(new_n506), .B2(G56), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n551), .B(new_n552), .C1(new_n617), .C2(new_n508), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n600), .A2(new_n605), .A3(new_n607), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(G559), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT79), .ZN(new_n621));
  MUX2_X1   g196(.A(new_n618), .B(new_n621), .S(G868), .Z(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n465), .A2(new_n473), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n478), .A2(G123), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n463), .A2(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G135), .ZN(new_n634));
  OAI221_X1 g209(.A(new_n631), .B1(new_n632), .B2(new_n633), .C1(new_n485), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n647), .A2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NOR2_X1   g230(.A1(G2072), .A2(G2078), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n445), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n658), .B2(KEYINPUT82), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(KEYINPUT82), .B2(new_n658), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n657), .B(KEYINPUT17), .ZN(new_n663));
  INV_X1    g238(.A(new_n655), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n660), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n662), .A2(new_n657), .A3(new_n664), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n664), .A3(new_n661), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n677), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT20), .Z(new_n681));
  AOI211_X1 g256(.A(new_n679), .B(new_n681), .C1(new_n674), .C2(new_n678), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G35), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT94), .Z(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n489), .B2(G29), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT29), .ZN(new_n693));
  INV_X1    g268(.A(G2090), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G29), .A2(G33), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n698));
  NAND3_X1  g273(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G139), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n485), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n463), .B1(new_n706), .B2(KEYINPUT90), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(KEYINPUT90), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n697), .B1(new_n709), .B2(new_n689), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(new_n443), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n695), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n689), .A2(G32), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n478), .A2(G129), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT26), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n465), .A2(G105), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n485), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G141), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n713), .B1(new_n721), .B2(new_n689), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n689), .A2(G26), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT28), .Z(new_n726));
  OR2_X1    g301(.A1(G104), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT86), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G128), .B2(new_n478), .ZN(new_n730));
  INV_X1    g305(.A(G140), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n485), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n726), .B1(new_n732), .B2(G29), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2067), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(G19), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n618), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G1341), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n724), .A2(new_n734), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT31), .B(G11), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT92), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(G28), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n689), .B1(new_n744), .B2(G28), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n743), .B1(new_n745), .B2(new_n746), .C1(new_n635), .C2(new_n689), .ZN(new_n747));
  NAND2_X1  g322(.A1(G160), .A2(G29), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G34), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(new_n689), .ZN(new_n751));
  AOI21_X1  g326(.A(G2084), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n748), .A2(G2084), .A3(new_n751), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n747), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n735), .A2(G5), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G171), .B2(new_n735), .ZN(new_n756));
  INV_X1    g331(.A(G1961), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n689), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n689), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(new_n444), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n754), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n741), .B(new_n762), .C1(new_n693), .C2(new_n694), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n735), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n735), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(G1966), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT93), .Z(new_n767));
  NAND2_X1  g342(.A1(G299), .A2(G16), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n735), .A2(G20), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT23), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1956), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n608), .A2(new_n735), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G4), .B2(new_n735), .ZN(new_n774));
  INV_X1    g349(.A(G1348), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n765), .A2(G1966), .ZN(new_n778));
  NOR4_X1   g353(.A1(new_n772), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n712), .A2(new_n763), .A3(new_n767), .A4(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G23), .B(G288), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT33), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1976), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n735), .A2(G6), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n588), .B2(new_n735), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT32), .B(G1981), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT84), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n785), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n735), .A2(G22), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT85), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n735), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1971), .Z(new_n793));
  NAND4_X1  g368(.A1(new_n783), .A2(new_n788), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n689), .A2(G25), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n720), .A2(G131), .ZN(new_n798));
  NOR2_X1   g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT83), .Z(new_n800));
  INV_X1    g375(.A(G2104), .ZN(new_n801));
  INV_X1    g376(.A(G107), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G2105), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n800), .A2(new_n803), .B1(new_n478), .B2(G119), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n797), .B1(new_n806), .B2(new_n689), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G1986), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n595), .A2(new_n735), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n735), .B2(G24), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n810), .B2(new_n812), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n795), .A2(new_n796), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT36), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n795), .A2(new_n817), .A3(new_n796), .A4(new_n814), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n780), .B1(new_n816), .B2(new_n818), .ZN(G311));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n820));
  XNOR2_X1  g395(.A(G311), .B(new_n820), .ZN(G150));
  NAND4_X1  g396(.A1(new_n527), .A2(new_n531), .A3(G55), .A4(G543), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n516), .A2(G93), .A3(new_n517), .A4(new_n511), .ZN(new_n823));
  NAND2_X1  g398(.A1(G80), .A2(G543), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n506), .B2(G67), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n822), .B(new_n823), .C1(new_n826), .C2(new_n508), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G860), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n608), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT96), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT38), .Z(new_n834));
  AND2_X1   g409(.A1(new_n618), .A2(new_n827), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n618), .A2(new_n827), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n834), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n831), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(new_n837), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n834), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n830), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(new_n635), .B(G160), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n489), .B(new_n847), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n704), .A2(new_n850), .A3(new_n708), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  INV_X1    g427(.A(G118), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(G2105), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n720), .A2(G142), .ZN(new_n855));
  AOI211_X1 g430(.A(new_n854), .B(new_n855), .C1(G130), .C2(new_n478), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n709), .A2(KEYINPUT99), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n732), .B(G164), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n721), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n732), .B(new_n498), .ZN(new_n863));
  INV_X1    g438(.A(new_n721), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n860), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n859), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n805), .B(new_n626), .Z(new_n868));
  AND2_X1   g443(.A1(new_n862), .A2(new_n865), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n869), .A2(new_n857), .A3(new_n860), .A4(new_n858), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT101), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n868), .B1(new_n867), .B2(new_n870), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n849), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n875), .A2(KEYINPUT101), .A3(new_n848), .A4(new_n871), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(KEYINPUT100), .B(G37), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g455(.A1(new_n827), .A2(new_n611), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n621), .B(new_n840), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n574), .B2(new_n575), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT76), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n569), .A2(new_n572), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n506), .A2(new_n561), .B1(G78), .B2(G543), .ZN(new_n887));
  INV_X1    g462(.A(G91), .ZN(new_n888));
  OAI22_X1  g463(.A1(new_n887), .A2(new_n508), .B1(new_n888), .B2(new_n540), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n567), .A2(KEYINPUT76), .A3(new_n573), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(KEYINPUT102), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n608), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n619), .A2(new_n890), .A3(KEYINPUT102), .A4(new_n891), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n882), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT103), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n898), .A3(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n893), .A2(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT41), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n882), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G303), .B(G288), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n588), .A2(new_n595), .ZN(new_n906));
  AOI21_X1  g481(.A(G290), .B1(new_n586), .B2(new_n587), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(G305), .A2(G290), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n588), .A2(new_n595), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n910), .A3(new_n904), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT42), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n903), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n881), .B1(new_n914), .B2(new_n611), .ZN(G295));
  OAI21_X1  g490(.A(new_n881), .B1(new_n914), .B2(new_n611), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  NAND2_X1  g492(.A1(G171), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n533), .B(KEYINPUT73), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n523), .ZN(new_n920));
  INV_X1    g495(.A(G67), .ZN(new_n921));
  AOI211_X1 g496(.A(new_n921), .B(new_n501), .C1(new_n503), .C2(new_n505), .ZN(new_n922));
  OAI21_X1  g497(.A(G651), .B1(new_n922), .B2(new_n825), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n822), .A2(new_n823), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n550), .A2(new_n553), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n617), .A2(new_n508), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n551), .A2(new_n552), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n516), .A2(G67), .A3(new_n517), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n508), .B1(new_n928), .B2(new_n824), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n822), .A2(new_n823), .ZN(new_n930));
  OAI22_X1  g505(.A1(new_n926), .A2(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT105), .B1(new_n542), .B2(new_n545), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n925), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n925), .B2(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n920), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n932), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n835), .B2(new_n836), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n542), .A2(new_n545), .A3(KEYINPUT105), .ZN(new_n938));
  NOR2_X1   g513(.A1(G286), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n925), .A2(new_n931), .A3(new_n932), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n893), .A2(new_n898), .A3(new_n894), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n898), .B1(new_n893), .B2(new_n894), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n893), .A2(new_n935), .A3(new_n941), .A4(new_n894), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n935), .A2(new_n941), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n895), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n945), .A2(new_n912), .A3(new_n947), .A4(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n946), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n901), .A2(KEYINPUT108), .A3(new_n899), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n944), .A2(new_n954), .B1(new_n941), .B2(new_n935), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n878), .B(new_n951), .C1(new_n956), .C2(new_n912), .ZN(new_n957));
  XOR2_X1   g532(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n946), .B(new_n949), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n912), .B1(new_n962), .B2(new_n945), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n963), .B2(G37), .ZN(new_n964));
  INV_X1    g539(.A(G37), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n950), .A2(new_n947), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n948), .B1(new_n901), .B2(new_n899), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT107), .B(new_n965), .C1(new_n968), .C2(new_n912), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n951), .A3(new_n969), .ZN(new_n970));
  AOI211_X1 g545(.A(KEYINPUT44), .B(new_n960), .C1(new_n970), .C2(new_n959), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n964), .A2(new_n969), .A3(new_n958), .A4(new_n951), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT109), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n970), .A2(new_n959), .ZN(new_n977));
  INV_X1    g552(.A(new_n960), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n972), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(new_n974), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT44), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n976), .A2(new_n983), .ZN(G397));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n498), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G160), .A2(G40), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(G1996), .A3(new_n864), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT110), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n732), .B(G2067), .Z(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G1996), .B2(new_n864), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n806), .A2(new_n808), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n806), .A2(new_n808), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n989), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n595), .B(new_n810), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n989), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n498), .A2(new_n985), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n498), .B2(new_n985), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n988), .ZN(new_n1007));
  INV_X1    g582(.A(G2084), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n986), .A2(new_n988), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1966), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n1013), .B2(G168), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G286), .A2(G8), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT124), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT123), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1012), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT123), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1014), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1013), .A2(new_n1026), .A3(new_n1015), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1001), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1023), .B2(G286), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1016), .B1(new_n1023), .B2(KEYINPUT123), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(KEYINPUT62), .A3(new_n1027), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n757), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n444), .A4(new_n1011), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1036), .A2(KEYINPUT125), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT125), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n987), .A2(new_n1042), .A3(new_n1011), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1003), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n988), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1041), .B1(new_n1047), .B2(G2078), .ZN(new_n1048));
  AOI21_X1  g623(.A(G301), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1029), .A2(new_n1034), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n988), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n1051), .A2(G1971), .B1(G2090), .B2(new_n1035), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G303), .A2(G8), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1055), .A2(KEYINPUT112), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT112), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1052), .A2(G8), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1052), .A2(new_n1059), .A3(KEYINPUT113), .A4(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n988), .A2(new_n1002), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n1020), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(G288), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT52), .B(new_n1068), .C1(new_n1067), .C2(G288), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n585), .B(G1981), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1020), .B(new_n1065), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1068), .A2(KEYINPUT52), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1069), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1007), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT116), .B1(new_n1006), .B2(new_n988), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1005), .ZN(new_n1080));
  OAI22_X1  g655(.A1(G1971), .A2(new_n1051), .B1(new_n1080), .B2(G2090), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1064), .A2(new_n1076), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT127), .B1(new_n1050), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  OR3_X1    g662(.A1(new_n1013), .A2(KEYINPUT117), .A3(G286), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT117), .B1(new_n1013), .B2(G286), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1052), .A2(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1083), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1064), .A2(new_n1092), .A3(new_n1076), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1064), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n585), .A2(G1981), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT114), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G288), .A2(G1976), .ZN(new_n1100));
  XOR2_X1   g675(.A(new_n1100), .B(KEYINPUT115), .Z(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1074), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1097), .A2(new_n1076), .B1(new_n1066), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1086), .A2(new_n1096), .A3(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1051), .A2(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT118), .B(G1956), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1080), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1109), .A2(KEYINPUT120), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n567), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n567), .A2(new_n573), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1109), .B2(KEYINPUT120), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1106), .A2(new_n1108), .A3(new_n1114), .ZN(new_n1116));
  AOI21_X1  g691(.A(G1348), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n988), .A2(new_n1002), .A3(G2067), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n619), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1110), .A2(new_n1115), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1106), .A2(new_n1108), .A3(new_n1114), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1114), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1116), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n618), .A2(KEYINPUT121), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1047), .A2(G1996), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1065), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n619), .B1(new_n1119), .B2(KEYINPUT60), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  NOR4_X1   g713(.A1(new_n1117), .A2(new_n1118), .A3(new_n1138), .A4(new_n608), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1137), .A2(new_n1139), .B1(KEYINPUT60), .B2(new_n1119), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT59), .B(new_n1130), .C1(new_n1131), .C2(new_n1133), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1136), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1121), .B1(new_n1129), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1033), .A2(new_n1027), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n472), .A2(KEYINPUT126), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n472), .A2(KEYINPUT126), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n444), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n476), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1045), .A2(new_n1145), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1048), .A2(new_n1036), .A3(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(G171), .B(KEYINPUT54), .Z(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1040), .A2(new_n1151), .A3(new_n1048), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1144), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1029), .A2(new_n1034), .A3(new_n1157), .A4(new_n1049), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1085), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1000), .B1(new_n1104), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n989), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(G1996), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT46), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n992), .B2(new_n721), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT47), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n994), .A2(new_n995), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n732), .A2(G2067), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1161), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n989), .A2(new_n810), .A3(new_n595), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT48), .Z(new_n1171));
  NOR2_X1   g746(.A1(new_n998), .A2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1166), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1160), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g749(.A1(new_n671), .A2(G319), .ZN(new_n1176));
  NOR3_X1   g750(.A1(G229), .A2(G401), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n977), .A2(new_n978), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n1177), .A2(new_n879), .A3(new_n1178), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


