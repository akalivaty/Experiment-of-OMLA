//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n460), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n482));
  OR2_X1    g057(.A1(G102), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n485), .A3(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n461), .B2(new_n462), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n462), .C2(new_n461), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(new_n500), .B1(new_n497), .B2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G62), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n495), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n498), .A2(new_n500), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n497), .A2(G543), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n505), .A2(G88), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n504), .A2(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(new_n501), .A2(G89), .A3(new_n508), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n505), .A2(G63), .A3(G651), .A4(new_n509), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n499), .B1(new_n506), .B2(new_n507), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n517), .A2(new_n518), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G168));
  NAND2_X1  g099(.A1(new_n521), .A2(G52), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n501), .A2(new_n508), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n499), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT68), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n509), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n529), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n495), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n521), .A2(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(KEYINPUT69), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n521), .B2(G53), .ZN(new_n553));
  OAI211_X1 g128(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n551), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT70), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n521), .A2(G53), .A3(new_n552), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n551), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n505), .A2(G65), .A3(new_n509), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n495), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n501), .A2(G91), .A3(new_n508), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n561), .A2(new_n567), .ZN(G299));
  AND3_X1   g143(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(new_n570), .A3(new_n517), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  OAI21_X1  g150(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n505), .A2(G87), .A3(new_n508), .A4(new_n509), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n521), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n505), .A2(G61), .A3(new_n509), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n495), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n505), .A2(G86), .A3(new_n508), .A4(new_n509), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n521), .A2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n521), .A2(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n526), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n501), .A2(G60), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n588), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n495), .B1(new_n593), .B2(new_n594), .ZN(new_n598));
  NOR3_X1   g173(.A1(new_n591), .A2(new_n598), .A3(KEYINPUT72), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n521), .A2(KEYINPUT73), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n514), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n605), .A3(G54), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT74), .B(G66), .Z(new_n607));
  AOI22_X1  g182(.A1(new_n501), .A2(new_n607), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n606), .B1(new_n608), .B2(new_n495), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n526), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n501), .A2(KEYINPUT10), .A3(G92), .A4(new_n508), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n602), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n602), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(G286), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n565), .B1(new_n619), .B2(new_n495), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n556), .B2(new_n560), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT75), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n618), .B1(new_n622), .B2(new_n617), .ZN(G297));
  AOI21_X1  g198(.A(new_n618), .B1(new_n622), .B2(new_n617), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n614), .B1(new_n625), .B2(G860), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT76), .Z(G148));
  OAI221_X1 g202(.A(new_n541), .B1(new_n526), .B2(new_n542), .C1(new_n539), .C2(new_n495), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n617), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n612), .A2(new_n613), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(new_n606), .C1(new_n495), .C2(new_n608), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n629), .B1(new_n632), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g209(.A(KEYINPUT3), .B(G2104), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(new_n468), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n474), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n476), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n460), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT77), .B(G2438), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n654), .A3(new_n652), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(KEYINPUT14), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n665), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT78), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(KEYINPUT78), .A3(new_n665), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n669), .B2(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT79), .Z(new_n674));
  XNOR2_X1  g249(.A(G2072), .B(G2078), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n672), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n675), .B(KEYINPUT17), .Z(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n678), .A3(new_n672), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(new_n639), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT80), .B(G2096), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n689), .A2(new_n690), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  MUX2_X1   g271(.A(new_n696), .B(new_n695), .S(new_n688), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT81), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n701), .A2(new_n703), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n701), .A2(new_n703), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n708), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(G229));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G20), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT23), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n621), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT102), .ZN(new_n716));
  INV_X1    g291(.A(G1956), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G35), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT101), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT29), .Z(new_n723));
  INV_X1    g298(.A(G2090), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n716), .A2(new_n717), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n718), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT103), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n712), .A2(G19), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n544), .B2(new_n712), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT89), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1341), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n733));
  NOR2_X1   g308(.A1(G4), .A2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT88), .Z(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n631), .B2(new_n712), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1348), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n719), .A2(G26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  AOI22_X1  g315(.A1(G128), .A2(new_n476), .B1(new_n474), .B2(G140), .ZN(new_n741));
  INV_X1    g316(.A(G104), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n742), .A2(new_n460), .A3(KEYINPUT90), .ZN(new_n743));
  AOI21_X1  g318(.A(KEYINPUT90), .B1(new_n742), .B2(new_n460), .ZN(new_n744));
  OAI221_X1 g319(.A(G2104), .B1(G116), .B2(new_n460), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(new_n719), .ZN(new_n748));
  INV_X1    g323(.A(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n737), .A2(new_n750), .ZN(new_n751));
  OR3_X1    g326(.A1(new_n732), .A2(new_n733), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n733), .B1(new_n732), .B2(new_n751), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n719), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G164), .B2(new_n719), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(G160), .A2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n760), .B2(KEYINPUT24), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(KEYINPUT24), .B2(new_n760), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(G2084), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n758), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n474), .A2(G139), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n635), .A2(G127), .ZN(new_n773));
  INV_X1    g348(.A(G115), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n467), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n772), .B1(G2105), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G29), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT94), .ZN(new_n778));
  OR2_X1    g353(.A1(G29), .A2(G33), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n782));
  OAI21_X1  g357(.A(G2072), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(G2072), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n784), .A2(new_n785), .A3(new_n780), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n767), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n712), .A2(G5), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G301), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1961), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT30), .B(G28), .ZN(new_n792));
  OR2_X1    g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  NAND2_X1  g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n792), .A2(new_n719), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n646), .B2(new_n719), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT98), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n719), .A2(G32), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT26), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G129), .B2(new_n476), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(new_n719), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT27), .B(G1996), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n791), .A2(new_n797), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(G2084), .B1(new_n759), .B2(new_n762), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n805), .B2(new_n807), .ZN(new_n811));
  INV_X1    g386(.A(new_n789), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G1961), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT99), .ZN(new_n814));
  NAND2_X1  g389(.A1(G168), .A2(G16), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(KEYINPUT96), .C1(G16), .C2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(KEYINPUT96), .B2(new_n815), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT97), .B(G1966), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n787), .A2(new_n809), .A3(new_n814), .A4(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT100), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n820), .A2(KEYINPUT100), .B1(new_n724), .B2(new_n723), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n728), .A2(new_n754), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT85), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n577), .A2(new_n578), .ZN(new_n826));
  INV_X1    g401(.A(G74), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n495), .B1(new_n533), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n825), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n576), .A2(KEYINPUT85), .A3(new_n577), .A4(new_n578), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  MUX2_X1   g406(.A(G23), .B(new_n831), .S(G16), .Z(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT33), .B(G1976), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT86), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(KEYINPUT86), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n712), .A2(G22), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n712), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1971), .ZN(new_n843));
  NOR2_X1   g418(.A1(G6), .A2(G16), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n586), .B2(G16), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT32), .B(G1981), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n839), .A2(new_n840), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT34), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(G25), .A2(G29), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n474), .A2(G131), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n476), .A2(G119), .ZN(new_n854));
  OR2_X1    g429(.A1(G95), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n852), .B1(new_n858), .B2(G29), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G1991), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT82), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(KEYINPUT87), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n712), .A2(G24), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT83), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT84), .ZN(new_n866));
  OAI21_X1  g441(.A(G16), .B1(G290), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n600), .A2(KEYINPUT84), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n863), .B1(new_n869), .B2(G1986), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(G1986), .B2(new_n869), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n824), .B1(new_n851), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n851), .A2(new_n824), .A3(new_n871), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n823), .B1(new_n873), .B2(new_n874), .ZN(G311));
  AND3_X1   g450(.A1(new_n754), .A2(new_n821), .A3(new_n822), .ZN(new_n876));
  INV_X1    g451(.A(new_n874), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n728), .B(new_n876), .C1(new_n877), .C2(new_n872), .ZN(G150));
  NAND3_X1  g453(.A1(new_n501), .A2(G93), .A3(new_n508), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT104), .B(G55), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n521), .A2(new_n880), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n879), .B(new_n881), .C1(new_n882), .C2(new_n495), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(G80), .A2(G543), .ZN(new_n886));
  INV_X1    g461(.A(G67), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n533), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(G651), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n889), .A2(KEYINPUT105), .A3(new_n879), .A4(new_n881), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G860), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT37), .Z(new_n893));
  NOR2_X1   g468(.A1(new_n628), .A2(new_n883), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n891), .B2(new_n628), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n614), .A2(G559), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(KEYINPUT39), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT106), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n898), .A2(KEYINPUT39), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(G860), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n893), .B1(new_n900), .B2(new_n902), .ZN(G145));
  XOR2_X1   g478(.A(new_n646), .B(G160), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n480), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n746), .B(G164), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(new_n803), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n803), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n776), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n776), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n637), .B(new_n857), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n460), .A2(KEYINPUT107), .A3(G118), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT107), .B1(new_n460), .B2(G118), .ZN(new_n918));
  OR2_X1    g493(.A1(G106), .A2(G2105), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n917), .A2(G2104), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n476), .A2(G130), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n474), .A2(G142), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n916), .A2(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT108), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n925), .B2(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n907), .B1(new_n915), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n915), .A2(new_n931), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n915), .A2(new_n931), .A3(new_n907), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n906), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n913), .A2(new_n914), .A3(new_n927), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT110), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n933), .A3(new_n906), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n938), .A2(KEYINPUT110), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT40), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(G395));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n504), .B2(new_n515), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n504), .A2(new_n515), .A3(new_n947), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n829), .B(new_n830), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n831), .A3(new_n948), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n586), .B1(new_n597), .B2(new_n599), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n592), .A2(new_n596), .A3(new_n588), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT72), .B1(new_n591), .B2(new_n598), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(G305), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n951), .A2(new_n955), .A3(new_n953), .A4(new_n958), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n960), .A2(new_n963), .A3(KEYINPUT42), .A4(new_n961), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n891), .A2(new_n628), .ZN(new_n969));
  INV_X1    g544(.A(new_n894), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n632), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n895), .B1(G559), .B2(new_n631), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n631), .A2(G299), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n621), .A2(new_n614), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT41), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT41), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n976), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n968), .B(new_n979), .C1(new_n981), .C2(new_n974), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(new_n981), .B2(new_n974), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n967), .A3(new_n966), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G868), .ZN(new_n986));
  INV_X1    g561(.A(new_n891), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(G868), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n946), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  AOI211_X1 g565(.A(KEYINPUT113), .B(new_n988), .C1(new_n985), .C2(G868), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(G295));
  NAND2_X1  g567(.A1(new_n986), .A2(new_n989), .ZN(G331));
  AOI22_X1  g568(.A1(new_n529), .A2(new_n536), .B1(new_n569), .B2(new_n517), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(G171), .B2(new_n573), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n895), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n994), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(G286), .B2(G301), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n980), .B1(new_n971), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n895), .A2(KEYINPUT114), .A3(new_n995), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n978), .A2(new_n977), .ZN(new_n1004));
  AOI21_X1  g579(.A(G301), .B1(new_n571), .B2(new_n572), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n544), .B1(new_n885), .B2(new_n890), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n1005), .A2(new_n994), .B1(new_n1006), .B2(new_n894), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n996), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1003), .A2(new_n1009), .A3(new_n962), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n895), .A2(KEYINPUT114), .A3(new_n995), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT114), .B1(new_n895), .B2(new_n995), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1013), .A2(new_n1001), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  INV_X1    g590(.A(new_n961), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n951), .A2(new_n953), .B1(new_n955), .B2(new_n958), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n960), .A2(KEYINPUT115), .A3(new_n961), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n937), .B(new_n1010), .C1(new_n1014), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n998), .A2(new_n1007), .A3(new_n1002), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1004), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1001), .A2(new_n996), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1020), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1010), .A2(new_n937), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1022), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT44), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1021), .A2(new_n1031), .A3(KEYINPUT43), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1021), .B2(KEYINPUT43), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1027), .A2(new_n1028), .A3(KEYINPUT43), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1030), .B1(new_n1035), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(G164), .B2(G1384), .ZN(new_n1038));
  INV_X1    g613(.A(G125), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n472), .B2(new_n473), .ZN(new_n1040));
  INV_X1    g615(.A(new_n464), .ZN(new_n1041));
  OAI21_X1  g616(.A(G2105), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1042), .A2(G40), .A3(new_n469), .A4(new_n466), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n746), .B(new_n749), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(new_n803), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1044), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1048), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n1050));
  INV_X1    g625(.A(G1996), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1047), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT47), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT48), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G290), .A2(G1986), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1055), .B1(new_n1057), .B2(new_n1048), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n803), .B(new_n1051), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n857), .A2(new_n861), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n857), .A2(new_n861), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1059), .A2(new_n1045), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1044), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1056), .A2(KEYINPUT48), .A3(new_n1044), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1058), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1059), .A2(new_n1045), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(new_n1044), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n746), .A2(G2067), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n1068), .A2(KEYINPUT127), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT127), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1044), .A3(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1054), .A2(new_n1066), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n580), .A2(new_n581), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G651), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n583), .A2(new_n584), .ZN(new_n1076));
  INV_X1    g651(.A(G1981), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(G1981), .B1(new_n582), .B2(new_n585), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(KEYINPUT49), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1078), .A2(new_n1079), .A3(KEYINPUT118), .A4(KEYINPUT49), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT49), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1085));
  INV_X1    g660(.A(G8), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n491), .A2(new_n493), .ZN(new_n1087));
  INV_X1    g662(.A(new_n487), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1384), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G40), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n465), .A2(new_n470), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1084), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G288), .A2(G1976), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1078), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1092), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n829), .A2(G1976), .A3(new_n830), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1092), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT52), .ZN(new_n1102));
  INV_X1    g677(.A(G1976), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(G288), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(new_n1104), .A3(new_n1092), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1084), .B2(new_n1094), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n504), .B2(new_n515), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT55), .B(G8), .C1(new_n504), .C2(new_n515), .ZN(new_n1111));
  INV_X1    g686(.A(G1971), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1037), .A2(G1384), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1091), .B1(G164), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n493), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n492), .B1(new_n635), .B2(new_n489), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n482), .B(new_n486), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1384), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT45), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1112), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT50), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1118), .A2(new_n1123), .A3(new_n1119), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1122), .A2(new_n1124), .A3(new_n724), .A4(new_n1091), .ZN(new_n1125));
  AOI221_X4 g700(.A(new_n1086), .B1(new_n1110), .B2(new_n1111), .C1(new_n1121), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1107), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1099), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(G8), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1043), .B1(new_n1118), .B2(new_n1113), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(KEYINPUT53), .A3(new_n1038), .A4(new_n757), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1123), .A2(new_n1119), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1091), .B1(G164), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1123), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n790), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1133), .A2(new_n757), .A3(new_n1038), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT53), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(G301), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1132), .A2(new_n1107), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G1966), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1146));
  INV_X1    g721(.A(G2084), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1122), .A2(new_n1124), .A3(new_n1147), .A4(new_n1091), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G8), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n523), .A2(KEYINPUT122), .A3(G8), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n523), .B2(G8), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1151), .B1(new_n1155), .B2(KEYINPUT124), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1150), .A2(new_n1156), .A3(new_n1155), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1154), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1152), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT51), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1086), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(new_n1159), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT123), .B1(new_n1149), .B2(new_n1159), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1149), .A2(KEYINPUT123), .A3(new_n1159), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1157), .B(new_n1163), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1144), .B1(KEYINPUT62), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1149), .A2(new_n1159), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1149), .A2(KEYINPUT123), .A3(new_n1159), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1157), .A4(new_n1163), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1128), .B1(new_n1167), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1139), .A2(KEYINPUT125), .A3(G301), .A4(new_n1142), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1142), .A2(G301), .A3(new_n1138), .A4(new_n1134), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1176), .B(new_n1177), .C1(new_n1180), .C2(new_n1143), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1136), .A2(new_n1137), .A3(G2090), .ZN(new_n1182));
  AOI21_X1  g757(.A(G1971), .B1(new_n1133), .B2(new_n1038), .ZN(new_n1183));
  OAI21_X1  g758(.A(G8), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1129), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1130), .A2(G8), .A3(new_n1129), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1186), .A2(new_n1187), .A3(new_n1095), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(G171), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1192), .A2(KEYINPUT54), .A3(new_n1178), .ZN(new_n1193));
  AND4_X1   g768(.A1(new_n1181), .A2(new_n1190), .A3(new_n1166), .A4(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n717), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1195));
  XNOR2_X1  g770(.A(KEYINPUT56), .B(G2072), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1133), .A2(new_n1038), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n561), .A2(new_n567), .A3(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n557), .A2(new_n559), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1199), .B(new_n565), .C1(new_n619), .C2(new_n495), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT57), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1198), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1201), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1195), .B(new_n1197), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(G1348), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1089), .A2(new_n749), .A3(new_n1091), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n631), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1198), .A2(new_n1203), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1205), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1208), .A2(KEYINPUT60), .A3(new_n1209), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n614), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1208), .A2(KEYINPUT60), .A3(new_n631), .A4(new_n1209), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(KEYINPUT60), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1118), .A2(new_n1113), .ZN(new_n1226));
  NAND4_X1  g801(.A1(new_n1038), .A2(new_n1051), .A3(new_n1091), .A4(new_n1226), .ZN(new_n1227));
  XOR2_X1   g802(.A(KEYINPUT58), .B(G1341), .Z(new_n1228));
  NAND2_X1  g803(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1228), .B1(new_n1229), .B2(new_n1043), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1231), .A2(KEYINPUT121), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT121), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1227), .A2(new_n1233), .A3(new_n1230), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1225), .B1(new_n1235), .B2(new_n544), .ZN(new_n1236));
  AND3_X1   g811(.A1(new_n1227), .A2(new_n1233), .A3(new_n1230), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1233), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1238));
  OAI211_X1 g813(.A(new_n1225), .B(new_n544), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1239));
  INV_X1    g814(.A(new_n1239), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1224), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1215), .A2(new_n1206), .ZN(new_n1242));
  INV_X1    g817(.A(KEYINPUT61), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g819(.A1(new_n1215), .A2(KEYINPUT61), .A3(new_n1206), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1217), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1194), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g823(.A(KEYINPUT63), .ZN(new_n1249));
  INV_X1    g824(.A(KEYINPUT119), .ZN(new_n1250));
  NAND3_X1  g825(.A1(new_n1162), .A2(new_n1250), .A3(new_n573), .ZN(new_n1251));
  INV_X1    g826(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1250), .B1(new_n1162), .B2(new_n573), .ZN(new_n1253));
  NOR2_X1   g828(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g829(.A(new_n1249), .B1(new_n1254), .B2(new_n1189), .ZN(new_n1255));
  NAND3_X1  g830(.A1(new_n1149), .A2(G8), .A3(new_n573), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1256), .A2(KEYINPUT119), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1257), .A2(new_n1251), .ZN(new_n1258));
  NAND4_X1  g833(.A1(new_n1258), .A2(new_n1132), .A3(KEYINPUT63), .A4(new_n1107), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g835(.A1(new_n1175), .A2(new_n1248), .A3(new_n1260), .ZN(new_n1261));
  XOR2_X1   g836(.A(new_n600), .B(G1986), .Z(new_n1262));
  OAI21_X1  g837(.A(new_n1044), .B1(new_n1262), .B2(new_n1063), .ZN(new_n1263));
  XNOR2_X1  g838(.A(new_n1263), .B(KEYINPUT117), .ZN(new_n1264));
  AOI21_X1  g839(.A(KEYINPUT126), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g840(.A1(new_n1157), .A2(new_n1163), .ZN(new_n1266));
  NOR2_X1   g841(.A1(new_n1165), .A2(new_n1164), .ZN(new_n1267));
  OAI21_X1  g842(.A(KEYINPUT62), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g843(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1269));
  NAND3_X1  g844(.A1(new_n1268), .A2(new_n1174), .A3(new_n1269), .ZN(new_n1270));
  AOI22_X1  g845(.A1(new_n1098), .A2(new_n1092), .B1(new_n1107), .B2(new_n1126), .ZN(new_n1271));
  NAND3_X1  g846(.A1(new_n1260), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g847(.A(new_n1222), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1273));
  OAI21_X1  g848(.A(new_n544), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1274));
  NAND2_X1  g849(.A1(new_n1274), .A2(KEYINPUT59), .ZN(new_n1275));
  AOI21_X1  g850(.A(new_n1273), .B1(new_n1275), .B2(new_n1239), .ZN(new_n1276));
  AND3_X1   g851(.A1(new_n1215), .A2(KEYINPUT61), .A3(new_n1206), .ZN(new_n1277));
  AOI21_X1  g852(.A(KEYINPUT61), .B1(new_n1215), .B2(new_n1206), .ZN(new_n1278));
  NOR2_X1   g853(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g854(.A(new_n1216), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g855(.A1(new_n1181), .A2(new_n1190), .A3(new_n1193), .A4(new_n1166), .ZN(new_n1281));
  NOR2_X1   g856(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g857(.A(KEYINPUT126), .B(new_n1264), .C1(new_n1272), .C2(new_n1282), .ZN(new_n1283));
  INV_X1    g858(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g859(.A(new_n1073), .B1(new_n1265), .B2(new_n1284), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g860(.A1(G227), .A2(new_n458), .ZN(new_n1287));
  AND3_X1   g861(.A1(new_n707), .A2(new_n710), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g862(.A(G401), .ZN(new_n1289));
  OAI211_X1 g863(.A(new_n1288), .B(new_n1289), .C1(new_n936), .C2(new_n942), .ZN(new_n1290));
  NOR2_X1   g864(.A1(new_n1035), .A2(new_n1290), .ZN(G308));
  OR3_X1    g865(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1292));
  INV_X1    g866(.A(new_n1290), .ZN(new_n1293));
  NAND2_X1  g867(.A1(new_n1292), .A2(new_n1293), .ZN(G225));
endmodule


