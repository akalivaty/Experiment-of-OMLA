//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n208), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n206), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n211), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n230), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  AND2_X1   g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n244), .A2(new_n222), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n232), .A2(G1698), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n251), .B(new_n252), .C1(G226), .C2(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G97), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n246), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT67), .B1(new_n244), .B2(new_n222), .ZN(new_n256));
  AND2_X1   g0056(.A1(G1), .A2(G13), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n256), .A2(new_n260), .A3(G238), .A4(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n256), .A2(G274), .A3(new_n260), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT66), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G41), .A2(G45), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G1), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n205), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n262), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT71), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n262), .B(new_n271), .C1(new_n263), .C2(new_n268), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n255), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT13), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT72), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n255), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n244), .A2(KEYINPUT67), .A3(new_n222), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n266), .A2(new_n267), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(G274), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n271), .B1(new_n281), .B2(new_n262), .ZN(new_n282));
  INV_X1    g0082(.A(new_n272), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT13), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n275), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G169), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT14), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT14), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n286), .A2(new_n290), .A3(G169), .A4(new_n287), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n273), .A2(new_n274), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n285), .A2(G179), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n289), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n222), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G68), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n206), .A2(G1), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n298), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(KEYINPUT73), .A3(new_n300), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT73), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n298), .B2(G68), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n304), .A2(KEYINPUT12), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(KEYINPUT12), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n302), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G20), .A2(G33), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G50), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n313), .A2(new_n314), .B1(new_n206), .B2(G68), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n206), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n202), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n296), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT11), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n310), .A2(new_n311), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n294), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(new_n284), .B2(KEYINPUT13), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n323), .B2(new_n292), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n286), .A2(G200), .A3(new_n287), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  INV_X1    g0128(.A(G150), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n316), .B1(new_n329), .B2(new_n313), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT70), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n330), .A2(new_n331), .B1(new_n206), .B2(new_n201), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n330), .A2(new_n331), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n296), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n299), .A2(new_n314), .A3(new_n301), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n314), .B2(new_n303), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT68), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n251), .B2(new_n202), .ZN(new_n339));
  AOI21_X1  g0139(.A(G1698), .B1(new_n249), .B2(new_n250), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G222), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(KEYINPUT68), .B2(new_n341), .ZN(new_n343));
  INV_X1    g0143(.A(G223), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G1698), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n251), .A2(KEYINPUT69), .A3(G1698), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n245), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n279), .A2(G226), .A3(new_n261), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n281), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n337), .B1(new_n358), .B2(G169), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n357), .A2(G179), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT9), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n357), .A2(G200), .B1(new_n337), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n357), .A2(new_n322), .B1(new_n362), .B2(new_n337), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT10), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n365), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT10), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(new_n363), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n361), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT17), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n328), .A2(new_n301), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n299), .B1(KEYINPUT77), .B2(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n372), .A2(KEYINPUT77), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(new_n303), .B2(new_n328), .ZN(new_n375));
  AND2_X1   g0175(.A1(G58), .A2(G68), .ZN(new_n376));
  NOR2_X1   g0176(.A1(G58), .A2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n312), .A2(G159), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(G20), .C1(new_n376), .C2(new_n377), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n348), .B2(new_n206), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n250), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT76), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n249), .A2(new_n206), .A3(new_n250), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n300), .B1(new_n392), .B2(new_n385), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT76), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT16), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n382), .A2(new_n380), .ZN(new_n396));
  XNOR2_X1  g0196(.A(G58), .B(G68), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n381), .B1(new_n397), .B2(G20), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n387), .A2(new_n399), .A3(KEYINPUT16), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n296), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n375), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n256), .A2(new_n260), .A3(G232), .A4(new_n261), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n263), .B2(new_n268), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n344), .A2(new_n349), .ZN(new_n405));
  INV_X1    g0205(.A(G226), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n407), .C1(new_n346), .C2(new_n347), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(KEYINPUT78), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n409), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n246), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n404), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G190), .ZN(new_n415));
  INV_X1    g0215(.A(G200), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n371), .B1(new_n402), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n375), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n399), .B1(new_n393), .B2(KEYINPUT76), .ZN(new_n421));
  AOI211_X1 g0221(.A(new_n388), .B(new_n300), .C1(new_n392), .C2(new_n385), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n393), .A2(new_n383), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n297), .B1(new_n424), .B2(KEYINPUT16), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n419), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n411), .A2(new_n412), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n245), .A3(new_n410), .ZN(new_n428));
  INV_X1    g0228(.A(new_n404), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n428), .A2(new_n429), .A3(G179), .ZN(new_n430));
  INV_X1    g0230(.A(G169), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT18), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n414), .A2(G179), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n431), .B2(new_n414), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n402), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n428), .A2(new_n429), .A3(G190), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n416), .B1(new_n428), .B2(new_n429), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n418), .A2(new_n434), .A3(new_n438), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n279), .A2(G244), .A3(new_n261), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n281), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n340), .A2(G232), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(new_n251), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n350), .A2(new_n351), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G238), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n447), .B1(new_n452), .B2(new_n246), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G200), .ZN(new_n454));
  INV_X1    g0254(.A(new_n328), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(new_n312), .B1(G20), .B2(G77), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT15), .B(G87), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n457), .A2(new_n316), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n297), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(G77), .B1(new_n206), .B2(G1), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n299), .A2(new_n460), .B1(G77), .B2(new_n298), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n454), .B(new_n462), .C1(new_n322), .C2(new_n453), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n453), .A2(G179), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n453), .B2(new_n431), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n370), .A2(new_n444), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n327), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n205), .B(G45), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n279), .A2(KEYINPUT80), .A3(G274), .A4(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n263), .B2(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n471), .A2(new_n256), .A3(new_n260), .ZN(new_n477));
  OAI211_X1 g0277(.A(G264), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n478));
  OAI211_X1 g0278(.A(G257), .B(new_n349), .C1(new_n346), .C2(new_n347), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n249), .A2(G303), .A3(new_n250), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n477), .A2(G270), .B1(new_n481), .B2(new_n245), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n205), .A2(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n298), .A2(new_n484), .A3(new_n222), .A4(new_n295), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G116), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G116), .B2(new_n303), .ZN(new_n487));
  AOI21_X1  g0287(.A(G20), .B1(G33), .B2(G283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n248), .A2(G97), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G116), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n295), .A2(new_n222), .B1(G20), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT20), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n492), .B1(new_n488), .B2(new_n489), .ZN(new_n499));
  OAI211_X1 g0299(.A(KEYINPUT20), .B(new_n496), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n487), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n483), .A2(new_n502), .A3(KEYINPUT21), .A4(G169), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT84), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n431), .B1(new_n476), .B2(new_n482), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT84), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT21), .A4(new_n502), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT21), .B1(new_n505), .B2(new_n502), .ZN(new_n509));
  INV_X1    g0309(.A(new_n502), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n476), .A2(new_n482), .A3(G179), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G257), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n514));
  OAI211_X1 g0314(.A(G250), .B(new_n349), .C1(new_n346), .C2(new_n347), .ZN(new_n515));
  INV_X1    g0315(.A(G294), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n248), .C2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(G264), .A2(new_n477), .B1(new_n517), .B2(new_n245), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n476), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n431), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n206), .B(G87), .C1(new_n346), .C2(new_n347), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT22), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n251), .A2(new_n523), .A3(new_n206), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  OR3_X1    g0326(.A1(new_n526), .A2(KEYINPUT85), .A3(G20), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n206), .B2(G107), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n449), .A2(KEYINPUT23), .A3(G20), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT85), .B1(new_n526), .B2(G20), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n527), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT24), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT24), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n525), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n297), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT79), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n297), .A2(new_n539), .A3(new_n298), .A4(new_n484), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n485), .A2(KEYINPUT79), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(G107), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n298), .A2(G107), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n543), .B(KEYINPUT25), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI221_X1 g0345(.A(new_n520), .B1(G179), .B2(new_n519), .C1(new_n538), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n508), .A2(new_n513), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  OAI211_X1 g0348(.A(G250), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n549));
  OAI211_X1 g0349(.A(G244), .B(new_n349), .C1(new_n346), .C2(new_n347), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT4), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT4), .B1(new_n340), .B2(G244), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n245), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n477), .A2(G257), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n476), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G200), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n540), .A2(new_n541), .A3(G97), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n298), .A2(G97), .ZN(new_n559));
  OAI21_X1  g0359(.A(G107), .B1(new_n384), .B2(new_n386), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  AND2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n449), .A2(KEYINPUT6), .A3(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(G20), .B1(G77), .B2(new_n312), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n559), .B1(new_n568), .B2(new_n296), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n476), .A2(G190), .A3(new_n554), .A4(new_n555), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n557), .A2(new_n558), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n537), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n536), .B1(new_n525), .B2(new_n533), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n296), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n545), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n518), .A2(new_n476), .A3(new_n322), .ZN(new_n576));
  AOI21_X1  g0376(.A(G200), .B1(new_n518), .B2(new_n476), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT19), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n206), .B1(new_n254), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n563), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n206), .B(G68), .C1(new_n346), .C2(new_n347), .ZN(new_n584));
  INV_X1    g0384(.A(G97), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n579), .B1(new_n316), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n296), .ZN(new_n588));
  INV_X1    g0388(.A(new_n457), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n298), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n540), .A2(new_n541), .A3(G87), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT82), .A4(G87), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(G244), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n596));
  OAI211_X1 g0396(.A(G238), .B(new_n349), .C1(new_n346), .C2(new_n347), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n597), .A3(new_n526), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n245), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n205), .A2(G45), .ZN(new_n600));
  INV_X1    g0400(.A(G250), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n600), .A2(G274), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n279), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n599), .A2(new_n604), .A3(new_n322), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n603), .A2(new_n602), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n279), .A2(new_n606), .B1(new_n598), .B2(new_n245), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n607), .B2(G200), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n599), .A2(new_n604), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n587), .A2(new_n296), .B1(new_n303), .B2(new_n457), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n457), .A2(KEYINPUT81), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n457), .A2(KEYINPUT81), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n540), .A2(new_n611), .A3(new_n541), .A4(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n609), .A2(new_n431), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(G179), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n595), .A2(new_n608), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n556), .A2(new_n431), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n568), .A2(new_n296), .ZN(new_n619));
  INV_X1    g0419(.A(new_n559), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n558), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n476), .A2(new_n615), .A3(new_n554), .A4(new_n555), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n571), .A2(new_n578), .A3(new_n617), .A4(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n502), .B1(new_n483), .B2(G200), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n476), .A2(new_n482), .A3(G190), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n547), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n468), .A2(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n366), .A2(new_n369), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT17), .B1(new_n426), .B2(new_n441), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n441), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n326), .A2(new_n464), .A3(new_n465), .ZN(new_n633));
  AOI211_X1 g0433(.A(new_n631), .B(new_n632), .C1(new_n321), .C2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n434), .A2(new_n438), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n630), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n361), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n614), .A2(new_n616), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n624), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n547), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(KEYINPUT26), .A3(new_n617), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT86), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT86), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n643), .A2(new_n646), .A3(KEYINPUT26), .A4(new_n617), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n595), .A2(new_n608), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n639), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n650), .B2(new_n623), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n645), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n468), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n637), .A2(new_n638), .A3(new_n654), .ZN(G369));
  INV_X1    g0455(.A(new_n627), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n508), .A2(new_n513), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(G213), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n510), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n665), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n508), .B2(new_n513), .ZN(new_n668));
  OAI211_X1 g0468(.A(G330), .B(new_n656), .C1(new_n666), .C2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n546), .A2(new_n663), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n663), .B1(new_n538), .B2(new_n545), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n578), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n546), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT87), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n673), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n657), .A2(new_n679), .A3(new_n546), .A4(new_n664), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT88), .B1(new_n680), .B2(new_n671), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT88), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n663), .B1(new_n508), .B2(new_n513), .ZN(new_n683));
  AOI211_X1 g0483(.A(new_n682), .B(new_n670), .C1(new_n683), .C2(new_n674), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n678), .B1(new_n681), .B2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n209), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n686), .A2(KEYINPUT89), .A3(G41), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT89), .B1(new_n686), .B2(G41), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n582), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n221), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n689), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n651), .A2(new_n644), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n508), .A2(new_n513), .A3(new_n546), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n695), .B(new_n639), .C1(new_n696), .C2(new_n624), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .A3(new_n664), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n663), .B1(new_n642), .B2(new_n652), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(KEYINPUT29), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n696), .A2(new_n641), .A3(new_n656), .A4(new_n664), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n518), .A2(new_n607), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n511), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n556), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n511), .A2(new_n556), .A3(new_n702), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT30), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n607), .A2(G179), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n556), .A2(new_n519), .A3(new_n710), .A4(new_n483), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n663), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT90), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT30), .B1(new_n703), .B2(new_n704), .ZN(new_n717));
  INV_X1    g0517(.A(new_n711), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT90), .B(new_n711), .C1(new_n708), .C2(KEYINPUT30), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(new_n709), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n664), .A2(new_n714), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n701), .A2(new_n715), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n700), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n694), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR2_X1   g0528(.A1(new_n666), .A2(new_n668), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n627), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT91), .ZN(new_n732));
  INV_X1    g0532(.A(new_n689), .ZN(new_n733));
  INV_X1    g0533(.A(G13), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n205), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n732), .B(new_n669), .C1(new_n733), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n209), .A2(new_n251), .ZN(new_n739));
  INV_X1    g0539(.A(G355), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n739), .A2(new_n740), .B1(G116), .B2(new_n209), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n686), .A2(new_n251), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G45), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n743), .B1(new_n221), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n239), .A2(new_n744), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n741), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n257), .B1(new_n206), .B2(G169), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT92), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(new_n733), .A3(new_n737), .ZN(new_n759));
  INV_X1    g0559(.A(new_n752), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n206), .B1(new_n761), .B2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n585), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n206), .A2(new_n615), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G58), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n416), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G20), .A3(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n581), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n765), .A2(new_n322), .A3(new_n416), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n348), .B(new_n773), .C1(G77), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n206), .A2(G190), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT94), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(KEYINPUT94), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n778), .A2(new_n771), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G107), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n777), .A2(G179), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT95), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n776), .B(new_n782), .C1(new_n300), .C2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n770), .B(new_n789), .C1(G50), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n778), .A2(new_n761), .A3(new_n779), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  INV_X1    g0596(.A(G326), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n790), .A2(new_n797), .B1(new_n762), .B2(new_n516), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G322), .B2(new_n767), .ZN(new_n799));
  INV_X1    g0599(.A(new_n793), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(G329), .ZN(new_n801));
  INV_X1    g0601(.A(new_n772), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n251), .B1(new_n802), .B2(G303), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n803), .B1(new_n804), .B2(new_n774), .C1(new_n805), .C2(new_n780), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n801), .B(new_n806), .C1(new_n787), .C2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n792), .A2(new_n796), .B1(new_n799), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n755), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n759), .B1(new_n760), .B2(new_n809), .C1(new_n730), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n738), .A2(new_n811), .ZN(G396));
  NOR2_X1   g0612(.A1(new_n733), .A2(new_n737), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n760), .A2(new_n754), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT96), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n788), .A2(KEYINPUT97), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n788), .A2(KEYINPUT97), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G283), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n251), .B1(new_n775), .B2(G116), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n449), .B2(new_n772), .C1(new_n804), .C2(new_n793), .ZN(new_n822));
  INV_X1    g0622(.A(G303), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n764), .B1(new_n823), .B2(new_n790), .C1(new_n768), .C2(new_n516), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n780), .A2(new_n581), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G137), .A2(new_n791), .B1(new_n775), .B2(G159), .ZN(new_n827));
  INV_X1    g0627(.A(G143), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(new_n768), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G150), .B2(new_n787), .ZN(new_n830));
  XOR2_X1   g0630(.A(KEYINPUT98), .B(KEYINPUT34), .Z(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n780), .A2(new_n300), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n251), .B1(new_n772), .B2(new_n314), .ZN(new_n835));
  INV_X1    g0635(.A(new_n762), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(G58), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n834), .B(new_n837), .C1(new_n838), .C2(new_n793), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n830), .B2(new_n831), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n820), .A2(new_n826), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n813), .B1(G77), .B2(new_n815), .C1(new_n841), .C2(new_n760), .ZN(new_n842));
  INV_X1    g0642(.A(new_n754), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n466), .A2(new_n663), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n663), .B1(new_n459), .B2(new_n461), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n463), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n466), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n842), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT99), .Z(new_n851));
  INV_X1    g0651(.A(new_n849), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n699), .B(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n725), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n813), .B1(new_n853), .B2(new_n725), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n735), .A2(new_n205), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n653), .A2(new_n852), .A3(new_n664), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n320), .A2(new_n663), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n321), .A2(new_n326), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n326), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n320), .B(new_n663), .C1(new_n294), .C2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n845), .A2(new_n860), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n420), .B1(new_n393), .B2(new_n383), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT100), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n867), .A3(new_n296), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n400), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n866), .B2(new_n296), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n375), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n661), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n443), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n402), .A2(KEYINPUT101), .A3(new_n437), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n426), .A2(new_n441), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n402), .A2(new_n872), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n426), .A2(new_n433), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(KEYINPUT101), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n871), .A2(new_n437), .B1(new_n426), .B2(new_n441), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n880), .B1(new_n884), .B2(new_n873), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n875), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n875), .B(KEYINPUT38), .C1(new_n883), .C2(new_n885), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n865), .A2(new_n890), .B1(new_n636), .B2(new_n661), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  INV_X1    g0692(.A(new_n889), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n402), .A2(new_n437), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n878), .A3(new_n877), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n882), .B2(new_n879), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n426), .A2(new_n661), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n443), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n892), .B1(new_n893), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n321), .A2(new_n663), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n888), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT102), .B1(new_n891), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n860), .A2(new_n845), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n862), .A2(new_n864), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(new_n890), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n636), .A2(new_n661), .ZN(new_n909));
  AND4_X1   g0709(.A1(KEYINPUT102), .A2(new_n904), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n468), .B(new_n698), .C1(KEYINPUT29), .C2(new_n699), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n637), .A3(new_n638), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n911), .B(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(G330), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT31), .B1(new_n712), .B2(new_n663), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n628), .B2(new_n664), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n712), .A2(new_n722), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n849), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT101), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT37), .B1(new_n894), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n402), .A2(new_n417), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(new_n898), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(new_n923), .A3(new_n876), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(new_n896), .B1(new_n443), .B2(new_n898), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n889), .B1(new_n925), .B2(KEYINPUT38), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n907), .A2(new_n919), .A3(KEYINPUT40), .A4(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(new_n921), .B1(KEYINPUT37), .B2(new_n895), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n632), .A2(new_n631), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n878), .B1(new_n635), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n887), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n930), .B1(new_n935), .B2(new_n889), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n936), .A2(new_n907), .A3(KEYINPUT103), .A4(new_n919), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n907), .A2(new_n890), .A3(new_n919), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n929), .A2(new_n937), .B1(new_n930), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n701), .A2(new_n715), .A3(new_n918), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n468), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n915), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n939), .B2(new_n941), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n859), .B1(new_n914), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n914), .B2(new_n943), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(G116), .A3(new_n223), .A4(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n692), .A2(new_n202), .A3(new_n376), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n300), .A2(G50), .ZN(new_n951));
  OAI211_X1 g0751(.A(G1), .B(new_n734), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n945), .A2(new_n949), .A3(new_n952), .ZN(G367));
  OAI21_X1  g0753(.A(new_n756), .B1(new_n209), .B2(new_n457), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n742), .A2(new_n229), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n813), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n762), .A2(new_n300), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n828), .B2(new_n790), .C1(new_n768), .C2(new_n329), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n348), .B1(new_n775), .B2(G50), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n769), .B2(new_n772), .C1(new_n202), .C2(new_n780), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(G137), .C2(new_n800), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n819), .A2(G159), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n819), .A2(G294), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n781), .A2(G97), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT46), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n772), .B2(new_n495), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT108), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n965), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n251), .B1(new_n775), .B2(G283), .ZN(new_n972));
  INV_X1    g0772(.A(G317), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n972), .B1(new_n804), .B2(new_n790), .C1(new_n973), .C2(new_n793), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n802), .A2(KEYINPUT46), .A3(G116), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n449), .B2(new_n762), .C1(new_n768), .C2(new_n823), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n962), .A2(new_n963), .B1(new_n964), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n760), .B1(new_n978), .B2(KEYINPUT47), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n956), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n595), .A2(new_n664), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT104), .Z(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(new_n650), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n640), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n755), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n643), .A2(new_n663), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n621), .A2(new_n663), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n571), .A2(new_n623), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n680), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n623), .B1(new_n990), .B2(new_n546), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n664), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT105), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n984), .A2(new_n985), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n999), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n678), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n991), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1006), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT107), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n681), .A2(new_n684), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n992), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n681), .A2(new_n684), .A3(KEYINPUT107), .A4(new_n991), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n991), .B1(new_n681), .B2(new_n684), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n680), .A2(new_n671), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n682), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n680), .A2(KEYINPUT88), .A3(new_n671), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n1021), .A3(new_n992), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT107), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1012), .A2(new_n1011), .A3(new_n992), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT44), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1015), .A2(new_n1018), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n1005), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n683), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n675), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n680), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n669), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n700), .A3(new_n725), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1015), .A2(new_n1018), .A3(new_n678), .A4(new_n1025), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1027), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n727), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n689), .B(KEYINPUT41), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n737), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n987), .B1(new_n1009), .B2(new_n1040), .ZN(G387));
  INV_X1    g0841(.A(KEYINPUT111), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1030), .B(new_n669), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n726), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1033), .A2(new_n733), .A3(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n739), .A2(new_n690), .B1(G107), .B2(new_n209), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT109), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n235), .A2(G45), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n690), .ZN(new_n1049));
  AOI211_X1 g0849(.A(G45), .B(new_n1049), .C1(G68), .C2(G77), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n328), .A2(G50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n743), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1047), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n813), .B1(new_n1054), .B2(new_n757), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n611), .A2(new_n612), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n836), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n314), .B2(new_n768), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT110), .Z(new_n1060));
  AOI21_X1  g0860(.A(new_n348), .B1(new_n775), .B2(G68), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n202), .B2(new_n772), .C1(new_n794), .C2(new_n790), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n965), .B1(new_n329), .B2(new_n793), .C1(new_n788), .C2(new_n328), .ZN(new_n1063));
  OR3_X1    g0863(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n251), .B1(new_n800), .B2(G326), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n772), .A2(new_n516), .B1(new_n762), .B2(new_n805), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n767), .A2(G317), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G303), .A2(new_n775), .B1(new_n791), .B2(G322), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n818), .C2(new_n804), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1065), .B1(new_n495), .B2(new_n780), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1064), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1055), .B1(new_n1076), .B2(new_n752), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n675), .A2(new_n755), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1077), .A2(new_n1078), .B1(new_n1032), .B2(new_n737), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1042), .B1(new_n1045), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1045), .A2(new_n1042), .A3(new_n1079), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(G393));
  INV_X1    g0883(.A(KEYINPUT112), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1035), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1027), .A2(new_n1035), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(KEYINPUT112), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n992), .A2(new_n755), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n756), .B1(new_n585), .B2(new_n209), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n743), .A2(new_n242), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n813), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n818), .A2(new_n823), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n768), .A2(new_n804), .B1(new_n790), .B2(new_n973), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n348), .B1(new_n772), .B2(new_n805), .C1(new_n516), .C2(new_n774), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G116), .B2(new_n836), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n800), .A2(G322), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n782), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n818), .A2(new_n314), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n768), .A2(new_n794), .B1(new_n790), .B2(new_n329), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n762), .A2(new_n202), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n251), .B1(new_n774), .B2(new_n328), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G68), .C2(new_n802), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n825), .B1(G143), .B2(new_n800), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1092), .A2(new_n1098), .B1(new_n1099), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1091), .B1(new_n1107), .B2(new_n752), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1087), .A2(new_n737), .B1(new_n1088), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1084), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1033), .B1(new_n1110), .B2(new_n1085), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1036), .A2(new_n733), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1109), .A2(new_n1113), .ZN(G390));
  OAI21_X1  g0914(.A(new_n813), .B1(new_n815), .B2(new_n455), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n251), .B1(new_n774), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n768), .A2(new_n838), .B1(new_n790), .B2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(G159), .C2(new_n836), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n802), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n772), .B2(new_n329), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n800), .A2(G125), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1120), .B(new_n1124), .C1(new_n314), .C2(new_n780), .ZN(new_n1125));
  INV_X1    g0925(.A(G137), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n818), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n818), .A2(new_n449), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n790), .A2(new_n805), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1102), .B(new_n1129), .C1(G116), .C2(new_n767), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n251), .B(new_n773), .C1(G97), .C2(new_n775), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n800), .A2(G294), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n834), .A4(new_n1132), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1125), .A2(new_n1127), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1115), .B1(new_n1134), .B2(new_n752), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n901), .A2(new_n903), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1135), .B1(new_n1137), .B2(new_n754), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n697), .A2(new_n664), .A3(new_n848), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT113), .B1(new_n1139), .B2(new_n845), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1139), .A2(KEYINPUT113), .A3(new_n845), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n907), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n902), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n926), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1136), .B1(new_n902), .B2(new_n865), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n724), .A2(G330), .A3(new_n852), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n907), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n906), .A2(new_n907), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1144), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1153), .A2(new_n1136), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n940), .A2(new_n852), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n915), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n907), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1151), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1138), .B1(new_n1158), .B2(new_n736), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT114), .B1(new_n1149), .B2(new_n907), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n724), .A2(G330), .A3(new_n852), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT114), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1161), .A2(new_n1162), .A3(new_n862), .A4(new_n864), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1160), .A2(new_n1157), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n906), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n862), .B(new_n864), .C1(new_n1155), .C2(new_n915), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1150), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1139), .A2(KEYINPUT113), .A3(new_n845), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n1140), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n468), .A2(G330), .A3(new_n940), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n912), .A2(new_n637), .A3(new_n638), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n689), .B1(new_n1176), .B2(new_n1158), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1145), .B1(new_n1169), .B2(new_n907), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1152), .A2(new_n1144), .B1(new_n901), .B2(new_n903), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n907), .B(new_n1156), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1172), .A2(new_n1180), .A3(new_n1151), .A4(new_n1175), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1159), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(G378));
  AOI22_X1  g0983(.A1(new_n906), .A2(new_n1164), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1175), .B1(new_n1158), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n929), .A2(new_n937), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n915), .B1(new_n938), .B2(new_n930), .ZN(new_n1187));
  XOR2_X1   g0987(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT116), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n337), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n661), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n370), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n370), .A2(new_n1193), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1190), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1196), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1198), .A2(KEYINPUT116), .A3(new_n1194), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1189), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT116), .B1(new_n1198), .B2(new_n1194), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1195), .A2(new_n1190), .A3(new_n1196), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(new_n1188), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1186), .A2(new_n1187), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT102), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n891), .A2(KEYINPUT102), .A3(new_n904), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1204), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1205), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1155), .B1(new_n862), .B2(new_n864), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT103), .B1(new_n1213), .B2(new_n936), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n937), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1187), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1204), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1186), .A2(new_n1187), .A3(new_n1204), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1218), .A2(new_n1219), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1185), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT57), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1210), .B1(new_n1205), .B2(new_n1211), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n911), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(KEYINPUT57), .A3(new_n1185), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n733), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1204), .A2(new_n843), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n813), .B1(G50), .B2(new_n814), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G58), .A2(new_n781), .B1(new_n800), .B2(G283), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n585), .B2(new_n788), .C1(new_n1056), .C2(new_n774), .ZN(new_n1232));
  INV_X1    g1032(.A(G41), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1233), .B(new_n348), .C1(new_n772), .C2(new_n202), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT115), .Z(new_n1235));
  OAI221_X1 g1035(.A(new_n958), .B1(new_n495), .B2(new_n790), .C1(new_n768), .C2(new_n449), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1232), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n774), .A2(new_n1126), .B1(new_n772), .B2(new_n1116), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G150), .B2(new_n836), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G128), .A2(new_n767), .B1(new_n791), .B2(G125), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n788), .C2(new_n838), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n781), .A2(G159), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G33), .B(G41), .C1(new_n800), .C2(G124), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G50), .B1(new_n248), .B2(new_n1233), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n251), .B2(G41), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1238), .A2(new_n1247), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1230), .B1(new_n1251), .B2(new_n752), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1226), .A2(new_n737), .B1(new_n1229), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1228), .A2(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n1184), .A2(new_n1174), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1176), .A2(new_n1255), .A3(new_n1039), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n862), .A2(new_n843), .A3(new_n864), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n813), .B1(new_n815), .B2(G68), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT117), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n790), .A2(new_n838), .B1(new_n762), .B2(new_n314), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n251), .B1(new_n329), .B2(new_n774), .C1(new_n768), .C2(new_n1126), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(G58), .C2(new_n781), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n793), .A2(new_n1118), .B1(new_n772), .B2(new_n794), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT120), .Z(new_n1264));
  OAI211_X1 g1064(.A(new_n1262), .B(new_n1264), .C1(new_n818), .C2(new_n1116), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n790), .A2(new_n516), .B1(new_n774), .B2(new_n449), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n819), .B2(G116), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT118), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n793), .A2(new_n823), .B1(new_n772), .B2(new_n585), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT119), .Z(new_n1270));
  NAND2_X1  g1070(.A1(new_n781), .A2(G77), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n251), .B1(new_n767), .B2(G283), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1058), .A4(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1265), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1259), .B1(new_n1274), .B2(new_n752), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1172), .A2(new_n737), .B1(new_n1257), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1256), .A2(new_n1276), .ZN(G381));
  INV_X1    g1077(.A(G396), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1081), .A2(new_n1278), .A3(new_n1082), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1279), .A2(G384), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1280), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT121), .Z(new_n1282));
  NAND2_X1  g1082(.A1(new_n1226), .A2(new_n737), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1229), .A2(new_n1252), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1224), .A2(new_n1225), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n689), .B1(new_n1286), .B2(KEYINPUT57), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1285), .B1(new_n1287), .B2(new_n1223), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1182), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1282), .A2(new_n1289), .ZN(G407));
  NAND2_X1  g1090(.A1(new_n662), .A2(G213), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT122), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G407), .B(G213), .C1(new_n1289), .C2(new_n1293), .ZN(G409));
  INV_X1    g1094(.A(new_n1082), .ZN(new_n1295));
  OAI21_X1  g1095(.A(G396), .B1(new_n1295), .B2(new_n1080), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1279), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1109), .A2(new_n1113), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1299));
  OAI21_X1  g1099(.A(G387), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1297), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1086), .A2(KEYINPUT112), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1085), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n737), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1088), .A2(new_n1108), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1301), .B1(new_n1302), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n736), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1311));
  AOI22_X1  g1111(.A1(new_n1310), .A2(new_n1311), .B1(new_n986), .B2(new_n981), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1109), .A2(new_n1113), .A3(new_n1297), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1308), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1300), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1300), .A2(new_n1314), .A3(KEYINPUT126), .A4(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1165), .A2(new_n1171), .A3(KEYINPUT60), .A4(new_n1174), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n733), .ZN(new_n1322));
  OAI21_X1  g1122(.A(KEYINPUT60), .B1(new_n1184), .B2(new_n1174), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1255), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1276), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n857), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1323), .A2(new_n1255), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G384), .B(new_n1276), .C1(new_n1327), .C2(new_n1322), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1326), .A2(new_n1328), .A3(KEYINPUT124), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT124), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1330));
  OR2_X1    g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1286), .A2(new_n1039), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1253), .A3(new_n1182), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1334), .B1(G375), .B2(G378), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1331), .A2(new_n1335), .A3(KEYINPUT63), .A4(new_n1293), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1320), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1292), .A2(G2897), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(G2897), .A3(new_n1292), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1339), .A2(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1333), .B1(new_n1288), .B2(new_n1182), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT123), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1292), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  OAI211_X1 g1145(.A(KEYINPUT123), .B(new_n1333), .C1(new_n1288), .C2(new_n1182), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1342), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1337), .A2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1182), .B1(new_n1228), .B2(new_n1253), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1344), .B1(new_n1349), .B2(new_n1334), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1350), .A2(new_n1293), .A3(new_n1331), .A4(new_n1346), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT63), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT125), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1351), .A2(KEYINPUT125), .A3(new_n1352), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1348), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1300), .A2(new_n1314), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1343), .A2(new_n1292), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1361), .A2(new_n1359), .ZN(new_n1362));
  AOI22_X1  g1162(.A1(new_n1351), .A2(new_n1359), .B1(new_n1360), .B2(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1315), .B1(new_n1360), .B2(new_n1342), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1358), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1357), .A2(new_n1365), .ZN(G405));
  INV_X1    g1166(.A(new_n1349), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(new_n1289), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1368), .A2(new_n1361), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1369), .B1(new_n1340), .B2(new_n1368), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1358), .ZN(new_n1371));
  XNOR2_X1  g1171(.A(new_n1371), .B(KEYINPUT127), .ZN(new_n1372));
  XNOR2_X1  g1172(.A(new_n1370), .B(new_n1372), .ZN(G402));
endmodule


