//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946;
  NOR2_X1   g000(.A1(G127gat), .A2(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT69), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n202), .B1(new_n207), .B2(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  NAND2_X1  g011(.A1(G113gat), .A2(G120gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(G113gat), .B2(G120gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n202), .ZN(new_n216));
  NAND2_X1  g015(.A1(G127gat), .A2(G134gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n210), .A2(KEYINPUT70), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n210), .A2(KEYINPUT70), .ZN(new_n220));
  OAI21_X1  g019(.A(G113gat), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n208), .A2(new_n214), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G141gat), .B(G148gat), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G155gat), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n223), .A2(KEYINPUT2), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(G155gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(G162gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT75), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n230), .B2(new_n231), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n233), .A2(new_n234), .A3(new_n223), .ZN(new_n235));
  AND2_X1   g034(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT76), .B(G155gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT2), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n229), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n222), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT75), .B1(new_n225), .B2(new_n227), .ZN(new_n244));
  XOR2_X1   g043(.A(G141gat), .B(G148gat), .Z(new_n245));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT2), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n224), .A2(KEYINPUT76), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G155gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT77), .B(G162gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n228), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT78), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n243), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(new_n241), .B2(new_n222), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n216), .A2(new_n217), .ZN(new_n265));
  INV_X1    g064(.A(new_n215), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT70), .B(G120gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n265), .B(new_n266), .C1(new_n267), .C2(new_n209), .ZN(new_n268));
  INV_X1    g067(.A(G134gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT69), .B(G127gat), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n214), .B(new_n216), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n255), .A2(KEYINPUT79), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n255), .A2(new_n272), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(KEYINPUT4), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT79), .B1(new_n255), .B2(new_n272), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n240), .A2(new_n245), .A3(new_n246), .A4(new_n244), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n222), .A2(new_n282), .A3(new_n263), .A4(new_n228), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT84), .B1(new_n284), .B2(new_n277), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n262), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n255), .A2(new_n272), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n281), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n260), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT81), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n294), .A3(new_n291), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n288), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n241), .B2(new_n242), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n256), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n291), .B1(new_n299), .B2(new_n243), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n276), .A2(new_n280), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT4), .B1(new_n281), .B2(new_n283), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT80), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI211_X1 g104(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n281), .C2(new_n283), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n300), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n296), .A2(KEYINPUT82), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT82), .B1(new_n296), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n287), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G1gat), .B(G29gat), .Z(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G57gat), .B(G85gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n310), .A2(KEYINPUT6), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT85), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n310), .A2(new_n319), .A3(KEYINPUT6), .A4(new_n316), .ZN(new_n320));
  INV_X1    g119(.A(new_n287), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n280), .B1(new_n264), .B2(new_n273), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n301), .B1(new_n323), .B2(KEYINPUT80), .ZN(new_n324));
  INV_X1    g123(.A(new_n306), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n261), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n290), .A2(new_n294), .A3(new_n291), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n294), .B1(new_n290), .B2(new_n291), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT5), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n322), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n296), .A2(new_n307), .A3(KEYINPUT82), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n321), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n315), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT6), .B1(new_n310), .B2(new_n316), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n318), .A2(new_n320), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G226gat), .ZN(new_n336));
  INV_X1    g135(.A(G233gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT67), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT26), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(KEYINPUT68), .A3(new_n342), .ZN(new_n346));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n340), .B2(new_n342), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT28), .B1(new_n352), .B2(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n355));
  INV_X1    g154(.A(G190gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360));
  INV_X1    g159(.A(new_n340), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n340), .A2(KEYINPUT23), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n347), .ZN(new_n365));
  OR3_X1    g164(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n354), .A2(KEYINPUT24), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n366), .A2(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n360), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n341), .A2(KEYINPUT23), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n370), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(G183gat), .B2(G190gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n347), .B(KEYINPUT66), .Z(new_n377));
  NAND4_X1  g176(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n350), .A2(new_n359), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n339), .B1(new_n379), .B2(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n350), .A2(new_n359), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n372), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n338), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G211gat), .B(G218gat), .Z(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT72), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n388));
  OR2_X1    g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(G197gat), .A2(G204gat), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n387), .B(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT73), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n380), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n339), .B1(new_n381), .B2(new_n382), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397));
  INV_X1    g196(.A(new_n382), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n348), .B1(new_n343), .B2(new_n344), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n358), .B1(new_n399), .B2(new_n346), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n397), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n396), .B1(new_n339), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n395), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n393), .B1(new_n403), .B2(new_n392), .ZN(new_n404));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n394), .B1(new_n380), .B2(new_n384), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT73), .B1(new_n401), .B2(new_n339), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n392), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n393), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n407), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT30), .A4(new_n407), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT74), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n410), .B(new_n417), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT86), .B1(new_n335), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n334), .A2(new_n333), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n330), .A2(new_n331), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n315), .B1(new_n425), .B2(new_n287), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n319), .B1(new_n426), .B2(KEYINPUT6), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n428));
  NOR4_X1   g227(.A1(new_n332), .A2(KEYINPUT85), .A3(new_n428), .A4(new_n315), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n424), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431));
  INV_X1    g230(.A(new_n422), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n383), .A2(new_n222), .ZN(new_n434));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT64), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n379), .A2(new_n272), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT32), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT71), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n442));
  XNOR2_X1  g241(.A(G15gat), .B(G43gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G71gat), .B(G99gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n438), .B(KEYINPUT32), .C1(new_n446), .C2(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n437), .ZN(new_n451));
  INV_X1    g250(.A(new_n436), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(KEYINPUT34), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(KEYINPUT34), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n454), .A2(new_n455), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n449), .A3(new_n448), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(KEYINPUT87), .A3(new_n459), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  INV_X1    g263(.A(new_n392), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT3), .B1(new_n465), .B2(new_n397), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT29), .B1(new_n241), .B2(new_n242), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n466), .A2(new_n241), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G78gat), .B(G106gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G228gat), .A2(G233gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G22gat), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT31), .B(G50gat), .Z(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n470), .B(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n423), .A2(new_n433), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n475), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n460), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n430), .A2(new_n432), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n430), .A2(new_n432), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n479), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n460), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n457), .A2(KEYINPUT36), .A3(new_n459), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n416), .B1(new_n415), .B2(KEYINPUT37), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n411), .A2(new_n412), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n392), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT37), .B1(new_n385), .B2(new_n465), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n408), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n407), .B1(new_n404), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n415), .A2(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n500), .B(new_n424), .C1(new_n427), .C2(new_n429), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n286), .A2(new_n259), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT39), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n291), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n504), .A2(new_n315), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n290), .A2(new_n291), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(new_n503), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n279), .A2(new_n285), .B1(new_n299), .B2(new_n243), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n260), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT40), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n504), .A2(new_n509), .A3(KEYINPUT40), .A4(new_n315), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n332), .B2(new_n315), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n479), .B1(new_n513), .B2(new_n422), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n488), .B1(new_n501), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n478), .A2(new_n482), .B1(new_n484), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G29gat), .A2(G36gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT88), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR3_X1   g320(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT15), .A3(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n519), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n522), .A2(new_n529), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n521), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n525), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT90), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n533), .A2(new_n534), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(G1gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(G1gat), .B2(new_n538), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G8gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n536), .A2(new_n543), .B1(new_n542), .B2(new_n533), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT18), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n544), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT12), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT18), .B1(new_n544), .B2(new_n545), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n542), .B(new_n533), .Z(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(new_n545), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n550), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n556), .B1(new_n550), .B2(new_n562), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n516), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT100), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT8), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n571), .B(new_n573), .C1(G85gat), .C2(G92gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n569), .B(new_n574), .Z(new_n575));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n575), .A2(new_n533), .B1(KEYINPUT41), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n537), .A2(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n536), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(KEYINPUT101), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(KEYINPUT101), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G190gat), .B(G218gat), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT99), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n583), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n591), .B(new_n577), .C1(new_n580), .C2(new_n581), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n585), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT104), .ZN(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT9), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT95), .Z(new_n603));
  NOR2_X1   g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(KEYINPUT93), .B2(new_n598), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n597), .B(KEYINPUT94), .ZN(new_n606));
  NOR2_X1   g405(.A1(KEYINPUT93), .A2(KEYINPUT9), .ZN(new_n607));
  OAI221_X1 g406(.A(new_n605), .B1(KEYINPUT93), .B2(new_n598), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(new_n575), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n574), .A2(KEYINPUT102), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n574), .A2(KEYINPUT102), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n569), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT103), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n569), .A2(new_n574), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n611), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n610), .A2(KEYINPUT10), .A3(new_n575), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n618), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n596), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n624), .A2(KEYINPUT104), .A3(new_n625), .A4(new_n629), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n631), .A2(new_n632), .B1(new_n626), .B2(new_n630), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n609), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT98), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n635), .B(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n542), .B1(new_n610), .B2(KEYINPUT21), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT20), .ZN(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G183gat), .B(G211gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n640), .B(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n589), .B1(new_n584), .B2(new_n592), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n595), .A2(new_n633), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n567), .A2(new_n335), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g453(.A1(new_n567), .A2(new_n652), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n432), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT16), .B(G8gat), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(G8gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  MUX2_X1   g459(.A(new_n658), .B(new_n660), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g460(.A(new_n488), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n655), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n462), .A2(new_n463), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n655), .B2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n655), .A2(new_n475), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n594), .A2(new_n649), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n633), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n648), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n567), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(G29gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n675), .A3(new_n335), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT45), .ZN(new_n677));
  NOR2_X1   g476(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n516), .B2(new_n670), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n680));
  AOI21_X1  g479(.A(new_n476), .B1(new_n483), .B2(KEYINPUT86), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n681), .A2(new_n433), .B1(KEYINPUT35), .B2(new_n481), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n515), .A2(new_n484), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n671), .B(new_n680), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n566), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n679), .A2(new_n684), .A3(new_n685), .A4(new_n673), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n686), .B2(new_n430), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n677), .A2(new_n687), .ZN(G1328gat));
  INV_X1    g487(.A(G36gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n689), .A3(new_n422), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT46), .Z(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n686), .B2(new_n432), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  OAI21_X1  g492(.A(G43gat), .B1(new_n686), .B2(new_n662), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT47), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(G43gat), .ZN(new_n697));
  INV_X1    g496(.A(new_n664), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n674), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n696), .B(new_n700), .ZN(G1330gat));
  OAI21_X1  g500(.A(G50gat), .B1(new_n686), .B2(new_n475), .ZN(new_n702));
  INV_X1    g501(.A(G50gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n674), .A2(new_n703), .A3(new_n479), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g506(.A(new_n648), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n594), .A2(new_n708), .A3(new_n649), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n566), .A3(new_n672), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n516), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(KEYINPUT108), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(KEYINPUT108), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n335), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g516(.A1(new_n714), .A2(new_n432), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  AND2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n718), .B2(new_n719), .ZN(G1333gat));
  OAI21_X1  g521(.A(G71gat), .B1(new_n714), .B2(new_n662), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n698), .A2(new_n599), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n714), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g525(.A1(new_n714), .A2(new_n475), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT109), .B(G78gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1335gat));
  AND2_X1   g528(.A1(new_n679), .A2(new_n684), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n685), .A2(new_n648), .A3(new_n633), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G85gat), .B1(new_n732), .B2(new_n430), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n478), .A2(new_n482), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n515), .A2(new_n484), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n685), .A2(new_n648), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n736), .A2(KEYINPUT51), .A3(new_n671), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n670), .B1(new_n734), .B2(new_n735), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT51), .A4(new_n737), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n736), .A2(new_n671), .A3(new_n737), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n739), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n430), .A2(new_n633), .A3(G85gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n733), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n422), .A3(new_n731), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G92gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n633), .A2(new_n432), .A3(G92gat), .ZN(new_n752));
  INV_X1    g551(.A(new_n745), .ZN(new_n753));
  INV_X1    g552(.A(new_n738), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n756), .A2(new_n757), .A3(KEYINPUT52), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n756), .B2(KEYINPUT52), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(new_n750), .B2(G92gat), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n752), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n758), .A2(new_n759), .B1(new_n763), .B2(new_n764), .ZN(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n732), .B2(new_n662), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n664), .A2(new_n633), .A3(G99gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n747), .B2(new_n767), .ZN(G1338gat));
  NOR3_X1   g567(.A1(new_n633), .A2(G106gat), .A3(new_n475), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n753), .B2(new_n754), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n679), .A2(new_n684), .A3(new_n479), .A4(new_n731), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT53), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n746), .A2(new_n775), .A3(new_n769), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n746), .B2(new_n769), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(G106gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n771), .B2(KEYINPUT114), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n730), .A2(new_n781), .A3(new_n479), .A4(new_n731), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT53), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT115), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n746), .A2(new_n769), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT113), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n746), .A2(new_n775), .A3(new_n769), .ZN(new_n787));
  AND4_X1   g586(.A1(KEYINPUT115), .A2(new_n783), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n774), .B1(new_n784), .B2(new_n788), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n651), .B2(new_n685), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n709), .A2(KEYINPUT116), .A3(new_n566), .A4(new_n633), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n558), .A2(new_n560), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n544), .B2(new_n545), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n554), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n563), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n594), .B2(new_n649), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n631), .A2(new_n632), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n620), .A2(new_n621), .B1(G230gat), .B2(G233gat), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n629), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n624), .A2(KEYINPUT54), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n622), .A2(new_n623), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n802), .B(KEYINPUT55), .C1(new_n803), .C2(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n799), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n798), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n563), .A2(new_n796), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n809), .A2(new_n566), .B1(new_n633), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n810), .B1(new_n812), .B2(new_n670), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n793), .B1(new_n813), .B2(new_n648), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n335), .A3(new_n480), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT117), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n814), .A2(new_n817), .A3(new_n335), .A4(new_n480), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n816), .A2(new_n432), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT118), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n209), .A3(new_n685), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n664), .A2(new_n479), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n335), .A2(new_n432), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n814), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n566), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n827), .ZN(G1340gat));
  NAND3_X1  g627(.A1(new_n820), .A2(new_n267), .A3(new_n672), .ZN(new_n829));
  OAI21_X1  g628(.A(G120gat), .B1(new_n826), .B2(new_n633), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1341gat));
  NAND3_X1  g630(.A1(new_n819), .A2(new_n270), .A3(new_n648), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n207), .B1(new_n826), .B2(new_n708), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1342gat));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n670), .A2(G134gat), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n819), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n816), .A2(new_n432), .A3(new_n818), .A4(new_n837), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n269), .B1(new_n825), .B2(new_n671), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(KEYINPUT56), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT119), .B1(new_n839), .B2(KEYINPUT56), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n838), .A2(new_n841), .A3(new_n842), .A4(KEYINPUT120), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1343gat));
  NAND2_X1  g646(.A1(new_n662), .A2(new_n479), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n432), .B1(new_n848), .B2(KEYINPUT123), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n814), .A2(new_n335), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n849), .B(new_n850), .C1(KEYINPUT123), .C2(new_n848), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n566), .A2(G141gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT124), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n824), .A2(new_n662), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT121), .Z(new_n857));
  AND3_X1   g656(.A1(new_n814), .A2(KEYINPUT57), .A3(new_n479), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n814), .B2(new_n479), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n685), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G141gat), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n851), .A2(new_n862), .A3(new_n852), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n854), .A2(new_n855), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n860), .A2(KEYINPUT122), .A3(G141gat), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n866), .A2(new_n867), .A3(new_n853), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n864), .B1(new_n868), .B2(new_n855), .ZN(G1344gat));
  INV_X1    g668(.A(G148gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n870), .A3(new_n672), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n672), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n812), .A2(new_n670), .ZN(new_n874));
  INV_X1    g673(.A(new_n810), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n648), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n651), .A2(new_n685), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT125), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879));
  INV_X1    g678(.A(new_n877), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n879), .B(new_n880), .C1(new_n813), .C2(new_n648), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n479), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n858), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n873), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n870), .B1(new_n886), .B2(KEYINPUT126), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n858), .B1(new_n882), .B2(new_n883), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n873), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n872), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n858), .A2(new_n859), .ZN(new_n892));
  INV_X1    g691(.A(new_n857), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI211_X1 g693(.A(KEYINPUT59), .B(new_n870), .C1(new_n894), .C2(new_n672), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n871), .B1(new_n891), .B2(new_n895), .ZN(G1345gat));
  NAND3_X1  g695(.A1(new_n851), .A2(new_n239), .A3(new_n648), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n648), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(new_n899), .B2(new_n239), .ZN(G1346gat));
  AOI21_X1  g699(.A(new_n253), .B1(new_n851), .B2(new_n671), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n670), .A2(new_n238), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n894), .B2(new_n902), .ZN(G1347gat));
  NAND4_X1  g702(.A1(new_n814), .A2(new_n430), .A3(new_n422), .A4(new_n822), .ZN(new_n904));
  INV_X1    g703(.A(G169gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(new_n566), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n814), .A2(new_n430), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n422), .A3(new_n480), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT127), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n685), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n906), .B1(new_n910), .B2(new_n905), .ZN(G1348gat));
  INV_X1    g710(.A(G176gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(new_n912), .A3(new_n672), .ZN(new_n913));
  OAI21_X1  g712(.A(G176gat), .B1(new_n904), .B2(new_n633), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  OAI21_X1  g714(.A(G183gat), .B1(new_n904), .B2(new_n708), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n648), .A2(new_n351), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n908), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n909), .A2(new_n356), .A3(new_n671), .ZN(new_n920));
  OAI21_X1  g719(.A(G190gat), .B1(new_n904), .B2(new_n670), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1351gat));
  AND4_X1   g722(.A1(new_n422), .A2(new_n907), .A3(new_n479), .A4(new_n662), .ZN(new_n924));
  AOI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n685), .ZN(new_n925));
  INV_X1    g724(.A(new_n889), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n488), .A2(new_n335), .A3(new_n432), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n685), .A2(G197gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  OAI21_X1  g730(.A(G204gat), .B1(new_n928), .B2(new_n633), .ZN(new_n932));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n924), .A2(new_n933), .A3(new_n672), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(G1353gat));
  INV_X1    g736(.A(G211gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n924), .A2(new_n938), .A3(new_n648), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n926), .A2(new_n648), .A3(new_n927), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n928), .B2(new_n670), .ZN(new_n944));
  INV_X1    g743(.A(G218gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n924), .A2(new_n945), .A3(new_n671), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1355gat));
endmodule


