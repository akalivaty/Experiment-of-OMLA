//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n210));
  XNOR2_X1  g0010(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n207), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n224));
  AND3_X1   g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n221), .A2(new_n225), .B1(G1), .B2(G20), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT1), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n211), .B(new_n219), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(new_n227), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  AND2_X1   g0045(.A1(G1), .A2(G13), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n257), .A2(G223), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT66), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n254), .A2(G222), .A3(new_n261), .ZN(new_n262));
  MUX2_X1   g0062(.A(new_n260), .B(KEYINPUT66), .S(new_n262), .Z(new_n263));
  OAI21_X1  g0063(.A(new_n249), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n247), .ZN(new_n265));
  OAI21_X1  g0065(.A(G274), .B1(new_n265), .B2(new_n217), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n249), .A2(new_n269), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(G226), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G200), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT68), .B1(new_n276), .B2(new_n217), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n206), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G50), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n207), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G50), .A2(G58), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n207), .B1(new_n292), .B2(new_n213), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n280), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n285), .B(new_n294), .C1(G50), .C2(new_n281), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT9), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n275), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT69), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n274), .B2(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n264), .A2(KEYINPUT69), .A3(G190), .A4(new_n273), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n297), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n274), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n264), .A2(new_n310), .A3(new_n273), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n295), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n281), .A2(KEYINPUT70), .A3(G68), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT12), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT70), .B1(new_n281), .B2(G68), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n317), .ZN(new_n319));
  INV_X1    g0119(.A(G50), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n290), .A2(new_n320), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n287), .A2(new_n259), .B1(new_n207), .B2(G68), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n280), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT11), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n318), .B(new_n319), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n283), .A2(G68), .A3(new_n284), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n324), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n231), .A2(G1698), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n254), .B(new_n331), .C1(G226), .C2(G1698), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G97), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n249), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n271), .B1(G238), .B2(new_n272), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT13), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n248), .B1(new_n332), .B2(new_n333), .ZN(new_n339));
  INV_X1    g0139(.A(G274), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n246), .B2(new_n247), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n269), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n270), .A2(new_n248), .ZN(new_n343));
  INV_X1    g0143(.A(G238), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT13), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(G169), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n310), .B2(new_n347), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n347), .B2(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n330), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n347), .A2(G200), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n329), .C1(new_n299), .C2(new_n347), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G244), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n342), .B1(new_n343), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n254), .A2(G232), .A3(new_n261), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n203), .B2(new_n254), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n257), .B2(G238), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n358), .B1(new_n361), .B2(new_n248), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G190), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n283), .A2(G77), .A3(new_n284), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G20), .A2(G77), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT15), .B(G87), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n286), .B2(new_n290), .C1(new_n287), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n280), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n282), .A2(new_n259), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n364), .B(new_n372), .C1(new_n373), .C2(new_n363), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n362), .B2(new_n308), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n310), .B(new_n358), .C1(new_n361), .C2(new_n248), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n381), .B2(new_n207), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n253), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n207), .B1(new_n214), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT71), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n289), .A2(G159), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n390), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT71), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n385), .A2(KEYINPUT16), .A3(new_n391), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n252), .A2(new_n207), .A3(new_n253), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n213), .B1(new_n398), .B2(new_n383), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n388), .A2(new_n390), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n394), .A2(new_n280), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n286), .B1(new_n206), .B2(G20), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n283), .A2(new_n403), .B1(new_n282), .B2(new_n286), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n342), .B1(new_n343), .B2(new_n231), .ZN(new_n406));
  OR2_X1    g0206(.A1(G223), .A2(G1698), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n407), .B1(G226), .B2(new_n261), .C1(new_n379), .C2(new_n380), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n248), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G179), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n406), .B2(new_n410), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n405), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  INV_X1    g0218(.A(new_n406), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n408), .A2(new_n409), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n249), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n421), .A3(new_n299), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G200), .B2(new_n411), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(new_n402), .A3(new_n404), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n423), .A2(new_n402), .A3(KEYINPUT17), .A4(new_n404), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n416), .A2(new_n418), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  OR3_X1    g0228(.A1(new_n355), .A2(new_n378), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n313), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT73), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(new_n267), .A3(KEYINPUT5), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT5), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(KEYINPUT73), .B2(G41), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n268), .A2(G1), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n436), .A2(new_n248), .ZN(new_n437));
  OAI211_X1 g0237(.A(G264), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n438));
  INV_X1    g0238(.A(G257), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1698), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n379), .B2(new_n380), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n252), .A2(G303), .A3(new_n253), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n437), .A2(G270), .B1(new_n443), .B2(new_n249), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT74), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n436), .B2(new_n266), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n206), .A2(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT73), .A2(G41), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(KEYINPUT5), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n449), .A2(KEYINPUT74), .A3(new_n341), .A4(new_n434), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n373), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT79), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n276), .A2(new_n217), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT20), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n277), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n206), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(G116), .A3(new_n281), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n282), .A2(new_n457), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n463), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OR3_X1    g0270(.A1(new_n452), .A2(new_n453), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n453), .B1(new_n452), .B2(new_n470), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n444), .A2(new_n451), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n471), .B(new_n472), .C1(new_n299), .C2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(G169), .A3(new_n470), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT77), .B(KEYINPUT21), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT78), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n475), .A2(KEYINPUT78), .A3(new_n476), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT21), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT76), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n308), .B1(new_n444), .B2(new_n451), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT76), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT21), .A4(new_n470), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n470), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n436), .A2(G270), .A3(new_n248), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n443), .A2(new_n249), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n451), .A2(G179), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n474), .A2(new_n481), .A3(new_n487), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n207), .B1(new_n333), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G87), .B2(new_n204), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n287), .B2(new_n202), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n207), .B(G68), .C1(new_n379), .C2(new_n380), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(new_n280), .B1(new_n282), .B2(new_n367), .ZN(new_n500));
  INV_X1    g0300(.A(new_n367), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n466), .A2(new_n281), .A3(new_n501), .A4(new_n467), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n435), .A2(new_n340), .ZN(new_n504));
  INV_X1    g0304(.A(G250), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n447), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n248), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n344), .A2(new_n261), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n356), .A2(G1698), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n509), .C1(new_n379), .C2(new_n380), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n507), .B1(new_n512), .B2(new_n248), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n308), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n248), .B1(new_n510), .B2(new_n511), .ZN(new_n515));
  INV_X1    g0315(.A(new_n507), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n310), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n503), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(G200), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(G190), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n283), .A2(G87), .A3(new_n467), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n500), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G257), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  OAI21_X1  g0326(.A(G250), .B1(new_n379), .B2(new_n380), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n249), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n437), .A2(G264), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n451), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G179), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n308), .B2(new_n531), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n282), .A2(new_n203), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT25), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n466), .A2(new_n281), .A3(new_n467), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n535), .B1(new_n537), .B2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n539));
  NAND2_X1  g0339(.A1(KEYINPUT80), .A2(KEYINPUT24), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(new_n207), .A3(G107), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT23), .B1(new_n203), .B2(G20), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n539), .B(new_n540), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n254), .A2(new_n207), .A3(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT22), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n254), .A2(new_n547), .A3(new_n207), .A4(G87), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(KEYINPUT80), .A2(KEYINPUT24), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n280), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n550), .B(new_n544), .C1(new_n546), .C2(new_n548), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n538), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n524), .B1(new_n533), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g0355(.A(G97), .B(G107), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n557), .A2(new_n202), .A3(G107), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n207), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n289), .A2(G77), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT72), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n203), .B1(new_n398), .B2(new_n383), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n466), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n281), .A2(G97), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n536), .B2(new_n202), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT75), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n571), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n562), .B(KEYINPUT72), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n559), .B1(new_n557), .B2(new_n556), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n207), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n280), .B1(new_n576), .B2(new_n566), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT75), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(KEYINPUT4), .A2(G244), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n261), .B(new_n581), .C1(new_n379), .C2(new_n380), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n356), .B1(new_n252), .B2(new_n253), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n454), .C1(new_n583), .C2(KEYINPUT4), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n261), .B1(new_n527), .B2(KEYINPUT4), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n249), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n437), .A2(G257), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n451), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G169), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n446), .A2(new_n450), .B1(new_n437), .B2(G257), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(G179), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n580), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n568), .A2(new_n571), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(G190), .A3(new_n586), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n588), .A2(G200), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n549), .A2(new_n551), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n549), .A2(new_n551), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n280), .A3(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n451), .A2(new_n529), .A3(new_n530), .A4(G190), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n531), .A2(G200), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n600), .A2(new_n538), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n555), .A2(new_n593), .A3(new_n597), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n493), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n430), .A2(new_n605), .ZN(G372));
  INV_X1    g0406(.A(KEYINPUT83), .ZN(new_n607));
  INV_X1    g0407(.A(new_n307), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n416), .A2(new_n418), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n354), .A2(new_n376), .A3(new_n375), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n352), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n426), .A2(new_n427), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n607), .B(new_n312), .C1(new_n608), .C2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n304), .B2(new_n306), .ZN(new_n615));
  INV_X1    g0415(.A(new_n312), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT83), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT81), .B1(new_n513), .B2(new_n308), .ZN(new_n619));
  OAI211_X1 g0419(.A(KEYINPUT81), .B(new_n308), .C1(new_n515), .C2(new_n516), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n518), .B(new_n503), .C1(new_n619), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n602), .A2(new_n601), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n622), .B(new_n523), .C1(new_n554), .C2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n572), .A2(new_n579), .B1(new_n589), .B2(new_n591), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n594), .A2(new_n596), .A3(new_n595), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n475), .A2(KEYINPUT78), .A3(new_n476), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT78), .B1(new_n475), .B2(new_n476), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n492), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n483), .A2(new_n486), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT82), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT82), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n481), .A2(new_n634), .A3(new_n487), .A4(new_n492), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n532), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n531), .A2(new_n308), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n554), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n628), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n593), .B2(new_n524), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n622), .A2(new_n523), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n591), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n308), .B1(new_n590), .B2(new_n586), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(new_n568), .B2(new_n571), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n643), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n641), .A2(new_n649), .A3(new_n622), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n640), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n430), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n618), .A2(new_n652), .ZN(G369));
  NAND3_X1  g0453(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n488), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n633), .A2(new_n635), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n493), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n554), .A2(new_n659), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n603), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n639), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n639), .A2(new_n659), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT84), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n667), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n631), .A2(new_n632), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n659), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n668), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(G399));
  NAND2_X1  g0482(.A1(new_n208), .A2(new_n267), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n215), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n688), .B(new_n660), .C1(new_n640), .C2(new_n650), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT26), .B1(new_n642), .B2(new_n646), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n519), .A2(new_n523), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n580), .A3(new_n648), .A4(new_n592), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n692), .A3(new_n622), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT86), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n481), .A2(new_n487), .A3(new_n492), .A4(new_n639), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n627), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n690), .A2(new_n692), .A3(KEYINPUT86), .A4(new_n622), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n660), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n689), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n491), .A2(KEYINPUT85), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n586), .A2(new_n451), .A3(new_n587), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT85), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n444), .A2(new_n706), .A3(G179), .A4(new_n451), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n517), .A2(new_n529), .A3(new_n530), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n704), .A2(new_n705), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n517), .A2(G179), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n588), .A2(new_n473), .A3(new_n712), .A4(new_n531), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n705), .A2(KEYINPUT30), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n659), .B1(new_n711), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n605), .B2(new_n660), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n718), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n703), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n702), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT87), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n687), .B1(new_n724), .B2(G1), .ZN(G364));
  AND2_X1   g0525(.A1(new_n207), .A2(G13), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n206), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n683), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n663), .B2(G330), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G330), .B2(new_n663), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n217), .B1(G20), .B2(new_n308), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT90), .Z(new_n741));
  NAND2_X1  g0541(.A1(new_n381), .A2(new_n208), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n268), .B2(new_n216), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n241), .B2(new_n268), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n254), .A2(new_n208), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n746), .B1(G116), .B2(new_n208), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n747), .A2(KEYINPUT88), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(KEYINPUT88), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n744), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n730), .B1(new_n741), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G20), .A3(new_n299), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n254), .B1(new_n754), .B2(G329), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n207), .B1(new_n752), .B2(G190), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(G20), .A2(G179), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT33), .B(G317), .Z(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n207), .A2(new_n373), .A3(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G190), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT91), .ZN(new_n769));
  AOI21_X1  g0569(.A(G200), .B1(new_n759), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n769), .B2(new_n759), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n758), .B(new_n768), .C1(G311), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT92), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n774), .A2(new_n775), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G326), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(new_n299), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT93), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT93), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G283), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n771), .A2(new_n299), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G322), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n773), .A2(new_n781), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n753), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  INV_X1    g0593(.A(new_n767), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G87), .ZN(new_n795));
  INV_X1    g0595(.A(new_n757), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n762), .A2(G68), .B1(new_n796), .B2(G97), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n793), .A2(new_n254), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n780), .A2(G50), .B1(G77), .B2(new_n772), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n786), .A2(G107), .ZN(new_n800));
  INV_X1    g0600(.A(new_n788), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n799), .B(new_n800), .C1(new_n212), .C2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n790), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT94), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n736), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n803), .B2(new_n804), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n751), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n739), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n663), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n732), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NOR2_X1   g0612(.A1(new_n736), .A2(new_n737), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n729), .B(new_n728), .C1(new_n813), .C2(new_n259), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n786), .A2(G87), .ZN(new_n815));
  INV_X1    g0615(.A(new_n772), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n457), .B2(new_n816), .C1(new_n779), .C2(new_n765), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n801), .A2(new_n756), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n381), .B1(new_n753), .B2(new_n819), .C1(new_n202), .C2(new_n757), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n763), .A2(new_n821), .B1(new_n203), .B2(new_n767), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n817), .A2(new_n818), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G143), .A2(new_n788), .B1(new_n772), .B2(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n825), .B2(new_n779), .C1(new_n288), .C2(new_n763), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n254), .B1(new_n828), .B2(new_n753), .C1(new_n767), .C2(new_n320), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n785), .A2(new_n213), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(G58), .C2(new_n796), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n823), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n374), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT95), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n377), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n371), .A2(new_n659), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n377), .A2(new_n834), .A3(new_n836), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n814), .B1(new_n806), .B2(new_n832), .C1(new_n840), .C2(new_n738), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n651), .A2(new_n660), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n838), .A2(new_n839), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n374), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n660), .B(new_n840), .C1(new_n640), .C2(new_n650), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n722), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT96), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n847), .ZN(new_n850));
  INV_X1    g0650(.A(new_n722), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n730), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n842), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  NOR2_X1   g0654(.A1(new_n329), .A2(new_n660), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n352), .A2(new_n354), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT97), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n352), .A2(KEYINPUT97), .A3(new_n354), .A4(new_n856), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n350), .A2(new_n351), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n855), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n840), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT31), .B1(new_n717), .B2(KEYINPUT102), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n866), .B(new_n659), .C1(new_n711), .C2(new_n716), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT103), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n865), .A2(KEYINPUT103), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n864), .B1(new_n872), .B2(new_n720), .ZN(new_n873));
  INV_X1    g0673(.A(new_n404), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT98), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n391), .A2(new_n393), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n399), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n385), .A2(KEYINPUT98), .A3(new_n391), .A4(new_n393), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n395), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n394), .A2(new_n280), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n414), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n424), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n657), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n657), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n405), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n888));
  NAND4_X1  g0688(.A1(new_n415), .A2(new_n887), .A3(new_n424), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n428), .A2(KEYINPUT99), .A3(new_n884), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT99), .B1(new_n428), .B2(new_n884), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT38), .B(new_n890), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n895), .A2(KEYINPUT101), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT101), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n873), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n428), .A2(new_n405), .A3(new_n886), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n415), .A2(new_n887), .A3(new_n424), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(new_n888), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n894), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n900), .B1(new_n896), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n873), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n593), .A2(new_n597), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n603), .A2(new_n639), .A3(new_n691), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(new_n678), .A3(new_n474), .A4(new_n660), .ZN(new_n912));
  INV_X1    g0712(.A(new_n719), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n870), .B2(new_n871), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n915), .A2(new_n313), .A3(new_n429), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n908), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n908), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n917), .A2(new_n918), .A3(new_n703), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n377), .A2(new_n659), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n920), .B1(new_n847), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n897), .B2(new_n898), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n609), .A2(new_n657), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n896), .A2(new_n905), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n861), .A2(new_n330), .A3(new_n660), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n702), .A2(new_n430), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n618), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n919), .A2(new_n937), .B1(new_n206), .B2(new_n726), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n919), .ZN(new_n939));
  INV_X1    g0739(.A(new_n575), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT35), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT35), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n941), .A2(G116), .A3(new_n218), .A4(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT36), .Z(new_n944));
  NAND3_X1  g0744(.A1(new_n216), .A2(G77), .A3(new_n386), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n320), .A2(G68), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n206), .B(G13), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n939), .A2(new_n944), .A3(new_n947), .ZN(G367));
  INV_X1    g0748(.A(KEYINPUT105), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n593), .B(new_n597), .C1(new_n594), .C2(new_n660), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n647), .A2(new_n659), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n949), .B1(new_n677), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n676), .A2(KEYINPUT105), .A3(new_n952), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT106), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n680), .A2(new_n952), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n593), .B1(new_n953), .B2(new_n639), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n957), .A2(KEYINPUT42), .B1(new_n660), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n522), .A2(new_n500), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n659), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n643), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT104), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT104), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(new_n622), .C2(new_n962), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n958), .A2(new_n960), .B1(KEYINPUT43), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n954), .A2(KEYINPUT106), .A3(new_n955), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n956), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n968), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n967), .A2(new_n972), .ZN(new_n974));
  AND4_X1   g0774(.A1(new_n970), .A2(new_n973), .A3(new_n974), .A4(new_n956), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n683), .B(KEYINPUT41), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n674), .A2(new_n679), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n669), .A3(new_n952), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT107), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(KEYINPUT107), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n681), .B2(new_n952), .ZN(new_n987));
  OAI211_X1 g0787(.A(KEYINPUT44), .B(new_n953), .C1(new_n680), .C2(new_n668), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(new_n985), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n676), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n674), .A2(new_n679), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n680), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n664), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n984), .A2(new_n677), .A3(new_n985), .A4(new_n989), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n991), .A2(new_n724), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n977), .B1(new_n996), .B2(new_n724), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n976), .B1(new_n997), .B2(new_n728), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n740), .B1(new_n208), .B2(new_n367), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n237), .A2(new_n742), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n730), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT108), .Z(new_n1002));
  NAND3_X1  g0802(.A1(new_n794), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT46), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n767), .B2(new_n457), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(new_n756), .C2(new_n763), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(KEYINPUT110), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT109), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n779), .A2(new_n819), .B1(new_n801), .B2(new_n765), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n381), .B1(new_n753), .B2(new_n1012), .C1(new_n203), .C2(new_n757), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n786), .B2(G97), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1006), .A2(KEYINPUT110), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n821), .C2(new_n816), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT112), .B(G137), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n753), .A2(new_n1017), .B1(new_n757), .B2(new_n213), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n763), .A2(new_n791), .B1(new_n212), .B2(new_n767), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(G150), .C2(new_n788), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n780), .A2(G143), .B1(G50), .B2(new_n772), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n254), .B1(new_n785), .B2(new_n259), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1020), .B(new_n1021), .C1(new_n1022), .C2(KEYINPUT111), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1011), .A2(new_n1016), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT47), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n806), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1002), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n809), .B2(new_n966), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n998), .A2(new_n1030), .ZN(G387));
  OAI22_X1  g0831(.A1(new_n745), .A2(new_n684), .B1(G107), .B2(new_n208), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n234), .A2(new_n268), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n684), .ZN(new_n1034));
  AOI211_X1 g0834(.A(G45), .B(new_n1034), .C1(G68), .C2(G77), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n286), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n742), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1032), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n730), .B1(new_n1040), .B2(new_n741), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n757), .A2(new_n367), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n254), .B1(new_n288), .B2(new_n753), .C1(new_n767), .C2(new_n259), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n286), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1043), .C1(new_n1044), .C2(new_n762), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n786), .A2(G97), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n780), .A2(G159), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G50), .A2(new_n788), .B1(new_n772), .B2(G68), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n767), .A2(new_n756), .B1(new_n821), .B2(new_n757), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n780), .A2(G322), .B1(G303), .B2(new_n772), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n819), .B2(new_n763), .C1(new_n1012), .C2(new_n801), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n1053), .B2(new_n1052), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT49), .Z(new_n1056));
  AOI21_X1  g0856(.A(new_n254), .B1(new_n754), .B2(G326), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n785), .B2(new_n457), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1049), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1041), .B1(new_n1059), .B2(new_n736), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n674), .B2(new_n809), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT114), .Z(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n728), .B2(new_n994), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n724), .A2(new_n994), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n729), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n724), .A2(new_n994), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  NAND3_X1  g0867(.A1(new_n991), .A2(new_n728), .A3(new_n995), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n740), .B1(new_n202), .B2(new_n208), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n244), .A2(new_n742), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n730), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n779), .A2(new_n1012), .B1(new_n801), .B2(new_n819), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT52), .Z(new_n1073));
  NOR2_X1   g0873(.A1(new_n767), .A2(new_n821), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n254), .B(new_n1074), .C1(G322), .C2(new_n754), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n772), .A2(G294), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n762), .A2(G303), .B1(new_n796), .B2(G116), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n800), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n779), .A2(new_n288), .B1(new_n801), .B2(new_n791), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT51), .Z(new_n1080));
  NOR2_X1   g0880(.A1(new_n767), .A2(new_n213), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n381), .B(new_n1081), .C1(G143), .C2(new_n754), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n772), .A2(new_n1044), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n762), .A2(G50), .B1(new_n796), .B2(G77), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n815), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1073), .A2(new_n1078), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1071), .B1(new_n1086), .B2(new_n736), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n952), .B2(new_n809), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n996), .A2(new_n729), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n991), .A2(new_n995), .B1(new_n724), .B2(new_n994), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1068), .B(new_n1088), .C1(new_n1089), .C2(new_n1090), .ZN(G390));
  NAND3_X1  g0891(.A1(new_n699), .A2(new_n840), .A3(new_n660), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n920), .B1(new_n1092), .B2(new_n922), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n928), .A2(new_n932), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT115), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n932), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n896), .B2(new_n905), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n694), .A2(new_n693), .B1(new_n696), .B2(new_n627), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n659), .B1(new_n1099), .B2(new_n698), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n921), .B1(new_n1100), .B2(new_n840), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1096), .B(new_n1098), .C1(new_n1101), .C2(new_n920), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1095), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n931), .B1(new_n923), .B2(new_n1097), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n915), .A2(new_n703), .A3(new_n864), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n722), .A2(new_n840), .A3(new_n863), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1103), .A2(new_n1104), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n728), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT116), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1107), .A2(new_n1112), .A3(new_n728), .A4(new_n1109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1109), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1106), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n915), .A2(new_n703), .A3(new_n845), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1108), .B(new_n1101), .C1(new_n1118), .C2(new_n863), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n847), .A2(new_n922), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n863), .B1(new_n722), .B2(new_n840), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1106), .B2(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n717), .A2(KEYINPUT102), .ZN(new_n1124));
  AND4_X1   g0924(.A1(KEYINPUT103), .A2(new_n1124), .A3(new_n718), .A4(new_n867), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT103), .B1(new_n865), .B2(new_n867), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n720), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n430), .A2(new_n1127), .A3(G330), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n935), .A2(new_n618), .A3(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n1115), .A2(new_n1117), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1107), .A2(new_n1109), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n729), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n931), .A2(new_n737), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n813), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n730), .B1(new_n1135), .B2(new_n1044), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n780), .A2(G128), .B1(G132), .B2(new_n788), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n767), .A2(new_n288), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n1139), .C1(new_n320), .C2(new_n785), .ZN(new_n1140));
  INV_X1    g0940(.A(G125), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n254), .B1(new_n753), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G159), .B2(new_n796), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1143), .B1(new_n763), .B2(new_n1017), .C1(new_n816), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n830), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n254), .B1(new_n754), .B2(G294), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n762), .A2(G107), .B1(new_n796), .B2(G77), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1146), .A2(new_n795), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n780), .A2(G283), .B1(G97), .B2(new_n772), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n457), .B2(new_n801), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1140), .A2(new_n1145), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1136), .B1(new_n1152), .B2(new_n736), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1134), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1114), .A2(new_n1133), .A3(new_n1154), .ZN(G378));
  OR2_X1    g0955(.A1(new_n925), .A2(new_n933), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n295), .A2(new_n886), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n313), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n306), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n305), .B1(new_n297), .B2(new_n302), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n312), .B(new_n1157), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1162), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1157), .B1(new_n307), .B2(new_n312), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n703), .B1(new_n873), .B2(new_n906), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n901), .B2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n857), .A2(new_n858), .B1(new_n861), .B2(new_n855), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n845), .B1(new_n860), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1127), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT101), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n428), .A2(new_n884), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT99), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n428), .A2(KEYINPUT99), .A3(new_n884), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT38), .B1(new_n1180), .B2(new_n890), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n896), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1175), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n895), .A2(KEYINPUT101), .A3(new_n896), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1174), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1170), .B(new_n1169), .C1(new_n1185), .C2(KEYINPUT40), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1156), .B1(new_n1171), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1169), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT40), .B1(new_n1190), .B2(new_n873), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1170), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n934), .A3(new_n1186), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1129), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1132), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1197), .A3(KEYINPUT57), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1194), .A2(new_n1188), .B1(new_n1132), .B2(new_n1196), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n729), .C1(KEYINPUT57), .C2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1144), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n794), .A2(new_n1201), .B1(new_n796), .B2(G150), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n828), .B2(new_n763), .ZN(new_n1203));
  INV_X1    g1003(.A(G128), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1204), .A2(new_n801), .B1(new_n816), .B2(new_n825), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G125), .C2(new_n780), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n786), .A2(G159), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n786), .A2(G58), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n203), .B2(new_n801), .C1(new_n779), .C2(new_n457), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n816), .A2(new_n367), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n254), .A2(G41), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n213), .B2(new_n757), .C1(new_n821), .C2(new_n753), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n763), .A2(new_n202), .B1(new_n259), .B2(new_n767), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT58), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1216), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n320), .C1(G33), .C2(G41), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1219), .A2(KEYINPUT58), .ZN(new_n1223));
  AND4_X1   g1023(.A1(new_n1212), .A2(new_n1220), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n730), .B1(G50), .B2(new_n1135), .C1(new_n1224), .C2(new_n806), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1189), .B2(new_n737), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1195), .B2(new_n728), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1200), .A2(new_n1227), .ZN(G375));
  OAI21_X1  g1028(.A(new_n730), .B1(new_n1135), .B2(G68), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n381), .B1(new_n753), .B2(new_n765), .C1(new_n763), .C2(new_n457), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G97), .B2(new_n794), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n780), .A2(G294), .B1(G107), .B2(new_n772), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(new_n259), .C2(new_n785), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1042), .B1(new_n788), .B2(G283), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT117), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n780), .A2(G132), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT118), .Z(new_n1237));
  OAI21_X1  g1037(.A(new_n254), .B1(new_n753), .B2(new_n1204), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n763), .A2(new_n1144), .B1(new_n320), .B2(new_n757), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(G159), .C2(new_n794), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1017), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G150), .A2(new_n772), .B1(new_n788), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1213), .A3(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1233), .A2(new_n1235), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT119), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n806), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1229), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n738), .B2(new_n863), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1123), .B2(new_n727), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1131), .A2(new_n977), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1119), .A2(new_n1129), .A3(new_n1122), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(G381));
  OR3_X1    g1055(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(G387), .A2(new_n1256), .A3(G384), .A4(G390), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1257), .B(KEYINPUT120), .Z(new_n1258));
  INV_X1    g1058(.A(G378), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1200), .A2(new_n1259), .A3(new_n1227), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1258), .A2(new_n1260), .ZN(G407));
  OAI211_X1 g1061(.A(G407), .B(G213), .C1(G343), .C2(new_n1260), .ZN(G409));
  AND2_X1   g1062(.A1(new_n658), .A2(G213), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1193), .A2(new_n934), .A3(new_n1186), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n934), .B1(new_n1193), .B2(new_n1186), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT57), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1132), .A2(new_n1196), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n729), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G378), .B(new_n1227), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT121), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1200), .A2(KEYINPUT121), .A3(G378), .A4(new_n1227), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n977), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1227), .A2(KEYINPUT122), .B1(new_n1275), .B2(new_n1199), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT122), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n727), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n1226), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G378), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1263), .B1(new_n1274), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1250), .B1(new_n853), .B2(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1253), .A2(KEYINPUT123), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1131), .A2(new_n683), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1285), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n853), .A2(new_n1284), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n1285), .B1(new_n1284), .B2(new_n853), .C1(new_n1288), .C2(new_n1290), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1263), .A2(G2897), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1280), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(new_n1301), .B2(new_n1263), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1283), .A2(new_n1299), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(G390), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT126), .B1(G387), .B2(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(G393), .B(new_n811), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G390), .B1(new_n998), .B2(new_n1030), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n998), .A2(new_n1030), .A3(G390), .ZN(new_n1309));
  OAI22_X1  g1109(.A1(new_n1305), .A2(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1308), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n998), .A2(new_n1030), .A3(G390), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1311), .A2(KEYINPUT126), .A3(new_n1312), .A4(new_n1306), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1314), .A2(KEYINPUT61), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1282), .A2(new_n1316), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1317), .A2(KEYINPUT63), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(KEYINPUT63), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1303), .B(new_n1315), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT62), .B1(new_n1282), .B2(new_n1316), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1316), .ZN(new_n1323));
  NOR4_X1   g1123(.A1(new_n1301), .A2(new_n1322), .A3(new_n1323), .A4(new_n1263), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1299), .B1(new_n1301), .B2(new_n1263), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1326), .A2(KEYINPUT127), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT127), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1325), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1314), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1320), .B1(new_n1330), .B2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1259), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1274), .A2(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1314), .B(new_n1334), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1335), .B(new_n1316), .ZN(G402));
endmodule


