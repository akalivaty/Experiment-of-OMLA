//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069;
  XOR2_X1   g000(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n187), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT66), .A2(G134), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT66), .A2(G134), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n197), .B(new_n198), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(G134), .B2(new_n198), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n199), .A2(new_n200), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G137), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n196), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT66), .A2(G134), .ZN(new_n212));
  AOI21_X1  g026(.A(G137), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n202), .B1(new_n213), .B2(new_n197), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n196), .B1(new_n215), .B2(new_n198), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n208), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(G131), .B1(new_n205), .B2(G137), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n204), .A2(new_n218), .A3(KEYINPUT67), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n207), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  AND2_X1   g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(KEYINPUT64), .A2(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT64), .A2(G143), .ZN(new_n226));
  AOI21_X1  g040(.A(G146), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n224), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(G146), .A3(new_n226), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G146), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(KEYINPUT65), .A3(G143), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n231), .A2(new_n234), .A3(new_n235), .A4(new_n222), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n220), .A2(new_n221), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n204), .A2(new_n206), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n204), .A2(new_n218), .A3(KEYINPUT67), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n204), .B2(new_n218), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n230), .A2(new_n236), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT68), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n233), .B2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n227), .B2(new_n229), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n231), .A2(new_n234), .A3(new_n235), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n213), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n210), .A2(G137), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n196), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n217), .B2(new_n219), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(KEYINPUT69), .ZN(new_n257));
  INV_X1    g071(.A(new_n255), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n241), .B2(new_n242), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n238), .A2(new_n245), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT71), .B(G116), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G119), .ZN(new_n264));
  INV_X1    g078(.A(G116), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G119), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G113), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT2), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G113), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n264), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(KEYINPUT70), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n269), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n266), .B1(new_n263), .B2(G119), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n262), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n243), .B2(new_n244), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n258), .B(new_n252), .C1(new_n241), .C2(new_n242), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n217), .A2(new_n219), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(KEYINPUT72), .A3(new_n258), .A4(new_n252), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n195), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT28), .B1(new_n281), .B2(new_n282), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n194), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n243), .A2(new_n244), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n284), .A2(new_n286), .A3(new_n291), .A4(KEYINPUT30), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n221), .B1(new_n220), .B2(new_n237), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n243), .A2(KEYINPUT68), .A3(new_n244), .ZN(new_n294));
  INV_X1    g108(.A(new_n252), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n259), .B2(new_n260), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n285), .A2(KEYINPUT69), .A3(new_n258), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n293), .A2(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n279), .B(new_n292), .C1(new_n298), .C2(KEYINPUT30), .ZN(new_n299));
  INV_X1    g113(.A(new_n287), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(new_n194), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT31), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT31), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n299), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n290), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT74), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n309), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n289), .A2(new_n194), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT29), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n284), .A2(new_n286), .A3(new_n291), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n279), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n195), .B1(new_n319), .B2(new_n287), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n315), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n323));
  INV_X1    g137(.A(new_n316), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n288), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n193), .B1(new_n299), .B2(new_n287), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n314), .B1(new_n327), .B2(G472), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n293), .A2(new_n294), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n259), .A2(new_n260), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n297), .A3(new_n252), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT30), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n279), .ZN(new_n333));
  INV_X1    g147(.A(new_n292), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n194), .B1(new_n335), .B2(new_n300), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n333), .B1(new_n329), .B2(new_n331), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT28), .B1(new_n337), .B2(new_n300), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n338), .B2(new_n316), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n321), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G472), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n340), .A2(KEYINPUT75), .A3(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n312), .B(new_n313), .C1(new_n328), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n344));
  INV_X1    g158(.A(G119), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(G128), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n249), .A2(KEYINPUT76), .A3(G119), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n346), .B(new_n347), .C1(G119), .C2(new_n249), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT24), .B(G110), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n350), .B(KEYINPUT77), .Z(new_n351));
  INV_X1    g165(.A(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G125), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(KEYINPUT16), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G140), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n352), .A2(G125), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n358), .B2(KEYINPUT16), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n359), .A2(G146), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(G146), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT78), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n345), .A2(KEYINPUT79), .A3(G128), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT23), .B1(new_n249), .B2(G119), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n345), .B2(G128), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n364), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G110), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n351), .A2(new_n362), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n359), .A2(G146), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n355), .A2(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n353), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT80), .B1(new_n374), .B2(G146), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n353), .A2(new_n373), .A3(new_n376), .A4(new_n228), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n348), .A2(new_n349), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n369), .B2(G110), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT81), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT81), .B1(new_n379), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n371), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT22), .B(G137), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n385), .B(new_n386), .Z(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n371), .B(new_n387), .C1(new_n382), .C2(new_n383), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n315), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT25), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n389), .A2(KEYINPUT25), .A3(new_n315), .A4(new_n390), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G217), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(G234), .B2(new_n315), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(G902), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT82), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n389), .A2(new_n401), .A3(new_n390), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n225), .A2(KEYINPUT13), .A3(G128), .A4(new_n226), .ZN(new_n406));
  AND2_X1   g220(.A1(KEYINPUT64), .A2(G143), .ZN(new_n407));
  NOR2_X1   g221(.A1(KEYINPUT64), .A2(G143), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n407), .A2(new_n408), .A3(new_n249), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n233), .A2(G128), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT13), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(KEYINPUT94), .B(new_n406), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n225), .A2(G128), .A3(new_n226), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT94), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n414), .B(new_n415), .C1(new_n411), .C2(new_n410), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n413), .A2(new_n416), .A3(G134), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n414), .B(new_n205), .C1(G128), .C2(new_n233), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT71), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G116), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n419), .A2(new_n421), .A3(G122), .ZN(new_n422));
  INV_X1    g236(.A(G122), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT93), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT93), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G122), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n265), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n422), .A2(new_n427), .A3(G107), .ZN(new_n428));
  INV_X1    g242(.A(G107), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n425), .A2(G122), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n423), .A2(KEYINPUT93), .ZN(new_n431));
  OAI21_X1  g245(.A(G116), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n419), .A2(new_n421), .A3(G122), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n418), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n405), .B1(new_n417), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n413), .A2(G134), .A3(new_n416), .ZN(new_n437));
  OAI21_X1  g251(.A(G107), .B1(new_n422), .B2(new_n427), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n429), .A3(new_n433), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n437), .A2(KEYINPUT95), .A3(new_n440), .A4(new_n418), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT14), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n432), .B1(new_n422), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n444));
  OAI21_X1  g258(.A(G107), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n215), .B1(new_n409), .B2(new_n410), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n418), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n436), .A2(new_n441), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT9), .B(G234), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(new_n396), .A3(G953), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n436), .A2(new_n441), .A3(new_n448), .A4(new_n451), .ZN(new_n454));
  AOI21_X1  g268(.A(G902), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT96), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n456), .ZN(new_n458));
  INV_X1    g272(.A(G478), .ZN(new_n459));
  OAI22_X1  g273(.A1(new_n457), .A2(new_n458), .B1(KEYINPUT15), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n456), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT15), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(G478), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G113), .B(G122), .ZN(new_n465));
  INV_X1    g279(.A(G104), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n356), .B2(new_n357), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n353), .A2(new_n373), .A3(KEYINPUT88), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT19), .A3(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n374), .A2(KEYINPUT19), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n228), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n372), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n188), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT64), .B(G143), .ZN(new_n478));
  INV_X1    g292(.A(G214), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n479), .A2(G237), .A3(G953), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n476), .B1(new_n481), .B2(G131), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n225), .A3(new_n226), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT90), .B(new_n196), .C1(new_n484), .C2(new_n477), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n196), .A3(new_n477), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n475), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(KEYINPUT18), .A2(G131), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n481), .B(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n470), .A2(G146), .A3(new_n471), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n378), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n378), .A2(KEYINPUT89), .A3(new_n491), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n468), .B1(new_n488), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n481), .A2(G131), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT90), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n481), .A2(new_n476), .A3(G131), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n499), .A2(new_n487), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n360), .A2(new_n361), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT17), .B1(new_n482), .B2(new_n485), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n490), .ZN(new_n506));
  INV_X1    g320(.A(new_n495), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT89), .B1(new_n378), .B2(new_n491), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n509), .A3(new_n467), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n497), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(G475), .A2(G902), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(KEYINPUT92), .B2(KEYINPUT20), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n512), .A2(KEYINPUT92), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n505), .A2(new_n509), .A3(new_n467), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n499), .A2(new_n501), .A3(new_n487), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n372), .A3(new_n474), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n467), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n516), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n497), .A2(new_n510), .A3(KEYINPUT91), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n512), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n515), .B1(new_n523), .B2(KEYINPUT20), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n505), .A2(new_n509), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n468), .ZN(new_n526));
  AOI21_X1  g340(.A(G902), .B1(new_n526), .B2(new_n510), .ZN(new_n527));
  INV_X1    g341(.A(G475), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n189), .A2(G952), .ZN(new_n531));
  INV_X1    g345(.A(G234), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n188), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n315), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT21), .B(G898), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n530), .A2(new_n538), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n464), .A2(new_n524), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G214), .B1(G237), .B2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G210), .B1(G237), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT3), .B1(new_n466), .B2(G107), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT3), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n429), .A3(G104), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n466), .A2(G107), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G101), .ZN(new_n550));
  INV_X1    g364(.A(G101), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n545), .A2(new_n547), .A3(new_n551), .A4(new_n548), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(KEYINPUT4), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT4), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n549), .A2(new_n554), .A3(G101), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n279), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n264), .A2(KEYINPUT5), .A3(new_n267), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT5), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n268), .B1(new_n266), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n466), .A2(G107), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n429), .A2(G104), .ZN(new_n562));
  OAI21_X1  g376(.A(G101), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n552), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n273), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n556), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G110), .B(G122), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n556), .A2(new_n566), .A3(new_n568), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n570), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(KEYINPUT6), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n568), .B1(new_n556), .B2(new_n566), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT6), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n567), .A2(new_n576), .A3(new_n569), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT86), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n572), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n237), .A2(G125), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(G125), .B2(new_n252), .ZN(new_n582));
  INV_X1    g396(.A(G224), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(G953), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n582), .B(new_n584), .Z(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(KEYINPUT87), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT7), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n582), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n568), .B(KEYINPUT8), .ZN(new_n591));
  INV_X1    g405(.A(new_n566), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n565), .B1(new_n560), .B2(new_n273), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n571), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n595), .A2(new_n315), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n587), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n578), .B(new_n577), .C1(new_n573), .C2(new_n574), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n585), .B1(new_n598), .B2(new_n572), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(KEYINPUT87), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n544), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n580), .A2(new_n586), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT87), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(new_n543), .A3(new_n587), .A4(new_n596), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n542), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n540), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G221), .B1(new_n450), .B2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G469), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n315), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT85), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n244), .A2(new_n553), .A3(new_n555), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n552), .A2(new_n563), .A3(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n252), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT1), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n478), .B2(new_n228), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n618), .B2(new_n249), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n564), .B1(new_n619), .B2(new_n251), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n613), .B(new_n615), .C1(KEYINPUT10), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT83), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n243), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n285), .A2(KEYINPUT83), .A3(new_n240), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(G110), .B(G140), .ZN(new_n626));
  INV_X1    g440(.A(G227), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(G953), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n612), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT12), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n248), .A2(new_n564), .A3(new_n251), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n620), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n631), .B1(new_n634), .B2(new_n220), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n228), .B1(new_n407), .B2(new_n408), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT1), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n234), .A2(new_n235), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n637), .A2(G128), .B1(new_n638), .B2(new_n231), .ZN(new_n639));
  INV_X1    g453(.A(new_n251), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n565), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n632), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(KEYINPUT12), .A3(new_n243), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n623), .A2(new_n624), .ZN(new_n645));
  INV_X1    g459(.A(new_n553), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n230), .A2(new_n555), .A3(new_n236), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n615), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n249), .B1(new_n636), .B2(KEYINPUT1), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n251), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT10), .B1(new_n651), .B2(new_n565), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n629), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT85), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n630), .A2(new_n644), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n653), .A2(new_n220), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n629), .B1(new_n625), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n611), .B1(new_n659), .B2(new_n610), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT84), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n625), .A2(new_n657), .A3(new_n629), .ZN(new_n662));
  INV_X1    g476(.A(new_n629), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n645), .A2(new_n653), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n644), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n661), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n634), .A2(new_n631), .A3(new_n220), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT12), .B1(new_n642), .B2(new_n243), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n629), .B1(new_n669), .B2(new_n625), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n654), .B1(new_n220), .B2(new_n653), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(KEYINPUT84), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G469), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n609), .B1(new_n660), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n343), .A2(new_n404), .A3(new_n607), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G101), .ZN(G3));
  NAND2_X1  g491(.A1(new_n606), .A2(new_n538), .ZN(new_n678));
  INV_X1    g492(.A(new_n515), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n497), .A2(KEYINPUT91), .A3(new_n510), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT91), .B1(new_n497), .B2(new_n510), .ZN(new_n681));
  INV_X1    g495(.A(new_n512), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT20), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n530), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n459), .A2(G902), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT33), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n453), .A2(new_n688), .A3(new_n454), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n688), .B1(new_n453), .B2(new_n454), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n455), .A2(G478), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n678), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n675), .A2(new_n404), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n341), .B1(new_n306), .B2(new_n315), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n309), .B2(new_n306), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT34), .B(G104), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G6));
  NOR2_X1   g515(.A1(new_n683), .A2(new_n684), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n523), .A2(KEYINPUT20), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT97), .ZN(new_n704));
  OR3_X1    g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n539), .B1(new_n460), .B2(new_n463), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n704), .B1(new_n702), .B2(new_n703), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT98), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT98), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n705), .A2(new_n706), .A3(new_n710), .A4(new_n707), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n606), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n698), .A3(new_n696), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT35), .B(G107), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G9));
  OR3_X1    g530(.A1(new_n384), .A2(KEYINPUT36), .A3(new_n388), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n384), .B1(KEYINPUT36), .B2(new_n388), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n398), .B1(new_n400), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n675), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n607), .A3(new_n698), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT37), .B(G110), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G12));
  NAND2_X1  g538(.A1(new_n675), .A2(new_n720), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n309), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT32), .B1(new_n306), .B2(new_n309), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n327), .A2(new_n314), .A3(G472), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT75), .B1(new_n340), .B2(new_n341), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n725), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n535), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n533), .B1(new_n733), .B2(G900), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n705), .A2(new_n530), .A3(new_n707), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n606), .ZN(new_n736));
  INV_X1    g550(.A(new_n464), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G128), .ZN(G30));
  XNOR2_X1  g554(.A(new_n734), .B(KEYINPUT39), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n675), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT40), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(KEYINPUT99), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(KEYINPUT99), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n335), .A2(new_n300), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n194), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n319), .A2(new_n287), .A3(new_n194), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n315), .ZN(new_n749));
  OAI21_X1  g563(.A(G472), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n312), .A2(new_n313), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n720), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n601), .A2(new_n605), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT38), .Z(new_n755));
  NOR2_X1   g569(.A1(new_n524), .A2(new_n529), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n755), .A2(new_n542), .A3(new_n737), .A4(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n744), .A2(new_n745), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n478), .ZN(G45));
  NAND4_X1  g573(.A1(new_n686), .A2(KEYINPUT100), .A3(new_n693), .A4(new_n734), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n693), .B(new_n734), .C1(new_n524), .C2(new_n529), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT100), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n763), .A3(new_n606), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT101), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n760), .A2(new_n763), .A3(new_n606), .A4(KEYINPUT101), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n343), .A3(new_n721), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT102), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT102), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n732), .A2(new_n770), .A3(new_n766), .A4(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G146), .ZN(G48));
  AOI21_X1  g587(.A(new_n403), .B1(new_n728), .B2(new_n731), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n656), .A2(new_n658), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n315), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT103), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(G469), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n659), .B1(KEYINPUT103), .B2(new_n610), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n608), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n774), .A2(new_n695), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT41), .B(G113), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G15));
  NAND3_X1  g598(.A1(new_n343), .A2(new_n404), .A3(new_n781), .ZN(new_n785));
  OR3_X1    g599(.A1(new_n785), .A2(new_n712), .A3(KEYINPUT104), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT104), .B1(new_n785), .B2(new_n712), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G116), .ZN(G18));
  NOR2_X1   g603(.A1(new_n736), .A2(new_n780), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n343), .A2(new_n540), .A3(new_n790), .A4(new_n720), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G119), .ZN(G21));
  AOI21_X1  g606(.A(new_n542), .B1(new_n460), .B2(new_n463), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n754), .A2(new_n686), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n780), .A3(new_n537), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n194), .B1(new_n320), .B2(new_n289), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n303), .A2(new_n305), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n697), .B1(new_n309), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n404), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G122), .ZN(G24));
  NAND2_X1  g614(.A1(new_n760), .A2(new_n763), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n309), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n299), .A2(new_n304), .A3(new_n301), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n304), .B1(new_n299), .B2(new_n301), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(G902), .B1(new_n805), .B2(new_n290), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n720), .B(new_n802), .C1(new_n806), .C2(new_n341), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT105), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n697), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(KEYINPUT105), .A3(new_n720), .A4(new_n802), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n801), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n790), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G125), .ZN(G27));
  XNOR2_X1  g628(.A(new_n727), .B(KEYINPUT111), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n731), .A3(new_n313), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n643), .A2(new_n635), .B1(new_n645), .B2(new_n653), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT106), .B1(new_n817), .B2(new_n663), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT106), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n629), .C1(new_n669), .C2(new_n625), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n820), .A3(G469), .A4(new_n671), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT107), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n609), .B1(new_n822), .B2(new_n660), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n601), .A2(new_n541), .A3(new_n605), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT108), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n601), .A2(new_n605), .A3(KEYINPUT108), .A4(new_n541), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n801), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(KEYINPUT42), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n816), .A2(new_n404), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n828), .A2(new_n343), .A3(new_n404), .A4(new_n829), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(KEYINPUT109), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n774), .A2(new_n834), .A3(new_n828), .A4(new_n829), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n831), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G131), .ZN(G33));
  NOR2_X1   g653(.A1(new_n735), .A2(new_n737), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n774), .A2(new_n840), .A3(new_n828), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G134), .ZN(G36));
  NAND2_X1  g656(.A1(new_n756), .A2(new_n693), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT43), .Z(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n720), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT44), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n845), .A2(new_n846), .A3(new_n698), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n826), .A2(new_n827), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n673), .A2(KEYINPUT45), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n818), .A2(new_n820), .A3(KEYINPUT45), .A4(new_n671), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(G469), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n850), .A2(new_n852), .B1(new_n610), .B2(new_n315), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT46), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n853), .A2(new_n854), .B1(new_n610), .B2(new_n659), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n856), .A2(new_n608), .A3(new_n741), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n846), .B1(new_n845), .B2(new_n698), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n847), .A2(new_n849), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(G137), .ZN(G39));
  NOR4_X1   g674(.A1(new_n343), .A2(new_n848), .A3(new_n404), .A4(new_n801), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n608), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT47), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT47), .B1(new_n856), .B2(new_n608), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(G140), .ZN(G42));
  AND2_X1   g681(.A1(new_n816), .A2(new_n404), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n848), .A2(new_n780), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n869), .A2(new_n534), .A3(new_n844), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT48), .Z(new_n872));
  AND4_X1   g686(.A1(new_n404), .A2(new_n844), .A3(new_n534), .A4(new_n798), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n790), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n404), .A2(new_n869), .A3(new_n534), .A4(new_n752), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n531), .B(new_n874), .C1(new_n876), .C2(new_n694), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(new_n686), .A3(new_n693), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n755), .A2(new_n542), .A3(new_n781), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(KEYINPUT118), .A3(KEYINPUT50), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n873), .B2(new_n879), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n878), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n864), .A2(new_n865), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n778), .A2(new_n779), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n608), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n849), .B(new_n873), .C1(new_n885), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n809), .A2(new_n811), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n870), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT119), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n872), .B(new_n877), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  INV_X1    g709(.A(new_n695), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n799), .B(new_n791), .C1(new_n785), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n786), .B2(new_n787), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n889), .A2(new_n829), .A3(new_n828), .ZN(new_n899));
  INV_X1    g713(.A(new_n458), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n900), .A2(new_n461), .B1(new_n462), .B2(G478), .ZN(new_n901));
  INV_X1    g715(.A(new_n463), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT112), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT112), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n460), .A2(new_n904), .A3(new_n463), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n848), .A2(new_n735), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n732), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n899), .A2(new_n841), .A3(new_n908), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n542), .B(new_n537), .C1(new_n601), .C2(new_n605), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT113), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n906), .A2(new_n910), .A3(new_n911), .A4(new_n756), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n903), .A2(new_n756), .A3(new_n905), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT113), .B1(new_n678), .B2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n914), .A3(new_n698), .A4(new_n696), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n915), .A2(new_n676), .A3(new_n699), .A4(new_n722), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n909), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n838), .A2(new_n898), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT52), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n812), .A2(new_n790), .B1(new_n732), .B2(new_n738), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n734), .B(KEYINPUT114), .Z(new_n921));
  NAND4_X1  g735(.A1(new_n754), .A2(new_n793), .A3(new_n686), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n720), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n751), .A2(new_n923), .A3(new_n924), .A4(new_n823), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT115), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n822), .A2(new_n660), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n608), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n922), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(KEYINPUT115), .A3(new_n924), .A4(new_n751), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n772), .A2(new_n919), .A3(new_n920), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n772), .A2(new_n920), .A3(new_n932), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n918), .A2(KEYINPUT53), .A3(new_n933), .A4(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n938));
  NAND4_X1  g752(.A1(new_n933), .A2(new_n838), .A3(new_n898), .A4(new_n917), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n934), .A2(KEYINPUT52), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT54), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n838), .A2(new_n933), .A3(new_n898), .A4(new_n917), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT53), .B1(new_n944), .B2(new_n936), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n939), .A2(new_n940), .A3(new_n938), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n943), .B1(new_n947), .B2(new_n942), .ZN(new_n948));
  OAI22_X1  g762(.A1(new_n895), .A2(new_n948), .B1(G952), .B2(G953), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n886), .A2(KEYINPUT49), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n886), .A2(KEYINPUT49), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n404), .A2(new_n541), .A3(new_n608), .ZN(new_n952));
  NOR4_X1   g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .A4(new_n843), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n752), .A3(new_n755), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n949), .A2(new_n954), .ZN(G75));
  NOR2_X1   g769(.A1(new_n189), .A2(G952), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n315), .B1(new_n937), .B2(new_n941), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT56), .B1(new_n958), .B2(G210), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n580), .A2(new_n586), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(new_n599), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT55), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n957), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n959), .B2(new_n962), .ZN(G51));
  OR2_X1    g778(.A1(new_n850), .A2(new_n852), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n958), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT120), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n611), .B(KEYINPUT57), .ZN(new_n970));
  INV_X1    g784(.A(new_n943), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n942), .B1(new_n937), .B2(new_n941), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n775), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n956), .B1(new_n969), .B2(new_n974), .ZN(G54));
  INV_X1    g789(.A(KEYINPUT122), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n680), .A2(new_n681), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(KEYINPUT58), .A2(G475), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n938), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n934), .A2(KEYINPUT52), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n944), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n934), .A2(new_n935), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT53), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n939), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(G902), .B(new_n980), .C1(new_n983), .C2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT121), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n958), .A2(KEYINPUT121), .A3(new_n980), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n315), .B(new_n979), .C1(new_n937), .C2(new_n941), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n957), .B1(new_n992), .B2(new_n977), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n976), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n937), .A2(new_n941), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n995), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n956), .B1(new_n996), .B2(new_n978), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n997), .A2(KEYINPUT122), .A3(new_n989), .A4(new_n990), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n994), .A2(new_n998), .ZN(G60));
  OR2_X1    g813(.A1(new_n689), .A2(new_n690), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G478), .A2(G902), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT59), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1000), .B(new_n1002), .C1(new_n971), .C2(new_n972), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n957), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1000), .B1(new_n948), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(G63));
  NAND2_X1  g820(.A1(G217), .A2(G902), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT60), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n937), .B2(new_n941), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n389), .A2(new_n390), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1009), .A2(new_n717), .A3(new_n718), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1012), .A2(new_n957), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT61), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1012), .A2(KEYINPUT61), .A3(new_n957), .A4(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G66));
  OAI21_X1  g832(.A(G953), .B1(new_n536), .B2(new_n583), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(KEYINPUT123), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n897), .B(new_n916), .C1(new_n786), .C2(new_n787), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(G953), .ZN(new_n1022));
  MUX2_X1   g836(.A(new_n1020), .B(KEYINPUT123), .S(new_n1022), .Z(new_n1023));
  OAI211_X1 g837(.A(new_n598), .B(new_n572), .C1(G898), .C2(new_n189), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT124), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1023), .B(new_n1025), .ZN(G69));
  NAND2_X1  g840(.A1(new_n859), .A2(new_n866), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n742), .B1(new_n694), .B2(new_n913), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1028), .A2(new_n774), .A3(new_n849), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n772), .A2(new_n920), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n758), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT62), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1031), .A2(new_n1034), .A3(new_n758), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1030), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(KEYINPUT125), .ZN(new_n1037));
  OR2_X1    g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n332), .A2(new_n334), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n472), .A2(new_n473), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1040), .A2(new_n189), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(G900), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1045), .B1(new_n1043), .B2(new_n627), .ZN(new_n1046));
  INV_X1    g860(.A(new_n794), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n868), .A2(new_n1047), .A3(new_n857), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(new_n841), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n1027), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1050), .A2(new_n838), .A3(new_n1031), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n1051), .A2(new_n189), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1043), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1053), .B1(G227), .B2(new_n189), .ZN(new_n1054));
  OAI221_X1 g868(.A(new_n1044), .B1(new_n189), .B2(new_n1046), .C1(new_n1052), .C2(new_n1054), .ZN(G72));
  INV_X1    g869(.A(new_n747), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1038), .A2(new_n1021), .A3(new_n1039), .ZN(new_n1057));
  NAND2_X1  g871(.A1(G472), .A2(G902), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n1058), .B(KEYINPUT63), .Z(new_n1059));
  XOR2_X1   g873(.A(new_n1059), .B(KEYINPUT126), .Z(new_n1060));
  AOI21_X1  g874(.A(new_n1056), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g875(.A1(new_n1050), .A2(new_n838), .A3(new_n1031), .A4(new_n1021), .ZN(new_n1062));
  INV_X1    g876(.A(KEYINPUT127), .ZN(new_n1063));
  AND3_X1   g877(.A1(new_n1062), .A2(new_n1063), .A3(new_n1060), .ZN(new_n1064));
  AOI21_X1  g878(.A(new_n1063), .B1(new_n1062), .B2(new_n1060), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n746), .A2(new_n194), .ZN(new_n1066));
  NOR3_X1   g880(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n1056), .A2(new_n1059), .A3(new_n1066), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n957), .B1(new_n947), .B2(new_n1068), .ZN(new_n1069));
  NOR3_X1   g883(.A1(new_n1061), .A2(new_n1067), .A3(new_n1069), .ZN(G57));
endmodule


