//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G232), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G97), .C2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT66), .Z(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n217), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n225), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G20), .ZN(new_n233));
  INV_X1    g0033(.A(new_n201), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n227), .B(new_n230), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n208), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT2), .ZN(new_n240));
  INV_X1    g0040(.A(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  INV_X1    g0044(.A(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n207), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT67), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G50), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(G107), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(KEYINPUT70), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G222), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n260), .B2(new_n265), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n268), .B1(new_n214), .B2(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n273), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n281), .B2(new_n241), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT69), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G190), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT74), .ZN(new_n287));
  INV_X1    g0087(.A(G200), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n286), .B(new_n287), .C1(new_n288), .C2(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  INV_X1    g0090(.A(G20), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n290), .A2(new_n291), .A3(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n202), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n231), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n291), .A2(G1), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n291), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(G150), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G20), .A2(G33), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n301), .A2(new_n302), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(G20), .B2(new_n203), .ZN(new_n307));
  INV_X1    g0107(.A(new_n295), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n293), .B1(new_n202), .B2(new_n300), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT9), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n286), .B(new_n310), .C1(new_n288), .C2(new_n285), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n289), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n284), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(G200), .B2(new_n284), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(new_n310), .C1(new_n287), .C2(KEYINPUT10), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n300), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G77), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT15), .B(G87), .Z(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n302), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n301), .A2(new_n305), .B1(new_n291), .B2(new_n214), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n295), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n292), .A2(new_n214), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n266), .A2(G232), .A3(new_n267), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT72), .B(G107), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n328), .B1(new_n266), .B2(new_n329), .C1(new_n270), .C2(new_n213), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n278), .B1(new_n330), .B2(new_n273), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n281), .A2(new_n215), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n327), .B1(new_n334), .B2(G179), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n278), .B(new_n332), .C1(new_n330), .C2(new_n273), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(G169), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(G200), .ZN(new_n340));
  INV_X1    g0140(.A(new_n327), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT73), .B1(new_n336), .B2(G190), .ZN(new_n342));
  AND4_X1   g0142(.A1(KEYINPUT73), .A2(new_n331), .A3(G190), .A4(new_n333), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n285), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n309), .C1(G169), .C2(new_n285), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n339), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n318), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT84), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT17), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT78), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n261), .ZN(new_n356));
  NAND2_X1  g0156(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(G33), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(new_n291), .A3(new_n263), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT7), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n358), .A2(new_n361), .A3(new_n291), .A4(new_n263), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(G68), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT79), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n360), .A2(KEYINPUT79), .A3(G68), .A4(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(G58), .B(G68), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(G20), .B1(G159), .B2(new_n304), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n371));
  NOR2_X1   g0171(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n262), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n373), .A2(KEYINPUT7), .A3(new_n291), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n260), .A2(new_n265), .A3(new_n291), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n374), .A2(new_n264), .B1(new_n375), .B2(new_n361), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n369), .B1(new_n376), .B2(new_n212), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(new_n295), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT81), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n358), .A2(new_n263), .B1(new_n271), .B2(new_n267), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n241), .A2(G1698), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT82), .B1(new_n385), .B2(new_n280), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n271), .A2(new_n267), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n371), .A2(new_n372), .A3(new_n262), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n384), .B(new_n387), .C1(new_n388), .C2(new_n259), .ZN(new_n389));
  INV_X1    g0189(.A(new_n382), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n280), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n281), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n278), .B1(new_n395), .B2(G232), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n314), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n396), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n288), .B1(new_n398), .B2(new_n391), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n297), .A2(G13), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n301), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n319), .B2(new_n301), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT80), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n380), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(KEYINPUT84), .A2(KEYINPUT17), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n354), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n380), .A2(new_n400), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n353), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT77), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n305), .A2(new_n202), .B1(new_n302), .B2(new_n214), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n291), .A2(G68), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n295), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT11), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n319), .A2(G68), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n292), .A2(new_n212), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT12), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n266), .A2(G226), .A3(new_n267), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n266), .A2(G232), .A3(G1698), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G97), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n273), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n281), .A2(new_n213), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  XOR2_X1   g0226(.A(new_n278), .B(KEYINPUT75), .Z(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT13), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n425), .B1(new_n423), .B2(new_n273), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT13), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n427), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n419), .B1(new_n433), .B2(G200), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n431), .A2(KEYINPUT76), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n435), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n430), .A2(new_n437), .A3(new_n427), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(G190), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n411), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  AND4_X1   g0240(.A1(new_n431), .A2(new_n424), .A3(new_n426), .A4(new_n427), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n431), .B1(new_n430), .B2(new_n427), .ZN(new_n442));
  OAI21_X1  g0242(.A(G200), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n419), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n411), .A2(new_n443), .A3(new_n439), .A4(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n389), .A2(new_n390), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n392), .B1(new_n447), .B2(new_n273), .ZN(new_n448));
  AOI211_X1 g0248(.A(KEYINPUT82), .B(new_n280), .C1(new_n389), .C2(new_n390), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n345), .B(new_n396), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT83), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G169), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n398), .B2(new_n391), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n394), .A2(KEYINPUT83), .A3(new_n345), .A4(new_n396), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n380), .A2(new_n404), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT18), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(G169), .B1(new_n441), .B2(new_n442), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT14), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT14), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n433), .A2(new_n465), .A3(G169), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n436), .A2(G179), .A3(new_n438), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n419), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n410), .A2(new_n446), .A3(new_n462), .A4(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT85), .B1(new_n350), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n410), .A2(new_n462), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n434), .A2(new_n411), .A3(new_n439), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n443), .A2(new_n439), .A3(new_n444), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT77), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n419), .B2(new_n468), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT85), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n473), .A2(new_n478), .A3(new_n349), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n267), .A2(G264), .ZN(new_n482));
  NOR2_X1   g0282(.A1(G257), .A2(G1698), .ZN(new_n483));
  AOI211_X1 g0283(.A(new_n482), .B(new_n483), .C1(new_n358), .C2(new_n263), .ZN(new_n484));
  XOR2_X1   g0284(.A(KEYINPUT88), .B(G303), .Z(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(new_n260), .A3(new_n265), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n273), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n493), .A2(new_n277), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n280), .A2(new_n493), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n245), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n488), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT21), .A3(G169), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n488), .A2(G179), .A3(new_n494), .A4(new_n497), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n502), .B(new_n291), .C1(G33), .C2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(new_n295), .C1(new_n291), .C2(G116), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT20), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n505), .B(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n308), .B(new_n401), .C1(G1), .C2(new_n262), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G116), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n507), .B(new_n510), .C1(G116), .C2(new_n401), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G169), .A3(new_n498), .ZN(new_n512));
  XNOR2_X1  g0312(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n501), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n495), .A2(new_n210), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n358), .A2(new_n263), .B1(new_n221), .B2(new_n267), .ZN(new_n517));
  INV_X1    g0317(.A(G257), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G1698), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n517), .A2(new_n519), .B1(G33), .B2(G294), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n516), .B(new_n494), .C1(new_n520), .C2(new_n280), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n453), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n521), .A2(G179), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n262), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n291), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n291), .A2(KEYINPUT23), .A3(G107), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n329), .A2(G20), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(KEYINPUT23), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT22), .ZN(new_n530));
  AOI21_X1  g0330(.A(G20), .B1(new_n358), .B2(new_n263), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n291), .ZN(new_n533));
  AOI211_X1 g0333(.A(new_n220), .B(new_n533), .C1(new_n260), .C2(new_n265), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n526), .B(new_n529), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n266), .A2(new_n530), .A3(new_n291), .A4(G87), .ZN(new_n537));
  AOI211_X1 g0337(.A(G20), .B(new_n220), .C1(new_n358), .C2(new_n263), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n530), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(new_n526), .A4(new_n529), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n308), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n209), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT25), .B1(new_n292), .B2(new_n209), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n508), .A2(new_n209), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n522), .B(new_n523), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n514), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n488), .A2(new_n494), .A3(new_n497), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n288), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n498), .A2(new_n314), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n549), .A2(new_n550), .A3(new_n511), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n521), .A2(new_n288), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT90), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT90), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n521), .A2(new_n554), .A3(new_n288), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n555), .C1(G190), .C2(new_n521), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n542), .A2(new_n545), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n551), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n304), .A2(G77), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n503), .A2(new_n209), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n560), .B1(new_n563), .B2(KEYINPUT6), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G20), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n559), .B(new_n565), .C1(new_n376), .C2(new_n329), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n295), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n258), .A2(new_n259), .A3(new_n257), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT70), .B1(new_n263), .B2(new_n264), .ZN(new_n569));
  OAI211_X1 g0369(.A(G250), .B(G1698), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n215), .A2(G1698), .ZN(new_n571));
  OAI211_X1 g0371(.A(KEYINPUT4), .B(new_n571), .C1(new_n568), .C2(new_n569), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n571), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n358), .B2(new_n263), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n502), .B1(new_n575), .B2(KEYINPUT4), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n273), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n494), .B1(new_n518), .B2(new_n495), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(G190), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n401), .A2(G97), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n509), .B2(G97), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n567), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT86), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n574), .B1(new_n260), .B2(new_n265), .ZN(new_n585));
  AOI22_X1  g0385(.A1(KEYINPUT4), .A2(new_n585), .B1(new_n269), .B2(G250), .ZN(new_n586));
  INV_X1    g0386(.A(new_n502), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n358), .A2(new_n263), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n571), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n280), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n584), .B1(new_n592), .B2(new_n578), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n577), .A2(KEYINPUT86), .A3(new_n579), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(G200), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n583), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n321), .A2(new_n401), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n508), .A2(new_n220), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n588), .A2(new_n291), .A3(G68), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n291), .B1(new_n422), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n329), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n220), .A2(new_n503), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n291), .A2(G33), .A3(G97), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT87), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n605), .A2(new_n606), .A3(new_n600), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n605), .B2(new_n600), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n599), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  AOI211_X1 g0410(.A(new_n597), .B(new_n598), .C1(new_n610), .C2(new_n295), .ZN(new_n611));
  INV_X1    g0411(.A(new_n490), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n277), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n280), .A2(G250), .A3(new_n612), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n358), .A2(new_n263), .B1(new_n215), .B2(G1698), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n213), .A2(new_n267), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n525), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n614), .B(new_n615), .C1(new_n618), .C2(new_n280), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n215), .A2(G1698), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n588), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n273), .B1(new_n622), .B2(new_n525), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n623), .A2(G190), .A3(new_n614), .A4(new_n615), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n611), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n619), .A2(new_n453), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n623), .A2(new_n345), .A3(new_n614), .A4(new_n615), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n610), .A2(new_n295), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n509), .A2(new_n321), .ZN(new_n629));
  INV_X1    g0429(.A(new_n597), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n592), .A2(new_n578), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n345), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n567), .A2(new_n582), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n577), .A2(new_n579), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n453), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n596), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n481), .A2(new_n547), .A3(new_n558), .A4(new_n640), .ZN(G372));
  INV_X1    g0441(.A(new_n632), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n633), .A3(KEYINPUT26), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n625), .A2(new_n632), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n639), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n642), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n514), .A2(new_n546), .B1(new_n556), .B2(new_n557), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n481), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n347), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n443), .A2(new_n439), .A3(new_n444), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n469), .B1(new_n339), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n410), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n462), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT91), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n318), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n313), .A2(new_n317), .A3(KEYINPUT91), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n653), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n652), .A2(new_n662), .ZN(G369));
  NOR2_X1   g0463(.A1(new_n290), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n275), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n511), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n514), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n514), .A2(new_n671), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n551), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n556), .A2(new_n557), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n670), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n557), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n546), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n546), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n514), .A2(new_n670), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n680), .A2(new_n686), .B1(new_n681), .B2(new_n678), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n228), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G1), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n329), .A2(new_n220), .A3(new_n503), .A4(new_n524), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n692), .A2(new_n693), .B1(new_n235), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT93), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n596), .A2(new_n696), .A3(new_n639), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n596), .B2(new_n639), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n633), .B(new_n649), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n648), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n700), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT29), .B1(new_n651), .B2(new_n678), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n640), .A2(new_n547), .A3(new_n558), .A4(new_n678), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n500), .A2(new_n619), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n520), .A2(new_n280), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n515), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n705), .A2(new_n634), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT92), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT30), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n498), .A2(new_n345), .A3(new_n619), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n521), .A3(new_n637), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n708), .A2(KEYINPUT92), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n670), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n704), .A2(new_n716), .A3(KEYINPUT31), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n718), .A3(new_n670), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n703), .B1(G330), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n695), .B1(new_n721), .B2(G1), .ZN(G364));
  OR2_X1    g0522(.A1(new_n674), .A2(G330), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n275), .B1(new_n664), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n690), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n723), .A2(new_n675), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT94), .Z(new_n729));
  INV_X1    g0529(.A(new_n266), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n689), .A2(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(G355), .B1(new_n524), .B2(new_n689), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  NOR2_X1   g0533(.A1(new_n689), .A2(new_n588), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n234), .A2(new_n489), .A3(G50), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n251), .B2(new_n489), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n733), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n231), .B1(G20), .B2(new_n453), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n727), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n742), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT96), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n291), .A2(new_n314), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(new_n749), .B2(G179), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n748), .A2(KEYINPUT96), .A3(new_n345), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n291), .A2(G190), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(new_n345), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n753), .A2(G50), .B1(G107), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n345), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n747), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n754), .A2(new_n758), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G58), .A2(new_n760), .B1(new_n762), .B2(G77), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n754), .A2(new_n345), .A3(new_n288), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G159), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n763), .B1(KEYINPUT32), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(KEYINPUT32), .B2(new_n766), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n754), .A2(G179), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G68), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n314), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n291), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n266), .B1(new_n503), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n748), .A2(G179), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G87), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n757), .A2(new_n768), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n765), .A2(G329), .ZN(new_n778));
  INV_X1    g0578(.A(new_n775), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G283), .B2(new_n756), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n753), .A2(G326), .ZN(new_n783));
  INV_X1    g0583(.A(new_n773), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G294), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n759), .A2(new_n786), .B1(new_n761), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n266), .B(new_n788), .C1(new_n770), .C2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n782), .A2(new_n783), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n777), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n741), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n744), .B1(new_n745), .B2(new_n792), .C1(new_n674), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n729), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT97), .ZN(G396));
  NAND2_X1  g0596(.A1(new_n651), .A2(new_n678), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n327), .A2(new_n670), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n338), .B1(new_n344), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n339), .A2(new_n670), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n797), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n720), .A2(G330), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n727), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n756), .A2(G87), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n806), .B1(new_n787), .B2(new_n764), .C1(new_n503), .C2(new_n773), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n266), .B(new_n807), .C1(G294), .C2(new_n760), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n775), .A2(G107), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n753), .A2(G303), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT98), .B(G283), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n812), .A2(new_n769), .B1(new_n761), .B2(new_n524), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT99), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G143), .ZN(new_n816));
  INV_X1    g0616(.A(G159), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n759), .A2(new_n816), .B1(new_n761), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(new_n753), .B2(G137), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n303), .B2(new_n769), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  INV_X1    g0621(.A(new_n588), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G50), .B2(new_n775), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n784), .A2(G58), .B1(new_n765), .B2(G132), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n755), .A2(new_n212), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n815), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n742), .A2(new_n739), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n827), .A2(new_n742), .B1(new_n214), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n726), .C1(new_n740), .C2(new_n801), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n805), .A2(new_n830), .ZN(G384));
  NOR2_X1   g0631(.A1(new_n469), .A2(new_n670), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT38), .ZN(new_n833));
  INV_X1    g0633(.A(new_n668), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n457), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n458), .A2(new_n835), .A3(new_n408), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT102), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(new_n668), .B1(new_n380), .B2(new_n404), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n842), .A2(KEYINPUT102), .A3(new_n836), .A4(new_n408), .ZN(new_n843));
  INV_X1    g0643(.A(new_n403), .ZN(new_n844));
  INV_X1    g0644(.A(new_n369), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n365), .B2(new_n366), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT16), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n308), .B1(new_n846), .B2(KEYINPUT16), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n408), .B1(new_n849), .B2(new_n840), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n668), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n839), .A2(new_n843), .B1(new_n852), .B2(KEYINPUT37), .ZN(new_n853));
  INV_X1    g0653(.A(new_n851), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n410), .B2(new_n462), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n833), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n850), .B2(new_n851), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n841), .A2(new_n405), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT102), .B1(new_n858), .B2(new_n836), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n841), .A2(new_n405), .A3(new_n838), .A4(KEYINPUT37), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n472), .A2(new_n851), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n836), .B1(new_n842), .B2(new_n408), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n839), .B2(new_n843), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n835), .B1(new_n410), .B2(new_n462), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n833), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n863), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n832), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n460), .A2(new_n461), .A3(new_n668), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT101), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n444), .A2(new_n678), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n468), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n446), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n876), .A2(KEYINPUT100), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(KEYINPUT100), .ZN(new_n881));
  AOI221_X4 g0681(.A(new_n654), .B1(new_n880), .B2(new_n881), .C1(new_n468), .C2(new_n419), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n875), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n876), .B1(new_n477), .B2(new_n468), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n881), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n469), .A2(new_n475), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT101), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n800), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n797), .B2(new_n799), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n864), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n873), .A2(new_n874), .A3(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT103), .Z(new_n893));
  NAND2_X1  g0693(.A1(new_n481), .A2(new_n703), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n662), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n717), .A2(new_n719), .A3(new_n801), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n883), .B2(new_n887), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n871), .B1(new_n898), .B2(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT40), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(KEYINPUT104), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n902), .B(new_n897), .C1(new_n883), .C2(new_n887), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n856), .A2(new_n863), .A3(new_n901), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n481), .A2(new_n720), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(G330), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n896), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n896), .A2(new_n909), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(KEYINPUT105), .B2(new_n911), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n912), .B1(KEYINPUT105), .B2(new_n911), .C1(new_n275), .C2(new_n664), .ZN(new_n913));
  OAI211_X1 g0713(.A(G20), .B(new_n232), .C1(new_n564), .C2(KEYINPUT35), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n524), .B(new_n914), .C1(KEYINPUT35), .C2(new_n564), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  OAI21_X1  g0716(.A(G77), .B1(new_n207), .B2(new_n212), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n235), .A2(new_n917), .B1(G50), .B2(new_n212), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(G1), .A3(new_n290), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n913), .A2(new_n916), .A3(new_n919), .ZN(G367));
  NOR2_X1   g0720(.A1(new_n697), .A2(new_n698), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n636), .A2(new_n670), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n639), .A2(new_n678), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n685), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n683), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n686), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT42), .B1(new_n930), .B2(new_n926), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n921), .A2(new_n546), .A3(new_n923), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n678), .B1(new_n932), .B2(new_n643), .ZN(new_n933));
  INV_X1    g0733(.A(new_n686), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n683), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT42), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n924), .C2(new_n925), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n931), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n611), .A2(new_n678), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n642), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n646), .B2(new_n940), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT106), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n931), .A2(new_n944), .A3(new_n933), .A4(new_n937), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n939), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n942), .B(KEYINPUT43), .Z(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n939), .B2(new_n945), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT107), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n949), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT107), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n946), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n928), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n953), .A3(new_n928), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n687), .B1(new_n924), .B2(new_n925), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT45), .Z(new_n958));
  NOR3_X1   g0758(.A1(new_n687), .A2(new_n924), .A3(new_n925), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n684), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n960), .A3(new_n685), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n929), .A2(new_n686), .ZN(new_n964));
  OAI211_X1 g0764(.A(G330), .B(new_n674), .C1(new_n964), .C2(new_n935), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n683), .A2(new_n934), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n930), .A2(new_n675), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n962), .A2(new_n721), .A3(new_n963), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n721), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n690), .B(KEYINPUT41), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n955), .B(new_n956), .C1(new_n972), .C2(new_n725), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n588), .B1(G97), .B2(new_n756), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT108), .B(G317), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n765), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(new_n752), .C2(new_n787), .ZN(new_n977));
  INV_X1    g0777(.A(new_n485), .ZN(new_n978));
  INV_X1    g0778(.A(G294), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n978), .A2(new_n759), .B1(new_n979), .B2(new_n769), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n779), .A2(new_n524), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(KEYINPUT46), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(KEYINPUT46), .B2(new_n981), .C1(new_n761), .C2(new_n812), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n977), .B(new_n983), .C1(new_n602), .C2(new_n784), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n266), .B1(new_n202), .B2(new_n761), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G159), .B2(new_n770), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n756), .A2(G77), .B1(new_n765), .B2(G137), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(new_n207), .C2(new_n779), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G143), .B2(new_n753), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n773), .A2(new_n212), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G150), .B2(new_n760), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT109), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n984), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  AOI21_X1  g0794(.A(new_n727), .B1(new_n994), .B2(new_n742), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n743), .B1(new_n228), .B2(new_n322), .C1(new_n735), .C2(new_n246), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n942), .A2(new_n793), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n973), .A2(new_n998), .ZN(G387));
  OR2_X1    g0799(.A1(new_n721), .A2(new_n968), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n721), .A2(new_n968), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n690), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n968), .A2(new_n725), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n242), .A2(new_n489), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1004), .A2(new_n734), .B1(new_n693), .B2(new_n731), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n301), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n202), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n212), .A2(new_n214), .ZN(new_n1009));
  NOR4_X1   g0809(.A1(new_n1008), .A2(G45), .A3(new_n1009), .A4(new_n693), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n1005), .A2(new_n1010), .B1(G107), .B2(new_n228), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n743), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G311), .A2(new_n770), .B1(new_n762), .B2(new_n485), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n752), .B2(new_n786), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n760), .B2(new_n975), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT48), .Z(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n979), .B2(new_n779), .C1(new_n773), .C2(new_n812), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT49), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n765), .A2(G326), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n588), .B1(G116), .B2(new_n756), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n779), .A2(new_n214), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n303), .B2(new_n764), .C1(new_n322), .C2(new_n773), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n588), .B1(new_n503), .B2(new_n755), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n759), .A2(new_n202), .B1(new_n761), .B2(new_n212), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n817), .B2(new_n752), .C1(new_n301), .C2(new_n769), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1023), .A2(new_n1030), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1012), .B1(new_n929), .B2(new_n793), .C1(new_n1031), .C2(new_n745), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1002), .B(new_n1003), .C1(new_n727), .C2(new_n1032), .ZN(G393));
  NAND2_X1  g0833(.A1(new_n962), .A2(new_n963), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n1001), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n690), .A3(new_n969), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n962), .A2(new_n725), .A3(new_n963), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n926), .A2(new_n741), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n588), .B1(new_n202), .B2(new_n769), .C1(new_n301), .C2(new_n761), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n806), .B1(new_n214), .B2(new_n773), .C1(new_n779), .C2(new_n212), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n752), .A2(new_n303), .B1(new_n817), .B2(new_n759), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT51), .Z(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT110), .B(KEYINPUT111), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1039), .B(new_n1040), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n816), .B2(new_n764), .C1(new_n1043), .C2(new_n1042), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n784), .A2(G116), .B1(new_n756), .B2(G107), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n779), .B2(new_n812), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n730), .B1(new_n979), .B2(new_n761), .C1(new_n978), .C2(new_n769), .ZN(new_n1048));
  INV_X1    g0848(.A(G317), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n752), .A2(new_n1049), .B1(new_n787), .B2(new_n759), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT52), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1047), .B(new_n1048), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .C1(new_n786), .C2(new_n764), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1045), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n727), .B1(new_n1054), .B2(new_n742), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n743), .B1(new_n503), .B2(new_n228), .C1(new_n255), .C2(new_n735), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1038), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1036), .A2(new_n1037), .A3(new_n1057), .ZN(G390));
  INV_X1    g0858(.A(KEYINPUT112), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n670), .B(new_n799), .C1(new_n699), .C2(new_n648), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n800), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n799), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n700), .A2(new_n678), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1063), .A2(KEYINPUT112), .A3(new_n889), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n888), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n832), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n871), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT113), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n884), .A2(KEYINPUT101), .A3(new_n886), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT101), .B1(new_n884), .B2(new_n886), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n890), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1066), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1074), .B(new_n865), .C1(KEYINPUT39), .C2(new_n871), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1065), .A2(KEYINPUT113), .A3(new_n871), .A4(new_n1066), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1069), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n717), .A2(new_n801), .A3(G330), .A4(new_n719), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n883), .B2(new_n887), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1078), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n888), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1069), .A2(new_n1075), .A3(new_n1076), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n481), .A2(G330), .A3(new_n720), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1085), .A2(new_n894), .A3(new_n662), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n888), .A2(new_n1081), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n890), .B1(new_n1087), .B2(new_n1079), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1072), .A2(new_n1078), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n1090), .A3(new_n1082), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT114), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1086), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1084), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1093), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1080), .A2(new_n1083), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n690), .A3(new_n1100), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n866), .A2(new_n740), .A3(new_n872), .ZN(new_n1102));
  INV_X1    g0902(.A(G125), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n266), .B1(new_n1103), .B2(new_n764), .C1(new_n817), .C2(new_n773), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  AOI22_X1  g0905(.A1(G137), .A2(new_n770), .B1(new_n762), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(G132), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n759), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1104), .B(new_n1108), .C1(G50), .C2(new_n756), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n775), .A2(G150), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT53), .Z(new_n1111));
  INV_X1    g0911(.A(G128), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1109), .B(new_n1111), .C1(new_n1112), .C2(new_n752), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT116), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n764), .A2(new_n979), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n826), .B(new_n1115), .C1(G77), .C2(new_n784), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n266), .B1(new_n775), .B2(G87), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n602), .A2(new_n770), .B1(new_n762), .B2(G97), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(G283), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1119), .B1(new_n524), .B2(new_n759), .C1(new_n1120), .C2(new_n752), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n745), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n828), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n726), .B1(new_n1006), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT115), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1102), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n725), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1101), .A2(new_n1128), .ZN(G378));
  OAI221_X1 g0929(.A(new_n1025), .B1(new_n207), .B2(new_n755), .C1(new_n1120), .C2(new_n764), .ZN(new_n1130));
  AOI21_X1  g0930(.A(G41), .B1(new_n760), .B2(G107), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n503), .B2(new_n769), .ZN(new_n1132));
  NOR4_X1   g0932(.A1(new_n1130), .A2(new_n588), .A3(new_n990), .A4(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n524), .B2(new_n752), .C1(new_n322), .C2(new_n761), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT58), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n202), .B1(new_n388), .B2(G41), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n773), .A2(new_n303), .ZN(new_n1137));
  INV_X1    g0937(.A(G137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n759), .A2(new_n1112), .B1(new_n761), .B2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1137), .B(new_n1139), .C1(new_n775), .C2(new_n1105), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n1103), .B2(new_n752), .C1(new_n1107), .C2(new_n769), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT59), .Z(new_n1142));
  AOI21_X1  g0942(.A(G41), .B1(new_n765), .B2(G124), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G33), .B1(new_n756), .B2(G159), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1135), .A2(new_n1136), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n727), .B1(new_n1146), .B2(new_n742), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n660), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT91), .B1(new_n313), .B2(new_n317), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n347), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n309), .A2(new_n834), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n661), .A2(new_n347), .A3(new_n1152), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT55), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1148), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT55), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(KEYINPUT56), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1147), .B1(G50), .B2(new_n1123), .C1(new_n1164), .C2(new_n740), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT117), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n899), .A2(KEYINPUT40), .B1(new_n903), .B2(new_n904), .ZN(new_n1167));
  INV_X1    g0967(.A(G330), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT118), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT118), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT104), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1072), .B2(new_n897), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n901), .B1(new_n1172), .B2(new_n871), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n902), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n904), .A2(new_n898), .A3(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1170), .B(G330), .C1(new_n1173), .C2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1169), .A2(new_n1176), .A3(new_n1164), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(new_n1170), .A3(G330), .A4(new_n906), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT119), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n892), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .A4(new_n892), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1166), .B1(new_n1185), .B2(new_n725), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1100), .A2(new_n1086), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n892), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1177), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1190), .A2(new_n1187), .A3(KEYINPUT57), .A4(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n690), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1186), .B1(new_n1188), .B2(new_n1193), .ZN(G375));
  OR2_X1    g0994(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1097), .A2(new_n971), .A3(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT120), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n726), .B1(G68), .B2(new_n1123), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT121), .Z(new_n1199));
  NOR2_X1   g0999(.A1(new_n779), .A2(new_n503), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n730), .B1(new_n214), .B2(new_n755), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n322), .A2(new_n773), .B1(new_n780), .B2(new_n764), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n524), .A2(new_n769), .B1(new_n759), .B2(new_n1120), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n979), .B2(new_n752), .C1(new_n329), .C2(new_n761), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n779), .A2(new_n817), .B1(new_n755), .B2(new_n207), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G50), .B2(new_n784), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n822), .B1(G150), .B2(new_n762), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n1112), .C2(new_n764), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT122), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(KEYINPUT122), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n753), .A2(G132), .B1(new_n770), .B2(new_n1105), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n759), .A2(new_n1138), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1205), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1199), .B1(new_n1215), .B2(new_n742), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT123), .Z(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1072), .B2(new_n739), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1092), .B2(new_n725), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1197), .A2(new_n1219), .ZN(G381));
  INV_X1    g1020(.A(G390), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n973), .A2(new_n998), .A3(new_n1221), .ZN(new_n1222));
  OR3_X1    g1022(.A1(new_n1222), .A2(G396), .A3(G393), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1183), .A2(new_n1184), .B1(new_n1086), .B2(new_n1100), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n690), .B(new_n1192), .C1(new_n1224), .C2(KEYINPUT57), .ZN(new_n1225));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1226), .A3(new_n1186), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n1223), .A2(new_n1227), .A3(G384), .A4(G381), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(G407));
  OAI21_X1  g1029(.A(G213), .B1(new_n1227), .B2(G343), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT124), .ZN(G409));
  INV_X1    g1032(.A(new_n956), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n725), .B1(new_n970), .B2(new_n971), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n954), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n998), .ZN(new_n1236));
  OAI21_X1  g1036(.A(G390), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1222), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT127), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(G396), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1237), .A2(KEYINPUT127), .A3(new_n1222), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G375), .A2(G378), .ZN(new_n1246));
  INV_X1    g1046(.A(G213), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(G343), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1190), .A2(new_n725), .A3(new_n1191), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n971), .B2(new_n1224), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1101), .A2(new_n1128), .A3(new_n1165), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1248), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n691), .B1(new_n1195), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1254), .B(new_n1093), .C1(new_n1253), .C2(new_n1195), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1219), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1246), .A2(new_n1252), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1246), .A2(new_n1252), .A3(KEYINPUT125), .A4(new_n1261), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1248), .A2(G2897), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1261), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G2897), .B(new_n1248), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1226), .B1(new_n1225), .B2(new_n1186), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1185), .A2(new_n971), .A3(new_n1187), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1190), .A2(new_n725), .A3(new_n1191), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1251), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1248), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1270), .B(new_n1271), .C1(new_n1272), .C2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1262), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1268), .B(new_n1278), .C1(new_n1279), .C2(new_n1265), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1245), .B1(new_n1267), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1272), .A2(new_n1277), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT125), .B1(new_n1283), .B2(new_n1261), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1266), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1282), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1278), .A2(new_n1268), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(new_n1245), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1279), .A2(KEYINPUT63), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1281), .A2(new_n1290), .ZN(G405));
  NAND2_X1  g1091(.A1(new_n1246), .A2(new_n1227), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1292), .A2(new_n1261), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1261), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1245), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1295), .B(new_n1296), .ZN(G402));
endmodule


