//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1198, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  OR3_X1    g0009(.A1(new_n209), .A2(KEYINPUT64), .A3(G13), .ZN(new_n210));
  OAI21_X1  g0010(.A(KEYINPUT64), .B1(new_n209), .B2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  AOI211_X1 g0020(.A(new_n218), .B(new_n220), .C1(G50), .C2(G226), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n221), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT65), .Z(new_n236));
  AOI211_X1 g0036(.A(new_n214), .B(new_n231), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n224), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  INV_X1    g0046(.A(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT68), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  OAI21_X1  g0058(.A(G303), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n260), .A2(new_n261), .A3(G257), .A4(new_n262), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n260), .A2(new_n261), .A3(G264), .A4(G1698), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n259), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  OAI211_X1 g0066(.A(G1), .B(G13), .C1(new_n257), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT5), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G41), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n271), .A2(new_n272), .A3(new_n274), .A4(G274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G270), .A3(new_n267), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n269), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G13), .A3(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n280), .A2(new_n232), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT78), .B1(new_n257), .B2(G1), .ZN(new_n283));
  OR3_X1    g0083(.A1(new_n257), .A2(KEYINPUT78), .A3(G1), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n282), .A2(G116), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n280), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(KEYINPUT79), .A3(new_n247), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT79), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n280), .B2(G116), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n281), .A2(new_n232), .B1(G20), .B2(new_n247), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G283), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n292), .B(new_n233), .C1(G33), .C2(new_n205), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n291), .A2(KEYINPUT20), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT20), .B1(new_n291), .B2(new_n293), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n285), .B(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n278), .A2(G169), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT21), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n269), .A2(new_n277), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(G179), .A3(new_n275), .A4(new_n296), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n278), .A2(new_n296), .A3(KEYINPUT21), .A4(G169), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(KEYINPUT80), .A2(G87), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n260), .A2(new_n261), .A3(new_n304), .A4(new_n233), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT22), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT3), .B(G33), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT22), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n233), .A4(new_n304), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n233), .A2(G33), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n233), .B2(G107), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n312), .A2(G116), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT24), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n281), .A2(new_n232), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n310), .A2(KEYINPUT24), .A3(new_n316), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT25), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n280), .B2(G107), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(new_n206), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT81), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT81), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n326), .B(new_n330), .C1(new_n327), .C2(new_n206), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n322), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n276), .A2(G264), .A3(new_n267), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT83), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT83), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n276), .A2(new_n336), .A3(G264), .A4(new_n267), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n260), .A2(new_n261), .A3(G257), .A4(G1698), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n260), .A2(new_n261), .A3(G250), .A4(new_n262), .ZN(new_n339));
  INV_X1    g0139(.A(G294), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT82), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT82), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G294), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n343), .A3(G33), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n335), .A2(new_n337), .B1(new_n268), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n275), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n333), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n347), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n303), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT69), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n279), .A2(G20), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n357), .B2(new_n202), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(KEYINPUT69), .A3(G50), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n282), .A3(new_n359), .ZN(new_n360));
  OR2_X1    g0160(.A1(KEYINPUT8), .A2(G58), .ZN(new_n361));
  NAND2_X1  g0161(.A1(KEYINPUT8), .A2(G58), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G150), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G20), .A2(G33), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n363), .A2(new_n311), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(G20), .B2(new_n203), .ZN(new_n368));
  INV_X1    g0168(.A(new_n320), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n360), .B1(G50), .B2(new_n280), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT9), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G222), .A2(G1698), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n262), .A2(G223), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n307), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n268), .C1(G77), .C2(new_n307), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n279), .B1(G41), .B2(G45), .ZN(new_n377));
  INV_X1    g0177(.A(G274), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G226), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n267), .A2(new_n377), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n376), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G200), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n370), .A2(new_n371), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n372), .A2(new_n383), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT10), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT13), .ZN(new_n389));
  INV_X1    g0189(.A(new_n379), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n380), .A2(new_n262), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n224), .A2(G1698), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n307), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n390), .B1(new_n395), .B2(new_n268), .ZN(new_n396));
  INV_X1    g0196(.A(new_n381), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G238), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n389), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n267), .B1(new_n393), .B2(new_n394), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n381), .A2(new_n227), .ZN(new_n401));
  NOR4_X1   g0201(.A1(new_n400), .A2(new_n401), .A3(new_n390), .A4(KEYINPUT13), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT14), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n391), .A2(new_n392), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n307), .B1(G33), .B2(G97), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n379), .B1(new_n406), .B2(new_n267), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT13), .B1(new_n407), .B2(new_n401), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n396), .A2(new_n389), .A3(new_n398), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(G169), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n409), .A3(G179), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n404), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n286), .A2(new_n226), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n282), .A2(G68), .A3(new_n356), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n366), .A2(new_n202), .B1(new_n233), .B2(G68), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n311), .A2(new_n216), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n320), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n420), .A2(KEYINPUT11), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(KEYINPUT11), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n416), .B(new_n417), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n410), .B2(G200), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n385), .B2(new_n410), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n382), .A2(new_n348), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n370), .B(new_n428), .C1(G179), .C2(new_n382), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n286), .A2(new_n216), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n282), .A2(G77), .A3(new_n356), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT71), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT71), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n282), .A2(new_n433), .A3(G77), .A4(new_n356), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G20), .A2(G77), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n436), .B1(new_n437), .B2(new_n311), .C1(new_n366), .C2(new_n363), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT70), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n438), .A2(new_n439), .A3(new_n320), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n438), .B2(new_n320), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n430), .B(new_n435), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G200), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n307), .A2(G232), .A3(new_n262), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n307), .A2(G238), .A3(G1698), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n446), .C1(new_n206), .C2(new_n307), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n390), .B1(new_n447), .B2(new_n268), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n397), .A2(G244), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n443), .A2(KEYINPUT72), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(G190), .A3(new_n449), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT72), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n442), .B2(new_n450), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n388), .A2(new_n427), .A3(new_n429), .A4(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(G223), .A2(G1698), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n380), .A2(G1698), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n307), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G87), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n267), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n267), .A2(G232), .A3(new_n377), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n379), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT75), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n379), .A3(KEYINPUT75), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n463), .A2(new_n467), .A3(new_n385), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT76), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n464), .A2(KEYINPUT75), .A3(new_n379), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT75), .B1(new_n464), .B2(new_n379), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT76), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(new_n385), .A4(new_n463), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n444), .B1(new_n462), .B2(new_n465), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n470), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n363), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n356), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n479), .A2(new_n320), .B1(new_n280), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n223), .A2(new_n226), .ZN(new_n481));
  OAI21_X1  g0281(.A(G20), .B1(new_n481), .B2(new_n201), .ZN(new_n482));
  INV_X1    g0282(.A(G159), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(new_n366), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT7), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n307), .B2(G20), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n260), .A2(new_n261), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT7), .A3(new_n233), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n484), .B1(new_n489), .B2(G68), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n369), .B1(new_n490), .B2(KEYINPUT16), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n260), .A2(KEYINPUT74), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT74), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n257), .A3(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n261), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(KEYINPUT7), .A3(new_n233), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n226), .B1(new_n498), .B2(new_n486), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n493), .B1(new_n499), .B2(new_n484), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n480), .B1(new_n491), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n477), .A2(new_n501), .A3(KEYINPUT17), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT17), .B1(new_n477), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n491), .A2(new_n500), .ZN(new_n505));
  INV_X1    g0305(.A(new_n480), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n473), .A2(new_n352), .A3(new_n463), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n348), .B1(new_n462), .B2(new_n465), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(KEYINPUT18), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT18), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n501), .B2(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n504), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n448), .A2(new_n449), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n348), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n448), .A2(new_n352), .A3(new_n449), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n442), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n457), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n276), .A2(new_n267), .ZN(new_n523));
  INV_X1    g0323(.A(G257), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n275), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n260), .A2(new_n261), .A3(G244), .A4(new_n262), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n307), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n307), .A2(G250), .A3(G1698), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n292), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n525), .B1(new_n531), .B2(new_n268), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G179), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n348), .B2(new_n532), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n206), .B1(new_n498), .B2(new_n486), .ZN(new_n535));
  NAND2_X1  g0335(.A1(KEYINPUT6), .A2(G97), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT77), .B1(new_n536), .B2(G107), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT77), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(new_n206), .A3(KEYINPUT6), .A4(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT6), .B1(new_n207), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n543), .A2(new_n233), .B1(new_n216), .B2(new_n366), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n320), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  MUX2_X1   g0345(.A(new_n280), .B(new_n327), .S(G97), .Z(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n534), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n346), .A2(new_n385), .A3(new_n275), .ZN(new_n549));
  AOI21_X1  g0349(.A(G200), .B1(new_n346), .B2(new_n275), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n332), .B(new_n322), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n227), .A2(new_n262), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n217), .A2(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n260), .A2(new_n552), .A3(new_n261), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n267), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n279), .A2(G45), .ZN(new_n557));
  AND2_X1   g0357(.A1(G33), .A2(G41), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(G250), .C1(new_n558), .C2(new_n232), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n557), .A2(new_n378), .ZN(new_n561));
  NOR4_X1   g0361(.A1(new_n556), .A2(new_n385), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n554), .A2(new_n555), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n268), .ZN(new_n564));
  INV_X1    g0364(.A(new_n561), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(new_n559), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(G200), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G87), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n327), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n233), .B1(new_n394), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n205), .A3(new_n206), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n233), .A2(G33), .A3(G97), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n571), .A2(new_n572), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n260), .A2(new_n261), .A3(new_n233), .A4(G68), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n369), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n437), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n280), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n569), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n571), .A2(new_n572), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n573), .A2(new_n570), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n578), .B1(new_n582), .B2(new_n320), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n282), .A2(new_n577), .A3(new_n283), .A4(new_n284), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n566), .A2(new_n348), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n556), .A2(new_n561), .A3(new_n560), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n352), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n567), .A2(new_n579), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AOI211_X1 g0388(.A(G190), .B(new_n525), .C1(new_n268), .C2(new_n531), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n531), .A2(new_n268), .ZN(new_n590));
  INV_X1    g0390(.A(new_n525), .ZN(new_n591));
  AOI21_X1  g0391(.A(G200), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n545), .B(new_n546), .C1(new_n589), .C2(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n548), .A2(new_n551), .A3(new_n588), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n300), .A2(G190), .A3(new_n275), .ZN(new_n595));
  INV_X1    g0395(.A(new_n296), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n278), .A2(G200), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n354), .A2(new_n522), .A3(new_n594), .A4(new_n598), .ZN(G372));
  NAND2_X1  g0399(.A1(new_n426), .A2(new_n521), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(new_n424), .A3(KEYINPUT86), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT86), .B1(new_n600), .B2(new_n424), .ZN(new_n603));
  INV_X1    g0403(.A(new_n504), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n515), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT87), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n603), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n504), .A3(new_n601), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n515), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n388), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n532), .A2(G179), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n532), .A2(new_n348), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT84), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n533), .B(new_n617), .C1(new_n348), .C2(new_n532), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n547), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n588), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n613), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  INV_X1    g0422(.A(new_n562), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n579), .B(new_n623), .C1(new_n444), .C2(new_n586), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n585), .A2(new_n587), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n534), .A2(new_n624), .A3(new_n625), .A4(new_n547), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n626), .B2(new_n613), .ZN(new_n627));
  INV_X1    g0427(.A(new_n548), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(KEYINPUT85), .A3(KEYINPUT26), .A4(new_n588), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n625), .ZN(new_n631));
  INV_X1    g0431(.A(new_n303), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n353), .A2(new_n333), .A3(new_n349), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n594), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n522), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n612), .A2(new_n429), .A3(new_n637), .ZN(G369));
  INV_X1    g0438(.A(G13), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n279), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n333), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n350), .A2(new_n353), .B1(new_n647), .B2(new_n551), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n633), .A2(new_n646), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n632), .A2(new_n646), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n632), .A2(new_n296), .A3(new_n646), .ZN(new_n653));
  INV_X1    g0453(.A(new_n646), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n303), .B1(new_n596), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n598), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G330), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n649), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n650), .A2(new_n651), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n212), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n279), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n572), .A2(G116), .ZN(new_n666));
  INV_X1    g0466(.A(new_n235), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n665), .A2(new_n666), .B1(new_n667), .B2(new_n664), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT28), .Z(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n671));
  INV_X1    g0471(.A(new_n619), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n588), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n673), .B2(KEYINPUT26), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n635), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n670), .B1(new_n675), .B2(new_n654), .ZN(new_n676));
  AOI211_X1 g0476(.A(KEYINPUT29), .B(new_n646), .C1(new_n630), .C2(new_n635), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n594), .A2(new_n354), .A3(new_n598), .A4(new_n654), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n278), .A2(new_n352), .A3(new_n566), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT88), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n532), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n278), .A2(KEYINPUT88), .A3(new_n352), .A4(new_n566), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n682), .A2(new_n347), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n300), .A2(new_n586), .A3(G179), .A4(new_n275), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n532), .A2(new_n346), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n688), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n278), .A2(new_n566), .A3(new_n352), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(KEYINPUT30), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n685), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n646), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n679), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT89), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n684), .A2(new_n683), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n561), .B1(new_n563), .B2(new_n268), .ZN(new_n700));
  AOI21_X1  g0500(.A(G179), .B1(new_n700), .B2(new_n559), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT88), .B1(new_n701), .B2(new_n278), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n699), .A2(new_n351), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT30), .B1(new_n690), .B2(new_n691), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n698), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n685), .A2(KEYINPUT89), .A3(new_n689), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n692), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n657), .B1(new_n697), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n678), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n669), .B1(new_n710), .B2(G1), .ZN(G364));
  INV_X1    g0511(.A(new_n658), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n656), .A2(new_n657), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n640), .A2(G45), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n665), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(KEYINPUT90), .A2(G169), .ZN(new_n717));
  NOR2_X1   g0517(.A1(KEYINPUT90), .A2(G169), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n717), .A2(new_n718), .A3(new_n233), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n232), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT91), .Z(new_n725));
  NOR2_X1   g0525(.A1(new_n236), .A2(G45), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n253), .B2(G45), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n212), .B1(new_n727), .B2(new_n307), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(G355), .B2(new_n307), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n725), .B(new_n729), .C1(G116), .C2(new_n663), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n233), .A2(new_n352), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT92), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G190), .A2(G200), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT92), .B1(new_n233), .B2(new_n352), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n385), .A2(G200), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n738), .A3(new_n736), .ZN(new_n739));
  INV_X1    g0539(.A(G322), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n731), .A2(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n233), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n735), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n307), .B(new_n741), .C1(G329), .C2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n385), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G283), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n732), .A2(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(G317), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT33), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n751), .A2(KEYINPUT33), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n749), .A2(new_n385), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G326), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n738), .A2(new_n352), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n341), .A2(new_n343), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n756), .A2(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(G303), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n745), .A2(new_n748), .A3(new_n754), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n759), .A2(G97), .ZN(new_n767));
  INV_X1    g0567(.A(new_n750), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n767), .B1(new_n768), .B2(new_n226), .C1(new_n202), .C2(new_n756), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n307), .B1(new_n746), .B2(new_n206), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(G87), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n771), .B1(new_n739), .B2(new_n223), .C1(new_n216), .C2(new_n737), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n744), .A2(G159), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT93), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT32), .Z(new_n776));
  OAI21_X1  g0576(.A(new_n766), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n730), .B1(new_n777), .B2(new_n720), .ZN(new_n778));
  INV_X1    g0578(.A(new_n715), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n656), .A2(new_n723), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n716), .A2(new_n781), .ZN(G396));
  AOI21_X1  g0582(.A(new_n646), .B1(new_n630), .B2(new_n635), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT96), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n520), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n518), .A2(new_n442), .A3(KEYINPUT96), .A4(new_n519), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(new_n456), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n442), .A2(new_n646), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n787), .A2(new_n456), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n521), .A2(new_n646), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n789), .B1(new_n783), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(new_n709), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n709), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(new_n798), .A3(new_n715), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n746), .A2(new_n568), .B1(new_n743), .B2(new_n731), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT94), .ZN(new_n801));
  INV_X1    g0601(.A(new_n737), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(G116), .B1(G283), .B2(new_n750), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n206), .B2(new_n763), .ZN(new_n804));
  INV_X1    g0604(.A(new_n739), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n801), .B(new_n804), .C1(G294), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n755), .A2(G303), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n806), .A2(new_n487), .A3(new_n767), .A4(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G137), .A2(new_n755), .B1(new_n750), .B2(G150), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT95), .ZN(new_n810));
  INV_X1    g0610(.A(G143), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n811), .B2(new_n739), .C1(new_n483), .C2(new_n737), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n813), .B1(new_n223), .B2(new_n760), .C1(new_n226), .C2(new_n746), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n307), .B1(new_n743), .B2(new_n815), .C1(new_n202), .C2(new_n763), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n808), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n720), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n793), .A2(new_n721), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n720), .A2(new_n721), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n216), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n818), .A2(new_n779), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n799), .A2(new_n822), .ZN(G384));
  NAND2_X1  g0623(.A1(new_n507), .A2(new_n511), .ZN(new_n824));
  INV_X1    g0624(.A(new_n644), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n507), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n477), .A2(new_n501), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n824), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n829), .A2(KEYINPUT98), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(KEYINPUT98), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n490), .A2(new_n492), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n480), .B1(new_n832), .B2(new_n491), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n511), .B2(new_n825), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(new_n828), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n830), .A2(new_n831), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n516), .A2(new_n825), .A3(new_n834), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n837), .A2(KEYINPUT38), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n477), .A2(new_n501), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n501), .A2(new_n510), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT98), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n827), .A4(new_n826), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n829), .A2(KEYINPUT98), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n843), .A2(new_n826), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n845), .A2(new_n846), .B1(new_n847), .B2(KEYINPUT37), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n826), .B1(new_n504), .B2(new_n515), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n839), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n423), .A2(new_n646), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n424), .A2(new_n426), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n414), .A2(new_n423), .A3(new_n646), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n853), .A2(new_n854), .B1(new_n791), .B2(new_n792), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n679), .A2(new_n696), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(KEYINPUT40), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n851), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n858), .B1(new_n839), .B2(new_n850), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT38), .B1(new_n837), .B2(new_n838), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n827), .B1(new_n835), .B2(new_n828), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n845), .B2(new_n846), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n644), .B(new_n833), .C1(new_n504), .C2(new_n515), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n868), .A2(new_n869), .A3(new_n840), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n857), .B(new_n855), .C1(new_n866), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT40), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT101), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n522), .A2(new_n857), .ZN(new_n876));
  OAI21_X1  g0676(.A(G330), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT102), .Z(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n876), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n787), .A2(new_n646), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n783), .B2(new_n788), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n853), .A2(new_n854), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n840), .B1(new_n868), .B2(new_n869), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n839), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n515), .B2(new_n825), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n414), .A2(new_n423), .A3(new_n654), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT39), .B1(new_n866), .B2(new_n870), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n839), .A2(new_n850), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n880), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n878), .A2(new_n895), .A3(new_n879), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n522), .B1(new_n676), .B2(new_n677), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n612), .A2(new_n900), .A3(new_n429), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT99), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n904), .B(new_n905), .C1(new_n279), .C2(new_n640), .ZN(new_n906));
  INV_X1    g0706(.A(new_n543), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n247), .B1(new_n907), .B2(KEYINPUT35), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n908), .B(new_n234), .C1(KEYINPUT35), .C2(new_n907), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT36), .ZN(new_n910));
  OAI21_X1  g0710(.A(G77), .B1(new_n223), .B2(new_n226), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n911), .A2(new_n235), .B1(G50), .B2(new_n226), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(G1), .A3(new_n639), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT97), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n906), .A2(new_n910), .A3(new_n914), .ZN(G367));
  NOR2_X1   g0715(.A1(new_n663), .A2(new_n307), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n725), .B1(new_n244), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n663), .A2(new_n577), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n715), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n723), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n579), .A2(new_n654), .ZN(new_n921));
  MUX2_X1   g0721(.A(new_n588), .B(new_n631), .S(new_n921), .Z(new_n922));
  OAI21_X1  g0722(.A(new_n307), .B1(new_n746), .B2(new_n216), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT106), .Z(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(G58), .B2(new_n764), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n744), .A2(G137), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G143), .A2(new_n755), .B1(new_n750), .B2(G159), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n202), .A2(new_n737), .B1(new_n739), .B2(new_n364), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n760), .A2(new_n226), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n764), .A2(G116), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT46), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT104), .Z(new_n935));
  OAI221_X1 g0735(.A(new_n935), .B1(new_n933), .B2(new_n932), .C1(new_n761), .C2(new_n768), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT105), .Z(new_n937));
  NOR2_X1   g0737(.A1(new_n746), .A2(new_n205), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n802), .A2(G283), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n805), .A2(G303), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n743), .A2(new_n751), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n307), .B(new_n942), .C1(G107), .C2(new_n759), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n756), .A2(new_n731), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n931), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  INV_X1    g0747(.A(new_n720), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n919), .B1(new_n920), .B2(new_n922), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n714), .A2(G1), .ZN(new_n950));
  INV_X1    g0750(.A(new_n710), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n652), .A2(new_n658), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(new_n661), .A3(new_n659), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n661), .A2(new_n660), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n548), .A2(new_n593), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n547), .A2(new_n646), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n672), .A2(new_n646), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT44), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n955), .A2(new_n958), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n954), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n710), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n664), .B(KEYINPUT41), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n950), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n650), .A2(new_n956), .A3(new_n651), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT42), .Z(new_n969));
  OAI21_X1  g0769(.A(new_n548), .B1(new_n958), .B2(new_n633), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n654), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n974), .B1(new_n972), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n659), .A2(new_n958), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n949), .B1(new_n967), .B2(new_n980), .ZN(G387));
  NAND4_X1  g0781(.A1(new_n952), .A2(new_n661), .A3(new_n659), .A4(new_n950), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G303), .A2(new_n802), .B1(new_n805), .B2(G317), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n731), .B2(new_n768), .C1(new_n740), .C2(new_n756), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT48), .ZN(new_n985));
  INV_X1    g0785(.A(G283), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n985), .B1(new_n986), .B2(new_n760), .C1(new_n761), .C2(new_n763), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT49), .Z(new_n988));
  OAI22_X1  g0788(.A1(new_n746), .A2(new_n247), .B1(new_n743), .B2(new_n757), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n988), .A2(new_n307), .A3(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n802), .A2(G68), .B1(new_n478), .B2(new_n750), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n202), .B2(new_n739), .C1(new_n483), .C2(new_n756), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n760), .A2(new_n437), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n216), .B2(new_n763), .C1(new_n364), .C2(new_n743), .ZN(new_n995));
  NOR4_X1   g0795(.A1(new_n992), .A2(new_n995), .A3(new_n487), .A4(new_n938), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n720), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n723), .B1(new_n648), .B2(new_n649), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n725), .B1(G107), .B2(new_n663), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n241), .A2(new_n270), .A3(new_n307), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n363), .A2(G50), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n270), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT50), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n1001), .A2(new_n1004), .B1(new_n226), .B2(new_n216), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n487), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1000), .B1(new_n666), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n999), .B1(new_n1007), .B2(new_n663), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n997), .A2(new_n779), .A3(new_n998), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n953), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n664), .B1(new_n710), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n982), .B(new_n1009), .C1(new_n954), .C2(new_n1011), .ZN(G393));
  XNOR2_X1  g0812(.A(new_n963), .B(new_n659), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n664), .B(new_n964), .C1(new_n1013), .C2(new_n954), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n950), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n756), .A2(new_n751), .B1(new_n731), .B2(new_n739), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT52), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n746), .A2(new_n206), .B1(new_n743), .B2(new_n740), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n307), .B(new_n1018), .C1(G283), .C2(new_n764), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n247), .B2(new_n760), .C1(new_n340), .C2(new_n737), .ZN(new_n1021));
  INV_X1    g0821(.A(G303), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n768), .A2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n746), .A2(new_n568), .B1(new_n743), .B2(new_n811), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G77), .B2(new_n759), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n226), .B2(new_n763), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n756), .A2(new_n364), .B1(new_n483), .B2(new_n739), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT51), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n487), .B1(new_n750), .B2(G50), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n363), .C2(new_n737), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1021), .A2(new_n1023), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT107), .Z(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n720), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n715), .B1(new_n958), .B2(new_n723), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n725), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n916), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1035), .B1(new_n205), .B2(new_n212), .C1(new_n250), .C2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1014), .A2(new_n1015), .A3(new_n1038), .ZN(G390));
  NAND3_X1  g0839(.A1(new_n855), .A2(G330), .A3(new_n857), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT109), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n855), .A2(new_n857), .A3(KEYINPUT109), .A4(G330), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n890), .B1(new_n882), .B2(new_n884), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n891), .A2(new_n1046), .A3(new_n893), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n890), .B(KEYINPUT108), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n646), .B1(new_n674), .B2(new_n635), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n881), .B1(new_n1049), .B2(new_n788), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n851), .B(new_n1048), .C1(new_n1050), .C2(new_n884), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1045), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT110), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n679), .A2(new_n696), .ZN(new_n1056));
  OAI211_X1 g0856(.A(G330), .B(new_n855), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT111), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n697), .A2(new_n708), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT111), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1059), .A2(new_n1060), .A3(G330), .A4(new_n855), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1047), .A2(new_n1051), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT110), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1054), .B1(new_n1064), .B2(new_n1052), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n857), .A2(KEYINPUT112), .A3(G330), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n794), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT112), .B1(new_n857), .B2(G330), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n884), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1062), .A2(new_n1050), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n882), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n883), .B1(new_n709), .B2(new_n794), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1071), .B1(new_n1044), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n522), .A2(G330), .A3(new_n857), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n612), .A2(new_n900), .A3(new_n429), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1065), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1065), .A2(new_n1079), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n664), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n891), .A2(new_n721), .A3(new_n893), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n771), .B1(new_n340), .B2(new_n743), .C1(new_n756), .C2(new_n986), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n805), .A2(G116), .B1(G77), .B2(new_n759), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT114), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(G107), .C2(new_n750), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n307), .B1(new_n747), .B2(G68), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n205), .C2(new_n737), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT115), .Z(new_n1090));
  AOI22_X1  g0890(.A1(new_n805), .A2(G132), .B1(G50), .B2(new_n747), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1091), .B(new_n307), .C1(new_n483), .C2(new_n760), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G128), .B2(new_n755), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n750), .A2(G137), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n744), .A2(G125), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT54), .B(G143), .Z(new_n1096));
  NAND2_X1  g0896(.A1(new_n802), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n763), .A2(new_n364), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1090), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(new_n720), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n715), .B(new_n1103), .C1(new_n363), .C2(new_n820), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1065), .A2(new_n950), .B1(new_n1083), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1082), .A2(new_n1105), .ZN(G378));
  INV_X1    g0906(.A(KEYINPUT57), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1076), .A2(KEYINPUT119), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1076), .A2(KEYINPUT119), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n1065), .C2(new_n1079), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n862), .A2(new_n863), .ZN(new_n1112));
  AOI211_X1 g0912(.A(KEYINPUT100), .B(new_n858), .C1(new_n839), .C2(new_n850), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n873), .B(G330), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n388), .A2(new_n429), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n370), .A2(new_n825), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n865), .A2(G330), .A3(new_n873), .A4(new_n1119), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n895), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n895), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1107), .B1(new_n1111), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1110), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1081), .A2(new_n1108), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n896), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1121), .A2(new_n1122), .A3(new_n895), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(KEYINPUT57), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1126), .A2(new_n664), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1120), .A2(new_n721), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n756), .A2(new_n247), .B1(new_n437), .B2(new_n737), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n929), .B(new_n1136), .C1(G97), .C2(new_n750), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n206), .B2(new_n739), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n266), .B(new_n487), .C1(new_n763), .C2(new_n216), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n743), .A2(new_n986), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n746), .A2(new_n223), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n266), .B1(new_n255), .B2(new_n257), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1142), .A2(KEYINPUT58), .B1(new_n202), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n755), .A2(G125), .B1(new_n759), .B2(G150), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT117), .Z(new_n1146));
  INV_X1    g0946(.A(new_n1096), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(new_n763), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1148), .A2(KEYINPUT116), .B1(new_n750), .B2(G132), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1146), .B(new_n1149), .C1(KEYINPUT116), .C2(new_n1148), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G137), .B2(new_n802), .ZN(new_n1151));
  INV_X1    g0951(.A(G128), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n739), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT59), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G33), .B1(new_n744), .B2(G124), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n266), .C1(new_n483), .C2(new_n746), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT118), .Z(new_n1157));
  OAI221_X1 g0957(.A(new_n1144), .B1(KEYINPUT58), .B2(new_n1142), .C1(new_n1154), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n720), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n820), .A2(new_n202), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1135), .A2(new_n779), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1132), .B2(new_n950), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1134), .A2(new_n1163), .ZN(G375));
  NAND3_X1  g0964(.A1(new_n1070), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n966), .B(KEYINPUT120), .Z(new_n1166));
  NAND3_X1  g0966(.A1(new_n1078), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n820), .A2(new_n226), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n802), .A2(G107), .B1(G77), .B2(new_n747), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n205), .B2(new_n763), .C1(new_n986), .C2(new_n739), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n994), .B1(new_n247), .B2(new_n768), .C1(new_n1022), .C2(new_n743), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n756), .A2(new_n340), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n307), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n487), .B1(new_n805), .B2(G137), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n815), .B2(new_n756), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1141), .B1(new_n802), .B2(G150), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n483), .B2(new_n763), .C1(new_n768), .C2(new_n1147), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G128), .C2(new_n744), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n759), .A2(G50), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1173), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT121), .Z(new_n1181));
  OAI211_X1 g0981(.A(new_n779), .B(new_n1168), .C1(new_n1181), .C2(new_n948), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n721), .B2(new_n884), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1074), .B2(new_n950), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1167), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT122), .ZN(G381));
  OR2_X1    g0986(.A1(G387), .A2(G390), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1187), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1188));
  INV_X1    g0988(.A(G384), .ZN(new_n1189));
  INV_X1    g0989(.A(G378), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n950), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1161), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n664), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n1194), .B2(new_n1107), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1192), .B1(new_n1195), .B2(new_n1133), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1196), .ZN(G407));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1190), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G407), .B(G213), .C1(G343), .C2(new_n1198), .ZN(G409));
  XNOR2_X1  g0999(.A(G393), .B(G396), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(G387), .A2(G390), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1187), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1200), .B1(new_n1187), .B2(new_n1201), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1190), .B1(new_n1134), .B2(new_n1163), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1128), .A2(new_n1132), .A3(new_n1166), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1163), .ZN(new_n1207));
  INV_X1    g1007(.A(G213), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1207), .A2(G378), .B1(new_n1208), .B2(G343), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n857), .A2(G330), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT112), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(new_n794), .A3(new_n1066), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n884), .A2(new_n1213), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n657), .B(new_n793), .C1(new_n697), .C2(new_n708), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1042), .B(new_n1043), .C1(new_n1215), .C2(new_n883), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1214), .A2(new_n1050), .B1(new_n1071), .B2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1217), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n1076), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT60), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1193), .B1(new_n1165), .B2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1070), .A2(new_n1076), .A3(new_n1073), .A4(KEYINPUT60), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT123), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1218), .A2(new_n1220), .A3(new_n1078), .A4(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1224), .A2(G384), .A3(new_n1184), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G384), .B1(new_n1224), .B2(new_n1184), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT124), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1165), .A2(new_n1219), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n664), .A3(new_n1078), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1184), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1189), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1224), .A2(G384), .A3(new_n1184), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT124), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1228), .A2(new_n1235), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1205), .A2(new_n1209), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT62), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1204), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1208), .A2(G343), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(G2897), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT126), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1241), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1241), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1227), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1233), .A2(KEYINPUT124), .A3(new_n1234), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT126), .B1(new_n1250), .B2(new_n1244), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1246), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G375), .A2(G378), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1110), .B1(new_n1065), .B2(new_n1079), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1254), .A2(new_n1108), .B1(new_n1131), .B2(new_n1130), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1192), .B1(new_n1255), .B2(new_n1166), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1240), .B1(new_n1256), .B2(new_n1190), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1252), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1257), .B(new_n1260), .C1(new_n1196), .C2(new_n1190), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1261), .B2(KEYINPUT62), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1239), .A2(new_n1259), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1253), .A2(new_n1264), .A3(new_n1257), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT125), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT127), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1246), .A2(new_n1251), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1261), .A2(KEYINPUT63), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1253), .A2(new_n1273), .A3(new_n1257), .A4(new_n1260), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1263), .B1(new_n1276), .B2(new_n1204), .ZN(G405));
  AOI22_X1  g1077(.A1(new_n1198), .A2(new_n1253), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1198), .A2(new_n1253), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1260), .B2(new_n1279), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(new_n1204), .ZN(G402));
endmodule


