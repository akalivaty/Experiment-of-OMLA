//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n206), .A2(new_n207), .B1(G155gat), .B2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G141gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n208), .A2(new_n209), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n207), .ZN(new_n220));
  NOR3_X1   g019(.A1(KEYINPUT73), .A2(G155gat), .A3(G162gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n215), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT74), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n212), .A2(KEYINPUT77), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(G141gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n211), .A2(KEYINPUT76), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(new_n210), .B2(G148gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n227), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n204), .A2(new_n205), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n215), .B1(new_n232), .B2(KEYINPUT2), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n219), .A2(new_n223), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT29), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G197gat), .B(G204gat), .ZN(new_n237));
  AND2_X1   g036(.A1(G211gat), .A2(G218gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(KEYINPUT22), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G211gat), .A2(G218gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n239), .B(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n236), .A2(new_n242), .B1(new_n244), .B2(new_n234), .ZN(new_n245));
  NAND2_X1  g044(.A1(G228gat), .A2(G233gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT84), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n249), .A2(G22gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(G22gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n247), .A2(new_n248), .ZN(new_n253));
  XNOR2_X1  g052(.A(G78gat), .B(G106gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT31), .B(G50gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n250), .B(new_n251), .C1(new_n256), .C2(new_n253), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT85), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT23), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(G169gat), .B2(G176gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  MUX2_X1   g068(.A(KEYINPUT24), .B(new_n268), .S(new_n269), .Z(new_n270));
  NAND2_X1  g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT25), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(KEYINPUT23), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n267), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT64), .B(G169gat), .ZN(new_n276));
  INV_X1    g075(.A(G176gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT23), .A3(new_n277), .ZN(new_n278));
  AND4_X1   g077(.A1(new_n267), .A2(new_n270), .A3(new_n271), .A4(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n275), .B1(new_n279), .B2(KEYINPUT25), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT27), .B(G183gat), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n283), .B(KEYINPUT28), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n273), .B(KEYINPUT26), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n271), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n269), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n243), .ZN(new_n289));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(G226gat), .A3(G233gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n293), .A2(new_n242), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n242), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G8gat), .B(G36gat), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT71), .ZN(new_n298));
  XOR2_X1   g097(.A(G64gat), .B(G92gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n263), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n293), .A2(new_n242), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n293), .A2(new_n242), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n300), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT72), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT70), .B1(new_n303), .B2(new_n304), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n300), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n305), .A2(KEYINPUT30), .A3(new_n306), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n308), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n315));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT0), .ZN(new_n317));
  XNOR2_X1  g116(.A(G57gat), .B(G85gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n209), .B(new_n215), .C1(new_n220), .C2(new_n221), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n218), .A2(new_n214), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n223), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G127gat), .B(G134gat), .Z(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT1), .ZN(new_n325));
  INV_X1    g124(.A(G120gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT66), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G120gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n327), .A2(new_n329), .A3(new_n330), .A4(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT66), .B(G120gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n330), .B1(new_n335), .B2(G113gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n325), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n231), .A2(new_n233), .ZN(new_n338));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n324), .B1(KEYINPUT1), .B2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n323), .A2(new_n337), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT79), .B1(new_n341), .B2(KEYINPUT4), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n337), .A2(new_n340), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .A4(new_n234), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n337), .A2(new_n340), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n321), .A2(new_n322), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n208), .A2(new_n209), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n338), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT4), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n348), .B1(new_n234), .B2(new_n235), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n323), .A2(new_n235), .A3(new_n338), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT5), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n353), .A2(new_n354), .A3(new_n359), .A4(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n351), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n341), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n366), .B2(new_n361), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n352), .A2(KEYINPUT78), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n341), .A2(new_n370), .A3(KEYINPUT4), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n360), .B1(new_n355), .B2(new_n357), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n358), .B1(new_n347), .B2(new_n352), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n354), .B1(new_n376), .B2(new_n362), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n320), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n359), .A3(new_n362), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT80), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n380), .A2(new_n319), .A3(new_n363), .A4(new_n374), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n381), .A2(KEYINPUT81), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT81), .B1(new_n381), .B2(new_n382), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n315), .B(new_n378), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n378), .A2(new_n382), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n375), .A2(new_n320), .A3(new_n377), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(KEYINPUT6), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n381), .A2(KEYINPUT81), .A3(new_n382), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n315), .B1(new_n392), .B2(new_n378), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n314), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT83), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n314), .B(new_n396), .C1(new_n387), .C2(new_n393), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n262), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n288), .B(new_n348), .ZN(new_n399));
  AND2_X1   g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n401), .A2(KEYINPUT32), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT69), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  XNOR2_X1  g204(.A(G15gat), .B(G43gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n404), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n399), .A2(new_n400), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n412), .B(KEYINPUT34), .Z(new_n413));
  OAI21_X1  g212(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n411), .B2(new_n414), .ZN(new_n416));
  OR3_X1    g215(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT36), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT36), .B1(new_n415), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n202), .B1(new_n398), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n260), .B(KEYINPUT85), .ZN(new_n421));
  INV_X1    g220(.A(new_n397), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT82), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n385), .A3(new_n386), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n396), .B1(new_n425), .B2(new_n314), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n421), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n419), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT86), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n308), .A2(new_n312), .A3(new_n313), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n376), .A2(new_n360), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(KEYINPUT39), .C1(new_n361), .C2(new_n366), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n319), .C1(KEYINPUT39), .C2(new_n432), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT40), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n435), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n430), .A2(new_n378), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n306), .B1(new_n305), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n310), .A2(new_n311), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n439), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT38), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT38), .B1(new_n296), .B2(KEYINPUT37), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n440), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n443), .A2(new_n301), .A3(new_n307), .A4(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n378), .A2(new_n382), .A3(new_n381), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n386), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n260), .B(new_n438), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n420), .A2(new_n429), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n260), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n451), .A2(new_n415), .A3(new_n416), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n395), .A2(new_n397), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT35), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n430), .A2(KEYINPUT35), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n448), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n450), .A2(new_n457), .ZN(new_n458));
  NOR3_X1   g257(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT89), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT90), .ZN(new_n463));
  INV_X1    g262(.A(G43gat), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT15), .B1(new_n464), .B2(G50gat), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n464), .B2(G50gat), .ZN(new_n466));
  INV_X1    g265(.A(G29gat), .ZN(new_n467));
  INV_X1    g266(.A(G36gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(G50gat), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT88), .B(G43gat), .Z(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(G50gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n466), .B(new_n469), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n459), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n466), .B1(new_n478), .B2(new_n469), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT17), .ZN(new_n483));
  XOR2_X1   g282(.A(G99gat), .B(G106gat), .Z(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT97), .ZN(new_n485));
  NAND2_X1  g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT7), .ZN(new_n487));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488));
  INV_X1    g287(.A(G85gat), .ZN(new_n489));
  INV_X1    g288(.A(G92gat), .ZN(new_n490));
  AOI22_X1  g289(.A1(KEYINPUT8), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n485), .B(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n483), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n480), .A2(new_n493), .ZN(new_n495));
  AND2_X1   g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(KEYINPUT41), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G190gat), .B(G218gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n496), .A2(KEYINPUT41), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT96), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n500), .B(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G134gat), .B(G162gat), .Z(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n500), .A2(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n502), .ZN(new_n507));
  INV_X1    g306(.A(new_n504), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(G71gat), .A2(G78gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(G71gat), .A2(G78gat), .ZN(new_n512));
  XOR2_X1   g311(.A(G57gat), .B(G64gat), .Z(new_n513));
  AOI211_X1 g312(.A(new_n511), .B(new_n512), .C1(new_n513), .C2(KEYINPUT9), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n511), .B1(KEYINPUT9), .B2(new_n512), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT94), .B(G57gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G64gat), .ZN(new_n517));
  INV_X1    g316(.A(G64gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G57gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT21), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G231gat), .A2(G233gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G127gat), .B(G155gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT95), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n528), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n533));
  AOI21_X1  g332(.A(G1gat), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n536), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n537), .A2(new_n538), .B1(KEYINPUT93), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(KEYINPUT93), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n540), .B(new_n541), .Z(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n523), .B2(new_n522), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n531), .B(new_n543), .Z(new_n544));
  XOR2_X1   g343(.A(G183gat), .B(G211gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n510), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n480), .A2(new_n542), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n483), .B2(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(KEYINPUT18), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n480), .B(new_n542), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n550), .B(KEYINPUT13), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT18), .B1(new_n549), .B2(new_n550), .ZN(new_n556));
  XOR2_X1   g355(.A(G113gat), .B(G141gat), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT11), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G169gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G197gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT12), .Z(new_n561));
  OR3_X1    g360(.A1(new_n555), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n555), .B2(new_n556), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT10), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n493), .A2(new_n566), .A3(new_n522), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n521), .A2(KEYINPUT98), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n521), .A2(KEYINPUT98), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n493), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(new_n493), .B2(new_n568), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n567), .B1(new_n571), .B2(new_n566), .ZN(new_n572));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n571), .B2(new_n573), .ZN(new_n576));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(G176gat), .B(G204gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n565), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n458), .A2(new_n547), .A3(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n425), .A2(KEYINPUT99), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n425), .A2(KEYINPUT99), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g389(.A1(new_n585), .A2(new_n430), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT16), .B(G8gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT42), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n592), .B(KEYINPUT101), .Z(new_n595));
  AOI22_X1  g394(.A1(new_n591), .A2(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n591), .B(KEYINPUT100), .Z(new_n597));
  NOR2_X1   g396(.A1(new_n593), .A2(G8gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(G1325gat));
  INV_X1    g398(.A(G15gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n415), .A2(new_n416), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n585), .A2(new_n419), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n600), .ZN(G1326gat));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n421), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT102), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT43), .B(G22gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(G1327gat));
  NAND2_X1  g407(.A1(new_n505), .A2(new_n509), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n584), .A2(new_n546), .ZN(new_n610));
  AOI211_X1 g409(.A(new_n609), .B(new_n610), .C1(new_n450), .C2(new_n457), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(new_n467), .A3(new_n588), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT45), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n450), .B2(new_n457), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT44), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n454), .A2(new_n456), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n427), .A2(new_n428), .A3(new_n449), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n510), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n619));
  OAI22_X1  g418(.A1(new_n614), .A2(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n588), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n621), .A2(new_n622), .A3(new_n610), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n613), .B1(new_n467), .B2(new_n623), .ZN(G1328gat));
  NAND3_X1  g423(.A1(new_n611), .A2(new_n468), .A3(new_n430), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT46), .Z(new_n626));
  NOR3_X1   g425(.A1(new_n621), .A2(new_n314), .A3(new_n610), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n468), .B2(new_n627), .ZN(G1329gat));
  NOR2_X1   g427(.A1(new_n621), .A2(new_n610), .ZN(new_n629));
  INV_X1    g428(.A(new_n471), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n419), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n611), .ZN(new_n632));
  INV_X1    g431(.A(new_n601), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n471), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g435(.A1(new_n262), .A2(G50gat), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT48), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n629), .A2(new_n451), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(new_n639), .B2(G50gat), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n632), .A2(new_n637), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n421), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(G50gat), .ZN(new_n646));
  OAI22_X1  g445(.A1(new_n642), .A2(new_n643), .B1(KEYINPUT48), .B2(new_n646), .ZN(G1331gat));
  NOR2_X1   g446(.A1(new_n616), .A2(new_n617), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n547), .A2(new_n565), .ZN(new_n650));
  INV_X1    g449(.A(new_n583), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n622), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n516), .ZN(G1332gat));
  INV_X1    g454(.A(KEYINPUT49), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n430), .B1(new_n656), .B2(new_n518), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT105), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n649), .A2(new_n652), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n518), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1333gat));
  OAI21_X1  g460(.A(G71gat), .B1(new_n653), .B2(new_n428), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n633), .A2(G71gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n653), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1334gat));
  NOR2_X1   g465(.A1(new_n653), .A2(new_n262), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT107), .B(G78gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1335gat));
  INV_X1    g468(.A(new_n546), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n670), .A2(new_n564), .A3(new_n651), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n615), .B1(new_n458), .B2(new_n510), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n618), .A2(new_n619), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n620), .A2(KEYINPUT108), .A3(new_n671), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G85gat), .B1(new_n678), .B2(new_n622), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n680), .B(new_n510), .C1(new_n616), .C2(new_n617), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n670), .A2(new_n564), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n618), .A2(KEYINPUT109), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT51), .ZN(new_n687));
  INV_X1    g486(.A(new_n685), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n683), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n690), .A2(KEYINPUT110), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(KEYINPUT110), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n583), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n588), .A2(new_n489), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n679), .B1(new_n693), .B2(new_n694), .ZN(G1336gat));
  NAND3_X1  g494(.A1(new_n430), .A2(new_n490), .A3(new_n583), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT111), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n686), .B2(new_n689), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT52), .ZN(new_n701));
  OAI21_X1  g500(.A(G92gat), .B1(new_n674), .B2(new_n314), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n620), .A2(KEYINPUT108), .A3(new_n671), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT108), .B1(new_n620), .B2(new_n671), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n704), .A2(new_n705), .A3(new_n314), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n700), .B1(new_n706), .B2(new_n490), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT112), .B1(new_n707), .B2(KEYINPUT52), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n676), .A2(new_n430), .A3(new_n677), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n699), .B1(new_n709), .B2(G92gat), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n711), .A3(new_n701), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n703), .B1(new_n708), .B2(new_n712), .ZN(G1337gat));
  OAI21_X1  g512(.A(G99gat), .B1(new_n678), .B2(new_n428), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n633), .A2(G99gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n693), .B2(new_n715), .ZN(G1338gat));
  NOR3_X1   g515(.A1(new_n651), .A2(new_n260), .A3(G106gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n690), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT53), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT113), .B(G106gat), .Z(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n674), .B2(new_n260), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n676), .A2(new_n421), .A3(new_n677), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n723), .A2(new_n720), .B1(new_n690), .B2(new_n717), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(new_n719), .ZN(G1339gat));
  OR3_X1    g524(.A1(new_n549), .A2(KEYINPUT114), .A3(new_n550), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT114), .B1(new_n549), .B2(new_n550), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n726), .B(new_n727), .C1(new_n552), .C2(new_n553), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n560), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(new_n562), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n572), .A2(new_n574), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n575), .A2(KEYINPUT54), .A3(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n732), .B(new_n579), .C1(KEYINPUT54), .C2(new_n575), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n735), .A2(new_n736), .A3(new_n580), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n510), .A2(new_n730), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n564), .A2(new_n737), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n729), .A2(new_n562), .A3(new_n583), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n609), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n743), .A2(new_n670), .B1(new_n583), .B2(new_n650), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(new_n314), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(new_n452), .A3(new_n588), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT115), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n332), .A3(new_n564), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n421), .A2(new_n633), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n745), .A2(new_n588), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G113gat), .B1(new_n750), .B2(new_n565), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1340gat));
  NAND3_X1  g551(.A1(new_n747), .A2(new_n335), .A3(new_n583), .ZN(new_n753));
  OAI21_X1  g552(.A(G120gat), .B1(new_n750), .B2(new_n651), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(G1341gat));
  NOR2_X1   g557(.A1(new_n746), .A2(new_n546), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n670), .A2(G127gat), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n759), .A2(G127gat), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT117), .ZN(G1342gat));
  INV_X1    g561(.A(new_n452), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n609), .A2(G134gat), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n745), .A2(new_n588), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G134gat), .B1(new_n750), .B2(new_n609), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(KEYINPUT118), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1343gat));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n650), .A2(new_n583), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n670), .B1(new_n738), .B2(new_n742), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n774), .B(new_n451), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n588), .A2(new_n314), .A3(new_n428), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT119), .Z(new_n779));
  AND2_X1   g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n740), .A2(KEYINPUT120), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n729), .A2(new_n782), .A3(new_n562), .A4(new_n583), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n739), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n781), .A2(KEYINPUT121), .A3(new_n739), .A4(new_n783), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n609), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n670), .B1(new_n788), .B2(new_n738), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n421), .B1(new_n789), .B2(new_n775), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT57), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n780), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n210), .B1(new_n793), .B2(new_n564), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n419), .A2(new_n260), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n745), .A2(new_n588), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n564), .A2(new_n210), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT58), .B1(new_n794), .B2(new_n798), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n792), .A2(KEYINPUT122), .A3(new_n565), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT122), .B1(new_n792), .B2(new_n565), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n210), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n798), .A2(KEYINPUT58), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(G1344gat));
  INV_X1    g603(.A(KEYINPUT123), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n805), .A3(new_n774), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n744), .A2(KEYINPUT57), .A3(new_n451), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n790), .B2(new_n774), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n583), .A3(new_n779), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n224), .A2(new_n226), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n796), .A2(new_n813), .A3(new_n651), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n792), .B2(new_n651), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n817), .ZN(G1345gat));
  OAI21_X1  g617(.A(G155gat), .B1(new_n792), .B2(new_n546), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n670), .A2(new_n204), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n796), .B2(new_n820), .ZN(G1346gat));
  OAI21_X1  g620(.A(G162gat), .B1(new_n792), .B2(new_n609), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n510), .A2(new_n205), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n796), .B2(new_n823), .ZN(G1347gat));
  NOR2_X1   g623(.A1(new_n588), .A2(new_n314), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n744), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n749), .ZN(new_n828));
  OAI21_X1  g627(.A(G169gat), .B1(new_n828), .B2(new_n565), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n826), .A2(new_n763), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n276), .A3(new_n564), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT124), .ZN(G1348gat));
  OAI21_X1  g632(.A(G176gat), .B1(new_n828), .B2(new_n651), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n277), .A3(new_n583), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1349gat));
  OAI21_X1  g635(.A(G183gat), .B1(new_n828), .B2(new_n546), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n830), .A2(new_n281), .A3(new_n670), .ZN(new_n838));
  NAND2_X1  g637(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n840), .B(new_n841), .Z(G1350gat));
  NAND3_X1  g641(.A1(new_n830), .A2(new_n282), .A3(new_n510), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(G190gat), .C1(new_n828), .C2(new_n609), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT126), .ZN(new_n846));
  OAI21_X1  g645(.A(G190gat), .B1(new_n828), .B2(new_n609), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT61), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n845), .A2(KEYINPUT126), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n843), .B1(new_n849), .B2(new_n850), .ZN(G1351gat));
  NAND2_X1  g650(.A1(new_n827), .A2(new_n795), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(G197gat), .B1(new_n853), .B2(new_n564), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n825), .A2(new_n428), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n810), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n564), .A2(G197gat), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(G1352gat));
  NAND3_X1  g658(.A1(new_n810), .A2(new_n583), .A3(new_n856), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G204gat), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT127), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n651), .A2(G204gat), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n852), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT127), .B(KEYINPUT62), .C1(new_n852), .C2(new_n863), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n866), .A2(new_n867), .B1(new_n865), .B2(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n861), .A2(new_n868), .ZN(G1353gat));
  OR3_X1    g668(.A1(new_n852), .A2(G211gat), .A3(new_n546), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n670), .B(new_n856), .C1(new_n808), .C2(new_n809), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n871), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT63), .B1(new_n871), .B2(G211gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(G1354gat));
  NAND3_X1  g673(.A1(new_n810), .A2(new_n510), .A3(new_n856), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G218gat), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n609), .A2(G218gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n852), .B2(new_n877), .ZN(G1355gat));
endmodule


