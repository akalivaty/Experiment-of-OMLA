//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n214), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n203), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n212), .B(new_n227), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n216), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n224), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n218), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n223), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G107), .ZN(new_n248));
  INV_X1    g0048(.A(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(new_n201), .ZN(new_n252));
  OAI21_X1  g0052(.A(G20), .B1(new_n252), .B2(new_n231), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT8), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT69), .B1(new_n258), .B2(G58), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n257), .B(new_n259), .C1(new_n260), .C2(KEYINPUT69), .ZN(new_n261));
  OR4_X1    g0061(.A1(KEYINPUT69), .A2(new_n257), .A3(new_n215), .A4(KEYINPUT8), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n229), .A2(G33), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n253), .B1(new_n254), .B2(new_n256), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n228), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n265), .A2(new_n271), .B1(new_n223), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n229), .A2(G1), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G50), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT67), .A2(G45), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT67), .A2(G45), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n272), .A3(G274), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G223), .A3(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G222), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n287), .B1(new_n202), .B2(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n228), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n285), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n296), .B1(new_n224), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n279), .B1(G179), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n299), .ZN(new_n302));
  INV_X1    g0102(.A(new_n279), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n303), .A2(KEYINPUT9), .B1(G200), .B2(new_n299), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n304), .B1(KEYINPUT9), .B2(new_n303), .C1(new_n305), .C2(new_n299), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n286), .A2(G232), .A3(G1698), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G97), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n311), .B(new_n312), .C1(new_n289), .C2(new_n224), .ZN(new_n313));
  INV_X1    g0113(.A(new_n298), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n295), .B1(G238), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n284), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n316), .B1(new_n315), .B2(new_n284), .ZN(new_n319));
  OAI21_X1  g0119(.A(G169), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT76), .A3(KEYINPUT14), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n315), .A2(new_n284), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n317), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(G169), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(G179), .A3(new_n317), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT77), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n328), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n321), .B(new_n326), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n274), .A2(KEYINPUT12), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n229), .A2(G68), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n256), .A2(new_n223), .B1(new_n264), .B2(new_n202), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n271), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT11), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT68), .B1(new_n266), .B2(new_n228), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n276), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(KEYINPUT72), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT12), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G68), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n273), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n272), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G68), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(KEYINPUT12), .A3(new_n348), .ZN(new_n349));
  AND4_X1   g0149(.A1(new_n332), .A2(new_n336), .A3(new_n343), .A4(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n331), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n324), .A2(G200), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n323), .A2(G190), .A3(new_n317), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n263), .A2(new_n274), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n339), .A2(new_n340), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n263), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n229), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NOR4_X1   g0165(.A1(new_n361), .A2(new_n362), .A3(new_n365), .A4(G20), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n215), .A2(new_n348), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n203), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n255), .A2(G159), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n367), .A2(new_n368), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n365), .B1(new_n286), .B2(G20), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n348), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n370), .A2(new_n371), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT16), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT78), .A2(KEYINPUT16), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n370), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n372), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n375), .A2(new_n376), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n339), .B1(new_n381), .B2(new_n378), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n360), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n294), .A2(G232), .A3(new_n297), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n284), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT80), .ZN(new_n386));
  OAI211_X1 g0186(.A(G226), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n387));
  OAI211_X1 g0187(.A(G223), .B(new_n288), .C1(new_n361), .C2(new_n362), .ZN(new_n388));
  INV_X1    g0188(.A(G33), .ZN(new_n389));
  INV_X1    g0189(.A(G87), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n387), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n295), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT80), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n284), .A2(new_n393), .A3(new_n384), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n386), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT79), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n391), .A2(new_n398), .A3(new_n295), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n398), .B1(new_n391), .B2(new_n295), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n386), .A2(new_n305), .A3(new_n394), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n397), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n383), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT17), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n383), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n380), .A2(new_n382), .ZN(new_n409));
  INV_X1    g0209(.A(new_n360), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G179), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n386), .A2(new_n412), .A3(new_n394), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n399), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n413), .A2(new_n415), .B1(new_n301), .B2(new_n395), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(KEYINPUT18), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n395), .A2(new_n301), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n418), .B1(new_n421), .B2(new_n383), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n406), .A2(new_n408), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n286), .A2(G238), .A3(G1698), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n286), .A2(G232), .A3(new_n288), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(new_n425), .C1(new_n217), .C2(new_n286), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n285), .B1(new_n426), .B2(new_n295), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n314), .A2(G244), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n301), .ZN(new_n430));
  INV_X1    g0230(.A(new_n429), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT75), .A3(new_n412), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n429), .B2(G179), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT15), .B(G87), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n436), .A2(new_n264), .B1(new_n260), .B2(new_n256), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n229), .A2(new_n202), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n271), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g0239(.A(new_n439), .B(KEYINPUT71), .Z(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT73), .B1(new_n341), .B2(new_n202), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT73), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n277), .A2(KEYINPUT72), .A3(new_n442), .A4(G77), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n441), .A2(new_n443), .B1(new_n202), .B2(new_n347), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(KEYINPUT74), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT74), .B1(new_n440), .B2(new_n444), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n430), .B(new_n435), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n431), .A2(G190), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n429), .A2(G200), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n449), .A2(new_n445), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n423), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n310), .A2(new_n353), .A3(new_n357), .A4(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(G257), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n455));
  OAI211_X1 g0255(.A(G250), .B(new_n288), .C1(new_n361), .C2(new_n362), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G294), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n295), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT5), .B(G41), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n460), .A2(new_n462), .B1(new_n292), .B2(new_n293), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G264), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n460), .A2(G274), .A3(new_n462), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n459), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G179), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT90), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n459), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n458), .A2(KEYINPUT90), .A3(new_n295), .ZN(new_n471));
  AND4_X1   g0271(.A1(new_n470), .A2(new_n464), .A3(new_n471), .A4(new_n465), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n468), .B1(new_n472), .B2(new_n301), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT88), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT22), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n286), .A2(new_n229), .A3(G87), .A4(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT23), .B1(new_n229), .B2(G107), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT89), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(KEYINPUT89), .B(KEYINPUT23), .C1(new_n229), .C2(G107), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n229), .A2(G107), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT23), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n477), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n229), .B(G87), .C1(new_n361), .C2(new_n362), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n474), .A2(new_n475), .ZN(new_n489));
  INV_X1    g0289(.A(new_n476), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n486), .A2(KEYINPUT24), .A3(new_n487), .A4(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n480), .A2(new_n481), .B1(new_n484), .B2(new_n483), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(new_n491), .A3(new_n487), .A4(new_n477), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT24), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n271), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n389), .A2(G1), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n337), .A2(new_n338), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(G107), .A3(new_n273), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n273), .A2(G107), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT25), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n497), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n473), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  NOR2_X1   g0305(.A1(KEYINPUT5), .A2(G41), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n462), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n507), .A2(G264), .A3(new_n294), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n459), .B2(new_n469), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(new_n305), .A3(new_n471), .A4(new_n465), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n466), .A2(new_n396), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(new_n500), .A3(new_n497), .A4(new_n502), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n514));
  OAI211_X1 g0314(.A(G238), .B(new_n288), .C1(new_n361), .C2(new_n362), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n295), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n272), .A2(G45), .A3(G274), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT83), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(new_n272), .A3(G45), .A4(G274), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n272), .A2(G45), .ZN(new_n524));
  AND2_X1   g0324(.A1(G33), .A2(G41), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(G250), .C1(new_n525), .C2(new_n228), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT84), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n526), .A2(KEYINPUT84), .A3(new_n520), .A4(new_n522), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G190), .B(new_n518), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n286), .A2(new_n229), .A3(G68), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n229), .B1(new_n312), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G87), .B2(new_n207), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n312), .B2(G20), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(new_n271), .B1(new_n347), .B2(new_n436), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n499), .A2(KEYINPUT85), .A3(G87), .A4(new_n273), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT85), .ZN(new_n539));
  INV_X1    g0339(.A(new_n498), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n269), .A2(new_n273), .A3(new_n270), .A4(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(new_n390), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n530), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n526), .A2(new_n520), .A3(new_n522), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT84), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n528), .B1(new_n295), .B2(new_n517), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n396), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n548), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n301), .ZN(new_n552));
  INV_X1    g0352(.A(new_n436), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n499), .A2(new_n273), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n548), .A2(new_n412), .B1(new_n537), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n544), .A2(new_n550), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n504), .A2(new_n513), .A3(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(new_n288), .C1(new_n361), .C2(new_n362), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G283), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G250), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT81), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n286), .A2(KEYINPUT81), .A3(G250), .A4(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n295), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n463), .A2(G257), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n465), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n301), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n569), .A2(new_n412), .A3(new_n465), .A4(new_n570), .ZN(new_n573));
  INV_X1    g0373(.A(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n274), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n499), .A2(G97), .A3(new_n273), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n217), .B1(new_n373), .B2(new_n374), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n256), .A2(new_n202), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT6), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n574), .A2(new_n217), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n579), .B1(new_n580), .B2(new_n206), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n229), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n577), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n575), .B(new_n576), .C1(new_n584), .C2(new_n339), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n572), .A2(new_n573), .A3(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n571), .A2(KEYINPUT82), .A3(G200), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT82), .B1(new_n571), .B2(G200), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n571), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n585), .B1(new_n590), .B2(G190), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n586), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n347), .A2(new_n249), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n266), .A2(new_n228), .B1(G20), .B2(new_n249), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n562), .B(new_n229), .C1(G33), .C2(new_n574), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n594), .A2(KEYINPUT20), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT20), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n269), .A2(new_n270), .A3(new_n540), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n345), .A2(G116), .A3(new_n346), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n301), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n507), .A2(G270), .A3(new_n294), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n604), .A2(new_n465), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(new_n288), .C1(new_n361), .C2(new_n362), .ZN(new_n606));
  INV_X1    g0406(.A(new_n362), .ZN(new_n607));
  NAND2_X1  g0407(.A1(KEYINPUT3), .A2(G33), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(G303), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G264), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n295), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT21), .B1(new_n603), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(G179), .A3(new_n612), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT86), .B1(new_n602), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n594), .A2(new_n595), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT20), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n594), .A2(KEYINPUT20), .A3(new_n595), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n345), .A2(G116), .A3(new_n346), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n499), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n623), .A3(new_n593), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n604), .A2(new_n465), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n295), .B2(new_n611), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT86), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n624), .A2(new_n626), .A3(new_n627), .A4(G179), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n624), .A2(new_n613), .A3(KEYINPUT21), .A4(G169), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n616), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n616), .A2(new_n628), .A3(new_n629), .A4(KEYINPUT87), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n614), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n613), .A2(G200), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n635), .B(new_n602), .C1(new_n305), .C2(new_n613), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n557), .A2(new_n592), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n454), .A2(new_n638), .ZN(G372));
  NOR2_X1   g0439(.A1(new_n630), .A2(new_n614), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n504), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n537), .A2(new_n554), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n412), .B(new_n518), .C1(new_n527), .C2(new_n529), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n551), .A2(KEYINPUT91), .A3(new_n301), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT91), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n548), .B2(G169), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n530), .A2(new_n537), .A3(new_n543), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n549), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n592), .A2(new_n641), .A3(new_n513), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n586), .A2(new_n556), .A3(KEYINPUT26), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n572), .A2(new_n573), .A3(new_n585), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n648), .A2(new_n654), .A3(new_n650), .ZN(new_n655));
  OAI211_X1 g0455(.A(KEYINPUT92), .B(new_n653), .C1(new_n655), .C2(KEYINPUT26), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n653), .A2(KEYINPUT92), .ZN(new_n657));
  INV_X1    g0457(.A(new_n648), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n652), .A2(new_n656), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n454), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n406), .A2(new_n408), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n357), .A2(new_n448), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n353), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n417), .A2(new_n422), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n307), .A2(new_n308), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n302), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n660), .A2(new_n667), .ZN(G369));
  XOR2_X1   g0468(.A(KEYINPUT93), .B(G330), .Z(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G13), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n272), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n634), .B(new_n636), .C1(new_n602), .C2(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n624), .B(new_n678), .C1(new_n630), .C2(new_n614), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n670), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n504), .A2(new_n513), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n503), .A2(new_n678), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n683), .A2(new_n684), .B1(new_n504), .B2(new_n679), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n634), .A2(new_n504), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n513), .A3(new_n679), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n210), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n232), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n548), .A2(new_n459), .A3(new_n464), .ZN(new_n697));
  INV_X1    g0497(.A(new_n615), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n590), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n467), .A2(G179), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(new_n551), .A3(new_n571), .A4(new_n613), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n590), .A2(new_n697), .A3(KEYINPUT30), .A4(new_n698), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n678), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT31), .B(new_n706), .C1(new_n637), .C2(new_n678), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n706), .A2(KEYINPUT31), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n669), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n707), .A2(KEYINPUT94), .A3(new_n669), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT26), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n586), .A2(new_n556), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n651), .A2(new_n586), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n648), .B1(new_n718), .B2(KEYINPUT26), .ZN(new_n719));
  INV_X1    g0519(.A(new_n687), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n592), .A2(new_n513), .A3(new_n651), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n717), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n715), .B1(new_n722), .B2(new_n679), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n659), .A2(new_n679), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n723), .B1(new_n715), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n714), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n696), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n690), .A2(new_n286), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n281), .A2(new_n282), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n233), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n730), .B(new_n732), .C1(new_n246), .C2(new_n461), .ZN(new_n733));
  INV_X1    g0533(.A(G355), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n286), .A2(new_n210), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n733), .B1(G116), .B2(new_n210), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n228), .B1(G20), .B2(new_n301), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT96), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n272), .B1(new_n672), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n691), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT95), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n229), .A2(new_n305), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n412), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n229), .A2(G190), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G179), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G322), .A2(new_n751), .B1(new_n755), .B2(G329), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n396), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G303), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n752), .A2(new_n757), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n761), .B1(G283), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n229), .B1(new_n753), .B2(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G294), .ZN(new_n767));
  NAND3_X1  g0567(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n305), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n363), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n752), .A2(new_n749), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(G311), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n768), .A2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(G317), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT33), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(KEYINPUT33), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n764), .A2(new_n767), .A3(new_n775), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n754), .A2(KEYINPUT32), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT32), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n755), .B2(G159), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(G68), .C2(new_n776), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n786), .B1(new_n223), .B2(new_n770), .C1(new_n574), .C2(new_n765), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G58), .A2(new_n751), .B1(new_n763), .B2(G107), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n759), .A2(G87), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n774), .A2(G77), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n788), .A2(new_n286), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n781), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n747), .B1(new_n792), .B2(new_n738), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n680), .A2(new_n681), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n741), .B(KEYINPUT97), .Z(new_n795));
  OAI211_X1 g0595(.A(new_n743), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n682), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n747), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n794), .A2(new_n669), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT98), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  AOI22_X1  g0602(.A1(new_n449), .A2(new_n445), .B1(new_n301), .B2(new_n429), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT100), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n803), .A2(new_n804), .A3(new_n435), .A4(new_n678), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT100), .B1(new_n448), .B2(new_n679), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n678), .B1(new_n446), .B2(new_n447), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n448), .A2(new_n452), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n724), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n659), .A2(new_n809), .A3(new_n679), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n713), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n747), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n774), .A2(G159), .B1(G137), .B2(new_n769), .ZN(new_n816));
  INV_X1    g0616(.A(G143), .ZN(new_n817));
  INV_X1    g0617(.A(new_n776), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n816), .B1(new_n817), .B2(new_n750), .C1(new_n254), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n763), .A2(G68), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n286), .B1(new_n754), .B2(new_n822), .C1(new_n223), .C2(new_n758), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G58), .B2(new_n766), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n770), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n363), .B1(new_n758), .B2(new_n217), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT99), .Z(new_n829));
  NOR2_X1   g0629(.A1(new_n762), .A2(new_n390), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n773), .A2(new_n249), .B1(new_n754), .B2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n830), .B(new_n832), .C1(G294), .C2(new_n751), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n766), .A2(G97), .B1(G283), .B2(new_n776), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n829), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n825), .B1(new_n827), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n747), .B1(new_n836), .B2(new_n738), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n738), .A2(new_n739), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(G77), .B2(new_n839), .C1(new_n809), .C2(new_n740), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n815), .A2(new_n840), .ZN(G384));
  INV_X1    g0641(.A(KEYINPUT40), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n351), .A2(new_n678), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n352), .A2(new_n356), .A3(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n351), .B(new_n678), .C1(new_n331), .C2(new_n357), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g0646(.A1(new_n707), .A2(new_n846), .A3(new_n708), .A4(new_n809), .ZN(new_n847));
  XOR2_X1   g0647(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n848));
  INV_X1    g0648(.A(new_n676), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n411), .B1(new_n416), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n405), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n411), .A2(new_n849), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n423), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n848), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n339), .B1(new_n372), .B2(new_n377), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n849), .B1(new_n857), .B2(new_n360), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n419), .B(new_n420), .C1(new_n857), .C2(new_n360), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n405), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n850), .A2(new_n852), .A3(new_n405), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(KEYINPUT38), .C1(new_n423), .C2(new_n858), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT104), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n661), .A2(new_n664), .ZN(new_n866));
  INV_X1    g0666(.A(new_n858), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT104), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT38), .A4(new_n863), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n856), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n842), .B1(new_n847), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n864), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n868), .B2(new_n863), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n842), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n707), .A2(new_n708), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n809), .A3(new_n846), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n454), .A2(new_n877), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n669), .ZN(new_n884));
  INV_X1    g0684(.A(new_n726), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n454), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n667), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n856), .A2(new_n865), .A3(new_n888), .A4(new_n870), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT39), .B1(new_n873), .B2(new_n874), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n352), .A2(new_n678), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n417), .A2(new_n422), .A3(new_n676), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n803), .A2(new_n435), .A3(new_n679), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n812), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n875), .A2(new_n896), .A3(new_n846), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n887), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n884), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n272), .B2(new_n672), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n232), .A2(new_n202), .A3(new_n369), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n252), .A2(new_n348), .ZN(new_n903));
  OAI211_X1 g0703(.A(G1), .B(new_n671), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n581), .A2(new_n582), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT101), .Z(new_n906));
  AOI21_X1  g0706(.A(new_n249), .B1(new_n906), .B2(KEYINPUT35), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n907), .B(new_n230), .C1(KEYINPUT35), .C2(new_n906), .ZN(new_n908));
  XOR2_X1   g0708(.A(KEYINPUT102), .B(KEYINPUT36), .Z(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n901), .A2(new_n904), .A3(new_n910), .ZN(G367));
  INV_X1    g0711(.A(G283), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n773), .A2(new_n912), .B1(new_n765), .B2(new_n217), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT111), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n759), .A2(G116), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT46), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n776), .A2(G294), .B1(new_n769), .B2(G311), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n286), .B1(new_n763), .B2(G97), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n755), .A2(G317), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n914), .B(new_n920), .C1(G303), .C2(new_n751), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT112), .Z(new_n922));
  NOR2_X1   g0722(.A1(new_n762), .A2(new_n202), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n215), .A2(new_n758), .B1(new_n750), .B2(new_n254), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(G137), .C2(new_n755), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n765), .A2(new_n348), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n286), .B1(new_n770), .B2(new_n817), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(G159), .C2(new_n776), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n925), .B(new_n928), .C1(new_n201), .C2(new_n773), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT47), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n747), .B1(new_n931), .B2(new_n738), .ZN(new_n932));
  INV_X1    g0732(.A(new_n730), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n742), .B1(new_n210), .B2(new_n436), .C1(new_n241), .C2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n679), .B1(new_n537), .B2(new_n543), .ZN(new_n935));
  MUX2_X1   g0735(.A(new_n651), .B(new_n648), .S(new_n935), .Z(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT106), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n932), .B(new_n934), .C1(new_n795), .C2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n634), .A2(new_n678), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(new_n504), .A3(new_n513), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n685), .B2(new_n939), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(new_n682), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n726), .A2(new_n711), .A3(new_n942), .A4(new_n712), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT108), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT45), .ZN(new_n946));
  INV_X1    g0746(.A(new_n688), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n654), .A2(new_n679), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT107), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n585), .A2(new_n678), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n592), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n946), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n953), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(KEYINPUT45), .A3(new_n688), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n954), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n956), .B2(new_n688), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n958), .A2(new_n686), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n686), .B1(new_n958), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n714), .A2(KEYINPUT108), .A3(new_n726), .A4(new_n942), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n945), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT109), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n945), .A2(new_n965), .A3(new_n966), .A4(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n728), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n691), .B(KEYINPUT41), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(KEYINPUT110), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT110), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n727), .B1(new_n969), .B2(new_n970), .ZN(new_n976));
  INV_X1    g0776(.A(new_n973), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n745), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n954), .A2(new_n940), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT42), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n654), .B1(new_n954), .B2(new_n504), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n679), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n981), .A2(new_n983), .B1(KEYINPUT43), .B2(new_n937), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n686), .A2(new_n954), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n984), .B(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n938), .B1(new_n979), .B2(new_n988), .ZN(G387));
  AOI22_X1  g0789(.A1(new_n774), .A2(G303), .B1(G322), .B2(new_n769), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n831), .B2(new_n818), .C1(new_n777), .C2(new_n750), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT48), .ZN(new_n992));
  INV_X1    g0792(.A(G294), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n912), .B2(new_n765), .C1(new_n993), .C2(new_n758), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT49), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n363), .B1(new_n754), .B2(new_n771), .C1(new_n249), .C2(new_n762), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT115), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n995), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n997), .A2(KEYINPUT115), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n766), .A2(new_n553), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n223), .B2(new_n750), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT114), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G97), .B2(new_n763), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n263), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n776), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n758), .A2(new_n202), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G150), .B2(new_n755), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n348), .B2(new_n773), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G159), .B2(new_n769), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1005), .A2(new_n286), .A3(new_n1007), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1001), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n747), .B1(new_n1013), .B2(new_n738), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n685), .B2(new_n795), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n260), .A2(G50), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT50), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n348), .A2(new_n202), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT113), .ZN(new_n1019));
  AOI211_X1 g0819(.A(G45), .B(new_n1018), .C1(new_n693), .C2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1017), .B(new_n1020), .C1(new_n1019), .C2(new_n693), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n730), .B(new_n1021), .C1(new_n238), .C2(new_n731), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(G107), .B2(new_n210), .C1(new_n693), .C2(new_n735), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1015), .B1(new_n742), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT116), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n745), .B2(new_n942), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n945), .A2(new_n966), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n728), .B2(new_n942), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1028), .B2(new_n692), .ZN(G393));
  INV_X1    g0829(.A(new_n965), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n969), .A2(new_n970), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1031), .A2(new_n691), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n742), .B1(new_n574), .B2(new_n210), .C1(new_n250), .C2(new_n933), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G68), .A2(new_n759), .B1(new_n755), .B2(G143), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n766), .A2(G77), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n260), .C2(new_n773), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n286), .B1(new_n762), .B2(new_n390), .C1(new_n818), .C2(new_n201), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n751), .A2(G159), .B1(G150), .B2(new_n769), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n770), .A2(new_n777), .B1(new_n750), .B2(new_n831), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT52), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G283), .A2(new_n759), .B1(new_n755), .B2(G322), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n286), .B1(new_n766), .B2(G116), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n763), .A2(G107), .B1(G303), .B2(new_n776), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n773), .A2(new_n993), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1038), .A2(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n747), .B1(new_n1048), .B2(new_n738), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n741), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1033), .B(new_n1049), .C1(new_n956), .C2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1030), .B2(new_n744), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1032), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(G390));
  NAND2_X1  g0854(.A1(new_n896), .A2(new_n846), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n892), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n889), .A2(new_n890), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n871), .A2(new_n1056), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n722), .A2(new_n679), .A3(new_n809), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n895), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n846), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1057), .A2(new_n1058), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT117), .ZN(new_n1064));
  AND4_X1   g0864(.A1(new_n1064), .A2(new_n713), .A3(new_n809), .A4(new_n846), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n810), .B1(new_n711), .B2(new_n712), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1064), .B1(new_n1066), .B2(new_n846), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1063), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1068), .A2(KEYINPUT118), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT118), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n713), .A2(new_n809), .A3(new_n846), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(KEYINPUT117), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1066), .A2(new_n1064), .A3(new_n846), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1070), .B1(new_n1074), .B2(new_n1063), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1063), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(G330), .A3(new_n847), .ZN(new_n1078));
  INV_X1    g0878(.A(G330), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n667), .B(new_n886), .C1(new_n882), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1061), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n877), .A2(new_n809), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n846), .B1(new_n1083), .B2(G330), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1082), .B(new_n1085), .C1(new_n1065), .C2(new_n1067), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1066), .A2(new_n846), .B1(new_n1079), .B2(new_n878), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1087), .A2(KEYINPUT119), .A3(new_n896), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT119), .B1(new_n1087), .B2(new_n896), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1076), .A2(new_n1078), .A3(new_n1081), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1081), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1068), .A2(KEYINPUT118), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1074), .A2(new_n1070), .A3(new_n1063), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n1078), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n691), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT120), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1091), .A2(new_n1096), .A3(KEYINPUT120), .A4(new_n691), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1093), .A2(new_n1094), .A3(new_n1078), .A4(new_n745), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n821), .B1(new_n249), .B2(new_n750), .C1(new_n993), .C2(new_n754), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G97), .B2(new_n774), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n776), .A2(G107), .B1(new_n769), .B2(G283), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n789), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1104), .A2(new_n363), .A3(new_n1035), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n770), .A2(new_n1108), .B1(new_n750), .B2(new_n822), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT121), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n286), .B1(new_n754), .B2(new_n1111), .C1(new_n201), .C2(new_n762), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT54), .B(G143), .Z(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n774), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n766), .A2(G159), .B1(G137), .B2(new_n776), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1110), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n759), .A2(G150), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1107), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n747), .B1(new_n1119), .B2(new_n738), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n1006), .B2(new_n839), .C1(new_n891), .C2(new_n740), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1102), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1101), .A2(new_n1123), .ZN(G378));
  NAND2_X1  g0924(.A1(new_n1087), .A2(new_n896), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1087), .A2(KEYINPUT119), .A3(new_n896), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1084), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1127), .A2(new_n1128), .B1(new_n1129), .B2(new_n1082), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1081), .B1(new_n1095), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n898), .B1(new_n880), .B2(new_n1079), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1133), .B(G330), .C1(new_n872), .C2(new_n879), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n303), .A2(new_n676), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n310), .A2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n302), .B(new_n1136), .C1(new_n307), .C2(new_n308), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT55), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1136), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n309), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT55), .B1(new_n1143), .B2(new_n1138), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1141), .A2(KEYINPUT56), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT56), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1135), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1131), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1131), .A2(new_n1151), .A3(KEYINPUT57), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n691), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n744), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1149), .A2(new_n739), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n838), .A2(new_n201), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n759), .A2(KEYINPUT122), .A3(new_n1113), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n774), .A2(G137), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n1108), .C2(new_n750), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT122), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1113), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n758), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n254), .B2(new_n765), .C1(new_n822), .C2(new_n818), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1162), .B(new_n1166), .C1(G125), .C2(new_n769), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT59), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G41), .B1(new_n763), .B2(G159), .ZN(new_n1169));
  INV_X1    g0969(.A(G124), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n754), .B1(KEYINPUT123), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(KEYINPUT123), .B2(new_n1170), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n389), .A3(new_n1169), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n223), .B1(new_n361), .B2(G41), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n926), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n770), .B2(new_n249), .C1(new_n574), .C2(new_n818), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1176), .A2(G41), .A3(new_n286), .A4(new_n1008), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n762), .A2(new_n215), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n436), .B2(new_n773), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G107), .B2(new_n751), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1177), .B(new_n1181), .C1(new_n912), .C2(new_n754), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT58), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1173), .A2(new_n1174), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n747), .B1(new_n1184), .B2(new_n738), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1158), .A2(new_n1159), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1157), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1156), .A2(new_n1187), .ZN(G375));
  INV_X1    g0988(.A(KEYINPUT124), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1130), .B2(new_n744), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n773), .A2(new_n254), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n758), .A2(new_n782), .B1(new_n754), .B2(new_n1108), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(G137), .C2(new_n751), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1164), .A2(new_n818), .B1(new_n223), .B2(new_n765), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G132), .B2(new_n769), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1193), .A2(new_n286), .A3(new_n1179), .A4(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n773), .A2(new_n217), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n574), .A2(new_n758), .B1(new_n750), .B2(new_n912), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(G303), .C2(new_n755), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n818), .A2(new_n249), .B1(new_n770), .B2(new_n993), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(new_n923), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1002), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1196), .B1(new_n1202), .B2(new_n286), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n747), .B1(new_n1203), .B2(new_n738), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(G68), .B2(new_n839), .C1(new_n846), .C2(new_n740), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1090), .A2(KEYINPUT124), .A3(new_n745), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1190), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1080), .B(new_n1086), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1092), .A2(new_n973), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(G381));
  NAND2_X1  g1011(.A1(new_n1097), .A2(new_n1123), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G375), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(G393), .A2(G396), .ZN(new_n1215));
  OR3_X1    g1015(.A1(G387), .A2(G390), .A3(new_n1215), .ZN(new_n1216));
  OR4_X1    g1016(.A1(G384), .A2(new_n1214), .A3(G381), .A4(new_n1216), .ZN(G407));
  OAI211_X1 g1017(.A(G407), .B(G213), .C1(G343), .C2(new_n1214), .ZN(G409));
  INV_X1    g1018(.A(new_n1212), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1131), .A2(new_n1151), .A3(new_n973), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1187), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1122), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(G375), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G213), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(G343), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(G384), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT60), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1209), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n691), .A3(new_n1092), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1209), .B2(new_n1229), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1130), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1080), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1231), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1228), .B1(new_n1235), .B2(new_n1207), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1208), .B(G384), .C1(new_n1237), .C2(new_n1231), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1224), .A2(new_n1227), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT62), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1226), .A2(G2897), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1236), .A2(new_n1238), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1243), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1212), .B1(new_n1187), .B2(new_n1220), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1187), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n692), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1155), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1248), .B1(G378), .B2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1244), .B(new_n1247), .C1(new_n1252), .C2(new_n1226), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1224), .A2(new_n1254), .A3(new_n1239), .A4(new_n1227), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1241), .A2(new_n1242), .A3(new_n1253), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(new_n1053), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G390), .B(new_n938), .C1(new_n979), .C2(new_n988), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G393), .A2(G396), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT126), .B1(new_n1215), .B2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1215), .A2(new_n1259), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1263));
  AND3_X1   g1063(.A1(G387), .A2(KEYINPUT126), .A3(new_n1053), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1261), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1256), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1257), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1224), .A2(KEYINPUT63), .A3(new_n1239), .A4(new_n1227), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1244), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1243), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1271), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1240), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1269), .B(new_n1270), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1266), .A2(new_n1278), .ZN(G405));
  NOR2_X1   g1079(.A1(G375), .A2(new_n1223), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1251), .A2(new_n1212), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1239), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G378), .A2(new_n1251), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G375), .A2(new_n1219), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n1284), .A3(new_n1245), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1267), .A2(new_n1282), .A3(new_n1268), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1265), .A2(KEYINPUT127), .A3(new_n1282), .A4(new_n1285), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1288), .A2(new_n1291), .A3(new_n1292), .ZN(G402));
endmodule


