//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT41), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  AND2_X1   g004(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT83), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT83), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G50gat), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT84), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n212), .ZN(new_n221));
  NAND2_X1  g020(.A1(G43gat), .A2(G50gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n211), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n217), .A2(new_n227), .A3(new_n218), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n210), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G99gat), .ZN(new_n232));
  INV_X1    g031(.A(G106gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G99gat), .A2(G106gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT95), .ZN(new_n237));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT7), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT95), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n234), .A2(new_n240), .A3(new_n235), .ZN(new_n241));
  INV_X1    g040(.A(G85gat), .ZN(new_n242));
  INV_X1    g041(.A(G92gat), .ZN(new_n243));
  AOI22_X1  g042(.A1(KEYINPUT8), .A2(new_n235), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND4_X1   g043(.A1(new_n237), .A2(new_n239), .A3(new_n241), .A4(new_n244), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n237), .A2(new_n241), .B1(new_n239), .B2(new_n244), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n204), .B1(new_n231), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n229), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n224), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n227), .B1(new_n217), .B2(new_n218), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n229), .B1(new_n251), .B2(new_n226), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n250), .A2(KEYINPUT17), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT17), .B1(new_n250), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n248), .B1(new_n255), .B2(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT96), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT96), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(new_n248), .C1(new_n255), .C2(new_n247), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n261), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n202), .A2(new_n203), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT94), .ZN(new_n267));
  XNOR2_X1  g066(.A(G190gat), .B(G218gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n262), .A2(new_n269), .A3(new_n264), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(G71gat), .B2(G78gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G64gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(G71gat), .A2(G78gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G71gat), .A2(G78gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  OAI221_X1 g082(.A(new_n276), .B1(new_n280), .B2(new_n281), .C1(new_n277), .C2(new_n278), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(KEYINPUT21), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G1gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT16), .ZN(new_n290));
  INV_X1    g089(.A(G15gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G22gat), .ZN(new_n292));
  INV_X1    g091(.A(G22gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G15gat), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(G1gat), .B1(new_n292), .B2(new_n294), .ZN(new_n296));
  OAI21_X1  g095(.A(G8gat), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n298));
  INV_X1    g097(.A(G8gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(G15gat), .B(G22gat), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n298), .B(new_n299), .C1(G1gat), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(KEYINPUT21), .B2(new_n285), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n288), .B(new_n303), .Z(new_n304));
  XNOR2_X1  g103(.A(G127gat), .B(G155gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT20), .ZN(new_n306));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n307), .B(KEYINPUT92), .Z(new_n308));
  XNOR2_X1  g107(.A(new_n306), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G183gat), .B(G211gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n304), .B(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n274), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n283), .B(new_n284), .C1(new_n245), .C2(new_n246), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n237), .A2(new_n239), .A3(new_n241), .A4(new_n244), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n237), .A2(new_n241), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n239), .A2(new_n244), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n285), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT10), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n247), .A2(KEYINPUT10), .A3(new_n285), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT97), .ZN(new_n324));
  NAND2_X1  g123(.A1(G230gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT97), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n326), .A3(new_n322), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n325), .B1(new_n314), .B2(new_n319), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n329), .A2(KEYINPUT98), .ZN(new_n330));
  XNOR2_X1  g129(.A(G120gat), .B(G148gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G176gat), .B(G204gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n329), .B2(KEYINPUT98), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT99), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n323), .B2(new_n325), .ZN(new_n338));
  INV_X1    g137(.A(new_n325), .ZN(new_n339));
  AOI211_X1 g138(.A(KEYINPUT99), .B(new_n339), .C1(new_n321), .C2(new_n322), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n338), .A2(new_n340), .A3(new_n329), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n336), .B1(new_n341), .B2(new_n333), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n313), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT64), .B(KEYINPUT24), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT66), .B(G183gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(G190gat), .ZN(new_n347));
  INV_X1    g146(.A(G183gat), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT65), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT23), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n358), .A2(G169gat), .A3(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n357), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n362), .A2(KEYINPUT25), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n353), .B1(new_n366), .B2(new_n350), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT25), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n370));
  NOR2_X1   g169(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n346), .B2(KEYINPUT27), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n372), .B2(G190gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT27), .B(G183gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(KEYINPUT28), .A3(new_n349), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n361), .A2(new_n356), .A3(KEYINPUT26), .ZN(new_n377));
  AOI211_X1 g176(.A(new_n350), .B(new_n377), .C1(KEYINPUT26), .C2(new_n356), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n364), .A2(new_n369), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G127gat), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT67), .B1(new_n380), .B2(G134gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G113gat), .B(G120gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(KEYINPUT1), .ZN(new_n383));
  XNOR2_X1  g182(.A(G127gat), .B(G134gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n383), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n383), .B(new_n384), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n376), .A2(new_n378), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n368), .B1(new_n355), .B2(new_n363), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G227gat), .A2(G233gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT34), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT34), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n387), .A2(new_n391), .A3(new_n395), .A4(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n398));
  INV_X1    g197(.A(new_n392), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n389), .A2(new_n390), .A3(new_n388), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n364), .A2(new_n369), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n376), .A2(new_n378), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n386), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n399), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405));
  XNOR2_X1  g204(.A(G15gat), .B(G43gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT68), .ZN(new_n407));
  XNOR2_X1  g206(.A(G71gat), .B(G99gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n410), .B2(new_n409), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(KEYINPUT32), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT71), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n404), .A2(new_n415), .A3(KEYINPUT32), .A4(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n404), .A2(new_n405), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n404), .A2(KEYINPUT32), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT69), .A4(new_n409), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT69), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n392), .B1(new_n387), .B2(new_n391), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n409), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(KEYINPUT33), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n398), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n418), .A2(new_n419), .A3(new_n409), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n431), .A2(new_n422), .B1(KEYINPUT72), .B2(new_n397), .ZN(new_n432));
  INV_X1    g231(.A(new_n398), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n420), .A4(new_n417), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436));
  XNOR2_X1  g235(.A(G197gat), .B(G204gat), .ZN(new_n437));
  INV_X1    g236(.A(G211gat), .ZN(new_n438));
  INV_X1    g237(.A(G218gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(KEYINPUT22), .B2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G211gat), .B(G218gat), .Z(new_n442));
  AND2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n441), .A2(new_n442), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n436), .B1(new_n445), .B2(KEYINPUT29), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n447));
  XNOR2_X1  g246(.A(G141gat), .B(G148gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT2), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(G155gat), .B2(G162gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g250(.A(G155gat), .B(G162gat), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n451), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n451), .A2(new_n452), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n451), .A2(new_n452), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n436), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n445), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G228gat), .ZN(new_n463));
  INV_X1    g262(.A(G233gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n441), .B(new_n442), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n458), .B2(new_n459), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n462), .B(new_n466), .C1(KEYINPUT77), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT77), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n455), .B(new_n461), .C1(new_n470), .C2(new_n465), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n293), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT78), .ZN(new_n473));
  XNOR2_X1  g272(.A(G78gat), .B(G106gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G50gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n471), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n468), .B1(new_n454), .B2(new_n446), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n466), .B1(new_n468), .B2(KEYINPUT77), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(G22gat), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n473), .A2(new_n476), .B1(new_n472), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT78), .ZN(new_n483));
  AND4_X1   g282(.A1(new_n483), .A2(new_n481), .A3(new_n472), .A4(new_n476), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n435), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G8gat), .B(G36gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G226gat), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n379), .A2(KEYINPUT29), .B1(new_n492), .B2(new_n464), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n401), .A2(new_n402), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n492), .A2(new_n464), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n467), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n467), .B1(new_n493), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n491), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n495), .B1(new_n494), .B2(new_n459), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n379), .A2(new_n492), .A3(new_n464), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n445), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n503), .A2(KEYINPUT30), .A3(new_n490), .A4(new_n497), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT73), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n500), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n490), .A3(new_n497), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G1gat), .B(G29gat), .Z(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G57gat), .B(G85gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n386), .B1(new_n456), .B2(new_n457), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n388), .A2(new_n454), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n518), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n454), .A2(KEYINPUT3), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n458), .A3(new_n388), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT4), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n388), .B2(new_n454), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n386), .B(KEYINPUT4), .C1(new_n456), .C2(new_n457), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n526), .A2(new_n522), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n528), .A2(new_n529), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(new_n518), .A3(new_n522), .A4(new_n526), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n531), .B1(new_n524), .B2(new_n530), .ZN(new_n536));
  OAI211_X1 g335(.A(KEYINPUT6), .B(new_n517), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n524), .A2(new_n530), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT75), .ZN(new_n540));
  INV_X1    g339(.A(new_n517), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n534), .A4(new_n532), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n534), .A3(new_n532), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n517), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n538), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n512), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT35), .B1(new_n487), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(KEYINPUT80), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT80), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n540), .A2(new_n551), .A3(new_n534), .A4(new_n532), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n517), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n538), .B1(new_n553), .B2(new_n544), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n511), .A2(new_n500), .A3(new_n504), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT81), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n485), .B1(new_n430), .B2(new_n434), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n559));
  INV_X1    g358(.A(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n543), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n541), .B1(new_n545), .B2(KEYINPUT80), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n552), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n559), .B(new_n560), .C1(new_n563), .C2(new_n538), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n430), .A2(KEYINPUT36), .A3(new_n434), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT36), .B1(new_n430), .B2(new_n434), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT37), .B1(new_n498), .B2(new_n499), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n503), .A2(new_n571), .A3(new_n497), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n491), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n573), .A2(KEYINPUT38), .ZN(new_n574));
  INV_X1    g373(.A(new_n509), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n573), .B2(KEYINPUT38), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n523), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(KEYINPUT79), .A3(new_n523), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT39), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(new_n517), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT40), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n581), .A2(KEYINPUT39), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n584), .B2(new_n587), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n555), .B(new_n553), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n577), .A2(new_n486), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n485), .B1(new_n512), .B2(new_n547), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n569), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n566), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT82), .B(G197gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT11), .B(G169gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT86), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n250), .A2(new_n302), .A3(new_n252), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n225), .B2(new_n230), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n250), .A2(KEYINPUT17), .A3(new_n252), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n302), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n603), .B1(new_n612), .B2(KEYINPUT18), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n253), .B2(new_n254), .ZN(new_n614));
  INV_X1    g413(.A(new_n606), .ZN(new_n615));
  AND4_X1   g414(.A1(new_n603), .A2(new_n614), .A3(KEYINPUT18), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n618));
  AOI21_X1  g417(.A(new_n302), .B1(new_n608), .B2(new_n609), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(new_n606), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT13), .Z(new_n621));
  AOI21_X1  g420(.A(new_n302), .B1(new_n250), .B2(new_n252), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT87), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n604), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI211_X1 g423(.A(KEYINPUT87), .B(new_n302), .C1(new_n250), .C2(new_n252), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n602), .B1(new_n617), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n614), .A2(KEYINPUT18), .A3(new_n615), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT86), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n603), .A3(KEYINPUT18), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n620), .A2(new_n626), .A3(new_n601), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT88), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT88), .B1(new_n632), .B2(new_n633), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n628), .B(KEYINPUT89), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT88), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n620), .A2(new_n626), .A3(new_n601), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n617), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT88), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT89), .B1(new_n642), .B2(new_n628), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n594), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT90), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT90), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n594), .A2(new_n648), .A3(new_n645), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n344), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n547), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT100), .B(G1gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1324gat));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT16), .B(G8gat), .Z(new_n655));
  NAND4_X1  g454(.A1(new_n650), .A2(new_n654), .A3(new_n555), .A4(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n344), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n648), .B1(new_n594), .B2(new_n645), .ZN(new_n658));
  AOI211_X1 g457(.A(KEYINPUT90), .B(new_n644), .C1(new_n566), .C2(new_n593), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n555), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n655), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT42), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n664));
  INV_X1    g463(.A(new_n660), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n665), .B2(new_n299), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n660), .A2(KEYINPUT101), .A3(G8gat), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n663), .A2(new_n670), .A3(new_n666), .A4(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(G1325gat));
  INV_X1    g471(.A(new_n650), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n569), .B(KEYINPUT103), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G15gat), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n650), .A2(new_n291), .A3(new_n435), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n650), .A2(new_n485), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n592), .A2(KEYINPUT105), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n685), .B(new_n485), .C1(new_n512), .C2(new_n547), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n569), .A2(new_n591), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n566), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n689), .A3(new_n274), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n273), .B1(new_n566), .B2(new_n593), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n690), .B(KEYINPUT106), .C1(new_n689), .C2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n688), .A2(new_n693), .A3(new_n689), .A4(new_n274), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n312), .A2(new_n343), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n547), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n647), .A2(new_n649), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n273), .A2(new_n698), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n547), .A2(new_n209), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n706), .A2(new_n703), .A3(new_n707), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n702), .A2(new_n708), .A3(new_n709), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n700), .B2(new_n560), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n695), .A2(KEYINPUT107), .A3(new_n555), .A4(new_n699), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(G36gat), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n704), .A2(new_n205), .A3(new_n555), .A4(new_n705), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT46), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(new_n700), .ZN(new_n718));
  INV_X1    g517(.A(new_n569), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n216), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n435), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(G43gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n704), .A2(new_n705), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT47), .ZN(new_n724));
  INV_X1    g523(.A(new_n723), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n695), .A2(new_n674), .A3(new_n699), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(G43gat), .ZN(new_n727));
  OAI22_X1  g526(.A1(new_n720), .A2(new_n724), .B1(new_n727), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n213), .A2(new_n215), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n486), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n704), .A2(new_n705), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n729), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n692), .A2(new_n485), .A3(new_n694), .A4(new_n699), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n731), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n736), .B(new_n738), .C1(new_n735), .C2(new_n734), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n737), .A2(KEYINPUT108), .A3(new_n731), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT108), .B1(new_n737), .B2(new_n731), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n740), .A2(new_n741), .A3(new_n734), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g542(.A1(new_n697), .A2(new_n688), .A3(new_n313), .A4(new_n342), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n547), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n555), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n674), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n721), .A2(G71gat), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n751), .A2(G71gat), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n485), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g555(.A1(new_n697), .A2(new_n312), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n343), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n695), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n701), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n688), .A2(new_n697), .A3(new_n312), .A4(new_n274), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n343), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n764), .B2(new_n763), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n547), .A2(new_n242), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  NOR2_X1   g567(.A1(new_n560), .A2(G92gat), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n761), .A2(new_n762), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n761), .A2(new_n762), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n342), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n692), .A2(new_n555), .A3(new_n694), .A4(new_n758), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n763), .A2(new_n776), .A3(new_n342), .A4(new_n769), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT52), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n775), .A2(new_n772), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n759), .B2(new_n675), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n435), .A2(new_n232), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n766), .B2(new_n784), .ZN(G1338gat));
  NAND4_X1  g584(.A1(new_n763), .A2(new_n233), .A3(new_n485), .A4(new_n342), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n692), .A2(new_n485), .A3(new_n694), .A4(new_n758), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G106gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g589(.A1(new_n313), .A2(new_n697), .A3(new_n343), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n321), .A2(new_n339), .A3(new_n322), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n328), .A2(KEYINPUT54), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n338), .B2(new_n340), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n334), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n793), .A2(new_n795), .A3(KEYINPUT55), .A4(new_n334), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n336), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n599), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n605), .B1(new_n614), .B2(new_n604), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n624), .A2(new_n625), .A3(new_n621), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n642), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n800), .A2(new_n273), .A3(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n342), .B(new_n804), .C1(new_n634), .C2(new_n635), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n642), .A2(KEYINPUT113), .A3(new_n342), .A4(new_n804), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n809), .B(new_n810), .C1(new_n697), .C2(new_n800), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n806), .B1(new_n811), .B2(new_n273), .ZN(new_n812));
  INV_X1    g611(.A(new_n312), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n791), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n547), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n487), .A2(new_n555), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n696), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n814), .A2(new_n557), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n701), .A2(new_n555), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n645), .A2(G113gat), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(G1340gat));
  AOI21_X1  g623(.A(G120gat), .B1(new_n818), .B2(new_n342), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n342), .A2(G120gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n822), .B2(new_n826), .ZN(G1341gat));
  NAND3_X1  g626(.A1(new_n822), .A2(G127gat), .A3(new_n813), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n830));
  AOI21_X1  g629(.A(G127gat), .B1(new_n818), .B2(new_n813), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(G1342gat));
  OR3_X1    g631(.A1(new_n817), .A2(G134gat), .A3(new_n273), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n822), .A2(new_n274), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G134gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(G1343gat));
  NOR3_X1   g637(.A1(new_n674), .A2(new_n486), .A3(new_n555), .ZN(new_n839));
  INV_X1    g638(.A(G141gat), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n645), .A4(new_n815), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n569), .A2(new_n821), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n486), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n807), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n642), .A2(KEYINPUT115), .A3(new_n342), .A4(new_n804), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n798), .A2(new_n336), .A3(new_n799), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n637), .B2(new_n643), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n854), .A3(KEYINPUT116), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT89), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n696), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n800), .B1(new_n858), .B2(new_n636), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n850), .A2(new_n851), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n855), .A2(new_n861), .A3(new_n273), .ZN(new_n862));
  INV_X1    g661(.A(new_n806), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n312), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n848), .B1(new_n865), .B2(new_n791), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n814), .B2(new_n485), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n645), .B(new_n845), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n840), .B1(new_n868), .B2(KEYINPUT117), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n813), .B1(new_n862), .B2(new_n863), .ZN(new_n870));
  INV_X1    g669(.A(new_n791), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n847), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n814), .A2(new_n485), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n846), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n644), .B(new_n844), .C1(new_n872), .C2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n843), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n845), .B1(new_n866), .B2(new_n867), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n697), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n842), .B1(new_n880), .B2(new_n841), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT118), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n843), .ZN(new_n883));
  OAI21_X1  g682(.A(G141gat), .B1(new_n875), .B2(new_n876), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n868), .A2(KEYINPUT117), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n844), .B1(new_n872), .B2(new_n874), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n840), .B1(new_n888), .B2(new_n696), .ZN(new_n889));
  INV_X1    g688(.A(new_n841), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT58), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n882), .A2(new_n892), .ZN(G1344gat));
  NAND2_X1  g692(.A1(new_n839), .A2(new_n815), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n894), .A2(G148gat), .A3(new_n343), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n657), .A2(new_n644), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT119), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n846), .B(new_n485), .C1(new_n898), .C2(new_n870), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n342), .A3(new_n845), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n896), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n896), .A2(G148gat), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n904), .B1(new_n888), .B2(new_n342), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n895), .B1(new_n903), .B2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n879), .B2(new_n312), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n894), .A2(G155gat), .A3(new_n312), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1346gat));
  NAND3_X1  g708(.A1(new_n839), .A2(new_n274), .A3(new_n815), .ZN(new_n910));
  INV_X1    g709(.A(G162gat), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n273), .A2(new_n911), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n910), .A2(new_n911), .B1(new_n888), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT120), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n547), .A2(new_n560), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n820), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(G169gat), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n916), .A2(new_n917), .A3(new_n644), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n814), .A2(new_n701), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(new_n557), .A3(new_n555), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n696), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n918), .B1(new_n917), .B2(new_n921), .ZN(G1348gat));
  INV_X1    g721(.A(G176gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n923), .A3(new_n342), .ZN(new_n924));
  OAI21_X1  g723(.A(G176gat), .B1(new_n916), .B2(new_n343), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  NAND3_X1  g725(.A1(new_n920), .A2(new_n374), .A3(new_n813), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n346), .B1(new_n916), .B2(new_n312), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n920), .A2(new_n349), .A3(new_n274), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n820), .A2(new_n274), .A3(new_n915), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  AND4_X1   g732(.A1(KEYINPUT121), .A2(new_n932), .A3(new_n933), .A4(G190gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n349), .B1(new_n935), .B2(KEYINPUT61), .ZN(new_n936));
  AOI22_X1  g735(.A1(new_n932), .A2(new_n936), .B1(KEYINPUT121), .B2(new_n933), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n931), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT122), .ZN(G1351gat));
  NAND2_X1  g738(.A1(new_n675), .A2(new_n915), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT124), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n901), .A2(new_n645), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G197gat), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n919), .A2(new_n675), .A3(new_n485), .A4(new_n555), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(G197gat), .A3(new_n697), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT123), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n946), .ZN(G1352gat));
  NAND3_X1  g746(.A1(new_n901), .A2(new_n342), .A3(new_n941), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G204gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n944), .A2(G204gat), .A3(new_n343), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n901), .A2(new_n813), .A3(new_n941), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n438), .B1(KEYINPUT125), .B2(new_n954), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n955), .B1(new_n953), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n813), .A2(new_n438), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n957), .A2(new_n958), .B1(new_n944), .B2(new_n959), .ZN(G1354gat));
  NAND2_X1  g759(.A1(new_n274), .A2(G218gat), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n901), .A2(new_n941), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n439), .B1(new_n944), .B2(new_n273), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


