//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G107), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(G101), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT83), .B1(new_n189), .B2(G104), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n189), .A3(G104), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n187), .A3(G107), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n192), .A2(new_n193), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n191), .B1(new_n198), .B2(G101), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(KEYINPUT69), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(KEYINPUT69), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n207), .B(G128), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  INV_X1    g026(.A(new_n203), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n199), .A2(new_n206), .A3(new_n211), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n211), .A2(new_n206), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n199), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT12), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  OAI211_X1 g034(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n220), .C2(G137), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(G134), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n220), .B2(G137), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n220), .A2(KEYINPUT66), .A3(G137), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n225), .A2(new_n228), .A3(new_n232), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n218), .A2(new_n219), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n219), .B1(new_n218), .B2(new_n234), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n193), .A2(new_n197), .ZN(new_n239));
  INV_X1    g053(.A(G101), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n192), .A4(new_n195), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n198), .A2(G101), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n207), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n207), .A2(KEYINPUT0), .A3(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n205), .A2(KEYINPUT0), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT0), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G128), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n204), .A2(new_n251), .A3(KEYINPUT64), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n246), .A2(new_n247), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n198), .A2(new_n254), .A3(G101), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n243), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT10), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n217), .B2(new_n199), .ZN(new_n258));
  INV_X1    g072(.A(new_n234), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n214), .A2(new_n211), .A3(new_n206), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n260), .A2(KEYINPUT10), .A3(new_n241), .A4(new_n191), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n256), .A2(new_n258), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G110), .B(G140), .ZN(new_n263));
  INV_X1    g077(.A(G227), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n263), .B(new_n265), .Z(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n238), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n256), .A2(new_n258), .A3(new_n261), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n234), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n262), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n266), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G469), .B1(new_n273), .B2(G902), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n267), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT84), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n218), .A2(new_n234), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT12), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n278), .A2(new_n262), .A3(new_n266), .A4(new_n235), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G469), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT74), .B(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n238), .A2(KEYINPUT84), .A3(new_n262), .A4(new_n266), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n280), .A2(new_n281), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n285), .A2(new_n286), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n274), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G140), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n290), .A2(KEYINPUT77), .A3(G125), .ZN(new_n291));
  XNOR2_X1  g105(.A(G125), .B(G140), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT16), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT78), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n290), .A3(G125), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n290), .A2(G125), .ZN(new_n298));
  INV_X1    g112(.A(G125), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G140), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n300), .A3(new_n293), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n290), .A2(KEYINPUT77), .A3(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT16), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n296), .A2(G146), .A3(new_n297), .A4(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G237), .A2(G953), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(G143), .A3(G214), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(G143), .B1(new_n307), .B2(G214), .ZN(new_n310));
  OAI21_X1  g124(.A(G131), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G237), .ZN(new_n312));
  INV_X1    g126(.A(G953), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G214), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n202), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n232), .A3(new_n308), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT19), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n292), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n200), .B(new_n319), .C1(new_n303), .C2(new_n318), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n306), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(new_n308), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT91), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT18), .B1(new_n322), .B2(KEYINPUT91), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(new_n232), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n292), .A2(new_n200), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n303), .B2(new_n200), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n322), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(G131), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G113), .B(G122), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(new_n187), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT92), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n296), .A2(new_n297), .A3(new_n305), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n200), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT17), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n311), .A2(new_n338), .A3(new_n316), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n322), .A2(KEYINPUT17), .A3(G131), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n306), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n332), .A3(new_n329), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n330), .A2(new_n344), .A3(new_n333), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n335), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G475), .ZN(new_n347));
  INV_X1    g161(.A(G902), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n342), .A2(new_n332), .A3(new_n329), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n332), .B1(new_n342), .B2(new_n329), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT93), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT93), .B(new_n348), .C1(new_n352), .C2(new_n353), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(G475), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G478), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT96), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(KEYINPUT15), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(KEYINPUT15), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT9), .B(G234), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT81), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n367), .A2(new_n368), .A3(G953), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G122), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT94), .B1(new_n371), .B2(G116), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT94), .ZN(new_n373));
  INV_X1    g187(.A(G116), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G122), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n374), .B2(G122), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G107), .ZN(new_n378));
  XNOR2_X1  g192(.A(G128), .B(G143), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(G134), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n374), .A2(G122), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(new_n376), .B2(KEYINPUT14), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT95), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n372), .A2(new_n375), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT95), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n372), .B2(new_n375), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(new_n381), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AOI211_X1 g203(.A(new_n378), .B(new_n380), .C1(new_n389), .C2(G107), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n379), .A2(new_n220), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n379), .A2(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n202), .A2(G128), .ZN(new_n393));
  OAI21_X1  g207(.A(G134), .B1(new_n393), .B2(KEYINPUT13), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n391), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n378), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n377), .A2(G107), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n370), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n389), .A2(G107), .ZN(new_n400));
  INV_X1    g214(.A(new_n380), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n398), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n369), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n365), .B1(new_n405), .B2(new_n283), .ZN(new_n406));
  AOI211_X1 g220(.A(new_n282), .B(new_n364), .C1(new_n399), .C2(new_n404), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n346), .A2(KEYINPUT20), .A3(new_n347), .A4(new_n348), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n351), .A2(new_n358), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n313), .A2(G952), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(G234), .B2(G237), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n313), .B(new_n283), .C1(G234), .C2(G237), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT21), .B(G898), .Z(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT97), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n367), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n348), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G221), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT82), .Z(new_n421));
  OAI21_X1  g235(.A(G214), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G116), .B(G119), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT5), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n374), .A2(KEYINPUT5), .A3(G119), .ZN(new_n428));
  INV_X1    g242(.A(G113), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT2), .B(G113), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n424), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n436), .B(new_n191), .C1(new_n198), .C2(G101), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT89), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n437), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT89), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n432), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n425), .A2(new_n430), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n199), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n438), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(G110), .B(G122), .Z(new_n446));
  XOR2_X1   g260(.A(new_n446), .B(KEYINPUT8), .Z(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n253), .A2(G125), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n260), .A2(new_n299), .ZN(new_n450));
  INV_X1    g264(.A(G224), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT7), .B1(new_n451), .B2(G953), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n452), .B1(new_n449), .B2(new_n450), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n435), .A2(new_n424), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n436), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n243), .A2(new_n460), .A3(new_n255), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n199), .B2(new_n443), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n462), .A2(new_n446), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n448), .A2(new_n455), .A3(KEYINPUT90), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n458), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n462), .A2(KEYINPUT86), .A3(new_n446), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n449), .A2(new_n450), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n451), .A2(G953), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT87), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n469), .B(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n463), .A2(KEYINPUT6), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n468), .B(new_n472), .C1(new_n473), .C2(new_n466), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n474), .A3(new_n348), .ZN(new_n475));
  OAI21_X1  g289(.A(G210), .B1(G237), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n465), .A2(new_n474), .A3(new_n348), .A4(new_n476), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n423), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n289), .A2(new_n417), .A3(new_n421), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT98), .ZN(new_n482));
  INV_X1    g296(.A(new_n421), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n279), .A2(new_n276), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT84), .B1(new_n271), .B2(new_n267), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n279), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n486), .A2(KEYINPUT85), .A3(new_n281), .A4(new_n283), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n285), .A2(new_n286), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n483), .B1(new_n489), .B2(new_n274), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT98), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n480), .A4(new_n417), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n482), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n337), .A2(new_n306), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT76), .ZN(new_n495));
  INV_X1    g309(.A(G119), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(G128), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n497), .A2(KEYINPUT23), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(KEYINPUT23), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n498), .B(new_n499), .C1(G119), .C2(new_n205), .ZN(new_n500));
  XNOR2_X1  g314(.A(G119), .B(G128), .ZN(new_n501));
  XOR2_X1   g315(.A(KEYINPUT24), .B(G110), .Z(new_n502));
  AOI22_X1  g316(.A1(new_n500), .A2(G110), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  OAI22_X1  g318(.A1(new_n500), .A2(G110), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n306), .A2(new_n505), .A3(new_n326), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT79), .B(KEYINPUT22), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(G137), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n313), .A2(G221), .A3(G234), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n504), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n504), .B2(new_n506), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT25), .B1(new_n513), .B2(new_n282), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n368), .B1(new_n283), .B2(G234), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n516), .B(new_n283), .C1(new_n511), .C2(new_n512), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT80), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n514), .A2(KEYINPUT80), .A3(new_n515), .A4(new_n517), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n515), .A2(G902), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n511), .B2(new_n512), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n527));
  NAND2_X1  g341(.A1(new_n307), .A2(G210), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(G101), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n260), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT67), .B1(new_n223), .B2(G134), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n220), .A3(G137), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n223), .A2(G134), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G131), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT68), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT68), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n540), .A3(G131), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n233), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT70), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n539), .A2(KEYINPUT70), .A3(new_n233), .A4(new_n541), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n532), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n234), .A2(new_n253), .ZN(new_n547));
  INV_X1    g361(.A(new_n460), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(KEYINPUT28), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n537), .A2(new_n540), .A3(G131), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n540), .B1(new_n537), .B2(G131), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n233), .A3(new_n260), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n548), .B1(new_n556), .B2(new_n547), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT28), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n531), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n531), .B1(new_n546), .B2(new_n549), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(KEYINPUT72), .B(new_n531), .C1(new_n546), .C2(new_n549), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT70), .B1(new_n555), .B2(new_n233), .ZN(new_n566));
  INV_X1    g380(.A(new_n545), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n260), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(new_n568), .B2(new_n547), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n556), .A2(new_n547), .A3(new_n565), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n460), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n564), .A2(new_n571), .A3(KEYINPUT31), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n559), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G472), .A2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n526), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT73), .ZN(new_n580));
  INV_X1    g394(.A(new_n559), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n564), .A2(KEYINPUT31), .A3(new_n571), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT31), .B1(new_n564), .B2(new_n571), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT32), .A3(new_n577), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n579), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n577), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT73), .A3(new_n526), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT29), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n552), .A2(new_n558), .A3(new_n531), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n569), .A2(new_n570), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n550), .B1(new_n593), .B2(new_n460), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n591), .B(new_n592), .C1(new_n594), .C2(new_n531), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n548), .B1(new_n568), .B2(new_n547), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n596), .A2(new_n550), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n551), .B1(new_n597), .B2(KEYINPUT28), .ZN(new_n598));
  INV_X1    g412(.A(new_n531), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n591), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n282), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n590), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT75), .B1(new_n589), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n605), .B(new_n602), .C1(new_n586), .C2(new_n588), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n493), .B(new_n525), .C1(new_n604), .C2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  AOI21_X1  g422(.A(new_n590), .B1(new_n584), .B2(new_n283), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n587), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n613), .A2(new_n525), .A3(new_n490), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT100), .ZN(new_n615));
  INV_X1    g429(.A(new_n480), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n416), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n390), .A2(new_n398), .A3(new_n370), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n369), .B1(new_n402), .B2(new_n403), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(KEYINPUT102), .B2(new_n404), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n282), .A2(new_n359), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n405), .A2(new_n618), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(KEYINPUT101), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(KEYINPUT101), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n624), .B(new_n625), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(G478), .B1(new_n405), .B2(new_n283), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT103), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n351), .A2(new_n358), .A3(new_n409), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n617), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n615), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n617), .ZN(new_n642));
  INV_X1    g456(.A(new_n408), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n615), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n504), .A2(new_n506), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n522), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n520), .A2(new_n521), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n493), .A2(new_n613), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT37), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G110), .ZN(G12));
  XNOR2_X1  g470(.A(new_n412), .B(KEYINPUT104), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n657), .B1(new_n413), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n644), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n660), .A2(new_n490), .A3(new_n480), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n653), .B(new_n661), .C1(new_n604), .C2(new_n606), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  INV_X1    g477(.A(new_n572), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n599), .B2(new_n597), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n665), .B2(G902), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n589), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT105), .Z(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n653), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n478), .A2(new_n479), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT38), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n659), .B(KEYINPUT39), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n490), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n643), .B(new_n634), .C1(new_n676), .C2(KEYINPUT40), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(KEYINPUT40), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n422), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n202), .ZN(G45));
  NOR3_X1   g495(.A1(new_n633), .A2(new_n635), .A3(new_n659), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n682), .A2(new_n490), .A3(new_n480), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n653), .B(new_n683), .C1(new_n604), .C2(new_n606), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  INV_X1    g499(.A(new_n486), .ZN(new_n686));
  OAI21_X1  g500(.A(G469), .B1(new_n686), .B2(new_n282), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n489), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n420), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n525), .B(new_n690), .C1(new_n604), .C2(new_n606), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n638), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT41), .B(G113), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  INV_X1    g509(.A(new_n645), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n374), .ZN(G18));
  NOR3_X1   g512(.A1(new_n616), .A2(new_n688), .A3(new_n689), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n699), .A2(new_n417), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(new_n653), .C1(new_n604), .C2(new_n606), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  NAND2_X1  g516(.A1(new_n634), .A2(new_n643), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(KEYINPUT106), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(KEYINPUT106), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n416), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n598), .A2(new_n531), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n574), .A2(new_n575), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n578), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n524), .A2(new_n710), .A3(new_n609), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n699), .A2(new_n706), .A3(new_n707), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n371), .ZN(G24));
  NOR2_X1   g529(.A1(new_n609), .A2(new_n710), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n716), .A2(KEYINPUT108), .A3(new_n653), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT108), .B1(new_n716), .B2(new_n653), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n682), .B(new_n699), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n274), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n273), .A2(KEYINPUT109), .A3(new_n348), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n722), .B1(new_n281), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n689), .B1(new_n724), .B2(new_n489), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n671), .A2(new_n423), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n525), .B(new_n727), .C1(new_n604), .C2(new_n606), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n682), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n603), .A2(new_n579), .A3(new_n585), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n732), .A2(new_n525), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n682), .A3(new_n727), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n729), .A2(new_n731), .B1(KEYINPUT42), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NAND2_X1  g550(.A1(new_n589), .A2(new_n603), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n605), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n589), .A2(KEYINPUT75), .A3(new_n603), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n525), .A3(new_n660), .A4(new_n727), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  INV_X1    g556(.A(new_n726), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n633), .A2(new_n634), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT43), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(new_n653), .C1(new_n611), .C2(new_n612), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n743), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n746), .A2(new_n747), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n273), .B(KEYINPUT45), .Z(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(G469), .ZN(new_n754));
  NAND2_X1  g568(.A1(G469), .A2(G902), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT110), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  AOI211_X1 g573(.A(new_n759), .B(KEYINPUT46), .C1(new_n754), .C2(new_n755), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n755), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n489), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n758), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n689), .A3(new_n674), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n752), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n751), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT112), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n223), .ZN(G39));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n758), .A2(new_n760), .ZN(new_n771));
  INV_X1    g585(.A(new_n762), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n770), .B1(new_n773), .B2(new_n420), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n763), .A2(KEYINPUT113), .A3(new_n689), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n769), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n770), .A3(new_n420), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT113), .B1(new_n763), .B2(new_n689), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT47), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n682), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n738), .A2(new_n739), .A3(new_n524), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n780), .A2(new_n743), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n290), .ZN(G42));
  OAI21_X1  g597(.A(new_n668), .B1(KEYINPUT49), .B2(new_n688), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n483), .B1(new_n688), .B2(KEYINPUT49), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n744), .A3(new_n525), .A4(new_n422), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT114), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n784), .A2(new_n672), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n688), .A2(new_n421), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n776), .B2(new_n779), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n745), .A2(new_n657), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n711), .ZN(new_n792));
  OR3_X1    g606(.A1(new_n790), .A2(new_n743), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n672), .A2(new_n422), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n791), .A2(new_n690), .A3(new_n711), .A4(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT50), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n743), .A2(new_n689), .A3(new_n688), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(new_n412), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n668), .A2(new_n525), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n635), .A3(new_n633), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n791), .A2(new_n797), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n717), .A2(new_n718), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n795), .A2(KEYINPUT50), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n801), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n793), .A2(new_n796), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT51), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n793), .A2(new_n806), .A3(new_n809), .A4(new_n796), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n411), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n800), .A2(new_n636), .ZN(new_n812));
  NAND2_X1  g626(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n802), .A2(new_n733), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n814), .B(new_n815), .Z(new_n816));
  NAND3_X1  g630(.A1(new_n791), .A2(new_n699), .A3(new_n711), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n811), .A2(new_n812), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n704), .A2(new_n705), .A3(new_n616), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n653), .A2(new_n659), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n667), .A2(new_n820), .A3(new_n725), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n662), .A2(new_n684), .A3(new_n719), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n823), .A2(new_n824), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n824), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n803), .A2(new_n682), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n727), .ZN(new_n835));
  INV_X1    g649(.A(new_n659), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n490), .A2(new_n408), .A3(new_n635), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n740), .A2(new_n653), .A3(new_n726), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n735), .A2(new_n835), .A3(new_n741), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n614), .A2(new_n645), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n654), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n614), .A2(new_n638), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n607), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n843), .B1(new_n607), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n692), .A2(new_n645), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n712), .B(KEYINPUT107), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n693), .A2(new_n848), .A3(new_n701), .A4(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n839), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n607), .A2(new_n844), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n607), .A2(new_n843), .A3(new_n844), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n841), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n701), .B1(new_n691), .B2(new_n637), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(new_n697), .A3(new_n714), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n740), .A2(new_n525), .A3(new_n727), .A4(new_n731), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n734), .A2(KEYINPUT42), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n859), .A2(new_n741), .A3(new_n838), .A4(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n856), .A2(new_n858), .A3(new_n861), .A4(new_n835), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n819), .B(new_n833), .C1(new_n852), .C2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n825), .B2(new_n826), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n828), .A2(KEYINPUT118), .A3(new_n830), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT53), .B1(new_n869), .B2(new_n862), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n865), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n851), .A2(KEYINPUT53), .A3(new_n827), .A4(new_n831), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n871), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n818), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n788), .B1(new_n880), .B2(new_n881), .ZN(G75));
  OAI21_X1  g696(.A(new_n819), .B1(new_n869), .B2(new_n862), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n283), .B1(new_n883), .B2(new_n872), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n477), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n468), .B1(new_n473), .B2(new_n466), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(new_n472), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n885), .B2(new_n886), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n313), .A2(G952), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  XOR2_X1   g707(.A(new_n755), .B(KEYINPUT57), .Z(new_n894));
  AOI21_X1  g708(.A(new_n873), .B1(new_n883), .B2(new_n872), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n867), .A2(new_n868), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT53), .B1(new_n896), .B2(new_n851), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n859), .A2(new_n741), .A3(new_n838), .A4(new_n860), .ZN(new_n898));
  INV_X1    g712(.A(new_n835), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(KEYINPUT53), .A3(new_n856), .A4(new_n858), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n832), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n897), .A2(new_n902), .A3(KEYINPUT54), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n894), .B1(new_n895), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(KEYINPUT121), .A3(new_n486), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n906));
  INV_X1    g720(.A(new_n894), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT54), .B1(new_n897), .B2(new_n902), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(new_n875), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n906), .B1(new_n909), .B2(new_n686), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n884), .A2(G469), .A3(new_n753), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n905), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n892), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(G54));
  NAND4_X1  g728(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .A4(new_n346), .ZN(new_n915));
  INV_X1    g729(.A(new_n346), .ZN(new_n916));
  OAI211_X1 g730(.A(KEYINPUT58), .B(new_n282), .C1(new_n897), .C2(new_n902), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n347), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT122), .ZN(G60));
  NOR2_X1   g734(.A1(new_n895), .A2(new_n903), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n627), .A2(new_n628), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n621), .B2(new_n623), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n913), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n877), .A2(new_n879), .A3(new_n926), .ZN(new_n929));
  INV_X1    g743(.A(new_n923), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(new_n883), .A2(new_n872), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n368), .A2(new_n348), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n651), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n932), .A2(new_n935), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n513), .B(KEYINPUT124), .Z(new_n938));
  OAI211_X1 g752(.A(new_n913), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G66));
  NAND2_X1  g755(.A1(new_n856), .A2(new_n858), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n313), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n415), .B2(new_n451), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n887), .B1(G898), .B2(new_n313), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT125), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G69));
  OAI21_X1  g762(.A(new_n319), .B1(new_n303), .B2(new_n318), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n593), .B(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n662), .A2(new_n719), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n684), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n782), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n764), .A2(new_n733), .A3(new_n820), .ZN(new_n954));
  AOI22_X1  g768(.A1(new_n751), .A2(new_n765), .B1(KEYINPUT126), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n735), .B1(new_n954), .B2(KEYINPUT126), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n953), .A2(new_n955), .A3(new_n741), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n950), .B1(new_n958), .B2(new_n313), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n264), .A2(G900), .A3(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n264), .A2(new_n658), .A3(new_n313), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n684), .B(new_n951), .C1(new_n679), .C2(new_n673), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n782), .B1(KEYINPUT62), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n740), .A2(new_n525), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n636), .B1(new_n643), .B2(new_n635), .ZN(new_n967));
  OR4_X1    g781(.A1(new_n966), .A2(new_n676), .A3(new_n743), .A4(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n964), .A2(new_n965), .A3(new_n766), .A4(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n950), .B1(new_n969), .B2(G953), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n961), .B1(new_n962), .B2(new_n970), .ZN(G72));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n969), .B2(new_n942), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n594), .A2(new_n599), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n973), .B1(new_n958), .B2(new_n942), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n599), .A3(new_n594), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n976), .A2(new_n913), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n865), .A2(new_n870), .ZN(new_n980));
  INV_X1    g794(.A(new_n973), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n594), .A2(new_n531), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n664), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT127), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n984), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n892), .B1(new_n974), .B2(new_n975), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n986), .A2(new_n987), .A3(new_n978), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n985), .A2(new_n989), .ZN(G57));
endmodule


