//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT79), .ZN(new_n203));
  OR2_X1    g002(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(G155gat), .A3(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT2), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n207), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT76), .B1(new_n210), .B2(G141gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n212));
  INV_X1    g011(.A(G141gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(G148gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(G141gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n208), .A2(new_n209), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n218), .B(KEYINPUT75), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(G148gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT2), .B1(new_n215), .B2(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n222), .A2(new_n217), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n203), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n216), .A2(new_n219), .ZN(new_n227));
  INV_X1    g026(.A(new_n205), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n229));
  INV_X1    g028(.A(G155gat), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT78), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT2), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n227), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  OR3_X1    g034(.A1(new_n222), .A2(new_n217), .A3(new_n224), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239));
  XOR2_X1   g038(.A(G211gat), .B(G218gat), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT71), .ZN(new_n241));
  XNOR2_X1  g040(.A(G197gat), .B(G204gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243));
  INV_X1    g042(.A(G211gat), .ZN(new_n244));
  INV_X1    g043(.A(G218gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n241), .B(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n239), .B1(new_n248), .B2(KEYINPUT29), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n236), .A3(new_n239), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT29), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n202), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n240), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n252), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n256), .A2(new_n240), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n239), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n235), .A2(new_n236), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n260), .A2(new_n261), .B1(G228gat), .B2(G233gat), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(G22gat), .B1(new_n255), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n265));
  INV_X1    g064(.A(G22gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(new_n262), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n238), .A2(new_n249), .B1(new_n253), .B2(new_n248), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n266), .B(new_n267), .C1(new_n268), .C2(new_n202), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G78gat), .B(G106gat), .Z(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n264), .A2(new_n265), .A3(new_n269), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT31), .B(G50gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n272), .A2(new_n276), .A3(new_n274), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT35), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OR3_X1    g084(.A1(new_n285), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(G169gat), .ZN(new_n290));
  INV_X1    g089(.A(G176gat), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT26), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(KEYINPUT26), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n290), .A2(new_n291), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n286), .A2(new_n288), .A3(new_n289), .A4(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n289), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n300), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT65), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n299), .A2(G169gat), .A3(G176gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(new_n294), .ZN(new_n310));
  OAI211_X1 g109(.A(KEYINPUT65), .B(new_n293), .C1(new_n296), .C2(new_n299), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n307), .A2(KEYINPUT66), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  OR2_X1    g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT24), .A3(new_n289), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n316), .A2(KEYINPUT25), .A3(new_n302), .A4(new_n300), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n313), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n293), .B1(new_n296), .B2(new_n299), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n306), .B1(new_n305), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT64), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g122(.A(KEYINPUT64), .B(new_n306), .C1(new_n305), .C2(new_n320), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n298), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327));
  OAI21_X1  g126(.A(G127gat), .B1(new_n327), .B2(KEYINPUT1), .ZN(new_n328));
  INV_X1    g127(.A(G120gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G113gat), .ZN(new_n330));
  INV_X1    g129(.A(G113gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G120gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n328), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G134gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n328), .A2(new_n336), .A3(G134gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G227gat), .A2(G233gat), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n312), .A2(new_n318), .A3(new_n323), .A4(new_n324), .ZN(new_n344));
  INV_X1    g143(.A(new_n340), .ZN(new_n345));
  AOI21_X1  g144(.A(G134gat), .B1(new_n328), .B2(new_n336), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(new_n347), .A3(new_n298), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT34), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT34), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n342), .A2(new_n351), .A3(new_n343), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT68), .B(G15gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(G43gat), .ZN(new_n355));
  XOR2_X1   g154(.A(G71gat), .B(G99gat), .Z(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n343), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n344), .A2(new_n347), .A3(new_n298), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n347), .B1(new_n344), .B2(new_n298), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n362), .B2(KEYINPUT32), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n357), .A2(KEYINPUT33), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(KEYINPUT32), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT69), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n362), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n366), .ZN(new_n370));
  AOI221_X4 g169(.A(new_n353), .B1(new_n363), .B2(new_n365), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n353), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(new_n365), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n371), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n342), .A2(new_n348), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(new_n359), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT69), .B1(new_n380), .B2(new_n366), .ZN(new_n381));
  INV_X1    g180(.A(new_n370), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n374), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n353), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n373), .A2(new_n372), .A3(new_n374), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT86), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n280), .B(new_n282), .C1(new_n377), .C2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT73), .ZN(new_n390));
  INV_X1    g189(.A(G8gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n248), .ZN(new_n393));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI211_X1 g194(.A(KEYINPUT29), .B(new_n395), .C1(new_n344), .C2(new_n298), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n344), .A2(new_n395), .A3(new_n298), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n393), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT72), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n326), .A2(new_n252), .A3(new_n394), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(new_n248), .A3(new_n397), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT72), .B(new_n393), .C1(new_n396), .C2(new_n398), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n392), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n405), .A2(KEYINPUT30), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n404), .ZN(new_n407));
  INV_X1    g206(.A(new_n392), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT74), .ZN(new_n411));
  AND4_X1   g210(.A1(new_n411), .A2(new_n407), .A3(KEYINPUT30), .A4(new_n408), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n405), .B2(KEYINPUT30), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n406), .B(new_n410), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n251), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n238), .B2(KEYINPUT3), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n347), .A2(KEYINPUT80), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n341), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n416), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n235), .A2(new_n339), .A3(new_n236), .A4(new_n340), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(KEYINPUT4), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n221), .A2(new_n225), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n429), .A2(KEYINPUT82), .A3(new_n347), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n423), .A2(new_n424), .A3(new_n425), .A4(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n235), .A2(KEYINPUT79), .A3(new_n236), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT79), .B1(new_n235), .B2(new_n236), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT3), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(new_n422), .A3(new_n251), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n427), .B2(KEYINPUT4), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n429), .A2(KEYINPUT81), .A3(new_n347), .A4(new_n430), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n432), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n442), .A3(new_n415), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n419), .A2(new_n421), .B1(new_n226), .B2(new_n237), .ZN(new_n444));
  INV_X1    g243(.A(new_n427), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n416), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(KEYINPUT5), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n438), .A2(new_n433), .A3(new_n425), .A4(new_n415), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT83), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT0), .B(G57gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(G85gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(G1gat), .B(G29gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(new_n455), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n434), .A2(new_n447), .A3(new_n449), .A4(new_n454), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n414), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n371), .B(new_n375), .C1(new_n278), .C2(new_n279), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n387), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n376), .B1(new_n371), .B2(new_n375), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n384), .A2(KEYINPUT86), .A3(new_n385), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT35), .ZN(new_n468));
  AND4_X1   g267(.A1(new_n281), .A2(new_n467), .A3(new_n468), .A4(new_n280), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n461), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n460), .A2(new_n456), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n408), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT74), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n405), .A2(new_n411), .A3(KEYINPUT30), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n409), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n406), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n280), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n371), .A2(new_n375), .ZN(new_n478));
  AND2_X1   g277(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n476), .A2(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n407), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n407), .A2(new_n484), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT38), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n484), .B1(new_n399), .B2(new_n402), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n489), .A2(KEYINPUT38), .A3(new_n408), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT38), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n403), .A2(new_n491), .A3(new_n404), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n485), .A2(new_n490), .B1(new_n408), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n488), .A2(new_n460), .A3(new_n456), .A4(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n414), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n415), .B1(new_n438), .B2(new_n433), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT39), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n454), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n444), .A2(new_n416), .A3(new_n445), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n496), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT40), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n496), .B(new_n505), .C1(new_n500), .C2(new_n502), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n457), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n280), .B(new_n494), .C1(new_n495), .C2(new_n507), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n464), .A2(new_n470), .B1(new_n483), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  INV_X1    g315(.A(G36gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n513), .A2(G36gat), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n519), .B(new_n521), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n518), .A2(new_n514), .ZN(new_n526));
  OR2_X1    g325(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(G36gat), .A3(new_n510), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n526), .B(new_n528), .C1(KEYINPUT15), .C2(new_n520), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n528), .A3(new_n524), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n522), .A3(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n525), .A2(new_n531), .A3(KEYINPUT17), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT17), .B1(new_n525), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(G15gat), .A2(G22gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(G15gat), .A2(G22gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT91), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G15gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n266), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  NAND2_X1  g339(.A1(G15gat), .A2(G22gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT16), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G1gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT92), .B1(new_n537), .B2(new_n542), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(G1gat), .ZN(new_n551));
  OAI21_X1  g350(.A(G8gat), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n550), .A2(G1gat), .B1(new_n543), .B2(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n548), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n391), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT93), .B1(new_n534), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n555), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n391), .B1(new_n553), .B2(new_n554), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n525), .A2(new_n531), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n525), .A2(new_n531), .A3(KEYINPUT17), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n556), .A2(new_n525), .A3(new_n531), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT94), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n557), .A2(new_n567), .A3(new_n568), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT95), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT18), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n560), .A2(new_n562), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n568), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n570), .B(KEYINPUT13), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT18), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n572), .A2(KEYINPUT95), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G169gat), .B(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT12), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n574), .A2(new_n578), .A3(new_n580), .A4(new_n587), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT96), .B1(new_n509), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n593));
  INV_X1    g392(.A(new_n591), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT35), .A2(new_n463), .B1(new_n469), .B2(new_n461), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n476), .A2(new_n477), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n480), .A2(new_n482), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n508), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  INV_X1    g401(.A(G57gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(G64gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT97), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n608), .A3(KEYINPUT9), .ZN(new_n609));
  XOR2_X1   g408(.A(G71gat), .B(G78gat), .Z(new_n610));
  INV_X1    g409(.A(G71gat), .ZN(new_n611));
  INV_X1    g410(.A(G78gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT9), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n609), .A2(new_n610), .B1(new_n614), .B2(new_n605), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n620));
  OR3_X1    g419(.A1(new_n556), .A2(KEYINPUT98), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT98), .B1(new_n556), .B2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G127gat), .B(G155gat), .Z(new_n624));
  OR2_X1    g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n624), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(new_n625), .B2(new_n630), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n619), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n618), .A3(new_n631), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  INV_X1    g438(.A(G85gat), .ZN(new_n640));
  INV_X1    g439(.A(G92gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(KEYINPUT8), .A2(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT7), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n640), .B2(new_n641), .ZN(new_n644));
  NAND3_X1  g443(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G99gat), .B(G106gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n566), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n646), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n525), .A3(new_n531), .ZN(new_n652));
  NAND3_X1  g451(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n652), .A2(KEYINPUT99), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT99), .B1(new_n652), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n649), .B(new_n659), .C1(new_n654), .C2(new_n655), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n638), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(new_n638), .A3(new_n660), .ZN(new_n663));
  XNOR2_X1  g462(.A(G134gat), .B(G162gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G190gat), .B(G218gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  AND3_X1   g465(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n662), .B2(new_n663), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n637), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT103), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n329), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n609), .A2(new_n610), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n614), .A2(new_n605), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n646), .B2(new_n647), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n648), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n651), .A2(new_n615), .A3(new_n681), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT10), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n651), .A2(new_n615), .A3(KEYINPUT10), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(G230gat), .A2(G233gat), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n683), .B2(new_n684), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n677), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(KEYINPUT104), .B(new_n677), .C1(new_n691), .C2(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n686), .A2(new_n698), .A3(new_n687), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n686), .B2(new_n687), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n689), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n692), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n676), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n672), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n600), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n471), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G1gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n706), .A2(new_n548), .A3(new_n707), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1324gat));
  NOR2_X1   g510(.A1(new_n544), .A2(new_n391), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n706), .A2(KEYINPUT42), .A3(new_n414), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n600), .A2(new_n414), .A3(new_n705), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(new_n712), .A3(new_n713), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n716), .B2(G8gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(G1325gat));
  AOI21_X1  g519(.A(G15gat), .B1(new_n706), .B2(new_n467), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n597), .A2(new_n538), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT105), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n706), .B2(new_n723), .ZN(G1326gat));
  XNOR2_X1  g523(.A(KEYINPUT43), .B(G22gat), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n706), .A2(new_n477), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n706), .B2(new_n477), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(G1327gat));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n509), .B2(new_n669), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT44), .B(new_n670), .C1(new_n595), .C2(new_n598), .ZN(new_n731));
  INV_X1    g530(.A(new_n637), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n704), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n591), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n730), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n513), .B1(new_n736), .B2(new_n471), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n734), .B1(new_n592), .B2(new_n599), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n670), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n471), .A2(new_n513), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND4_X1   g541(.A1(new_n738), .A2(new_n739), .A3(new_n670), .A4(new_n741), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(G1328gat));
  NAND4_X1  g543(.A1(new_n739), .A2(new_n517), .A3(new_n414), .A4(new_n670), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n746));
  OAI21_X1  g545(.A(G36gat), .B1(new_n736), .B2(new_n495), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(G1329gat));
  OAI21_X1  g548(.A(G43gat), .B1(new_n736), .B2(new_n597), .ZN(new_n750));
  INV_X1    g549(.A(new_n467), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n739), .A2(new_n670), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n753), .A3(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1330gat));
  NAND4_X1  g557(.A1(new_n730), .A2(new_n477), .A3(new_n731), .A4(new_n735), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G50gat), .ZN(new_n760));
  INV_X1    g559(.A(G50gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n600), .A2(new_n761), .A3(new_n670), .A4(new_n733), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n762), .B2(new_n280), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(KEYINPUT48), .B(new_n760), .C1(new_n762), .C2(new_n280), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1331gat));
  NAND2_X1  g566(.A1(new_n483), .A2(new_n508), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n465), .A2(new_n466), .B1(new_n278), .B2(new_n279), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n476), .B1(new_n769), .B2(new_n282), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n468), .B1(new_n770), .B2(new_n462), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n387), .A2(KEYINPUT87), .A3(new_n476), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n704), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n594), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(new_n671), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n471), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n603), .ZN(G1332gat));
  AOI21_X1  g577(.A(new_n495), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT106), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n776), .A2(KEYINPUT107), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT107), .B1(new_n776), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1333gat));
  OAI21_X1  g584(.A(new_n611), .B1(new_n776), .B2(new_n751), .ZN(new_n786));
  AND4_X1   g585(.A1(G71gat), .A2(new_n773), .A3(new_n671), .A4(new_n775), .ZN(new_n787));
  INV_X1    g586(.A(new_n597), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT108), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n790));
  NOR4_X1   g589(.A1(new_n776), .A2(new_n790), .A3(new_n611), .A4(new_n597), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n793), .B(new_n786), .C1(new_n789), .C2(new_n791), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1334gat));
  NOR2_X1   g596(.A1(new_n776), .A2(new_n280), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(new_n612), .ZN(G1335gat));
  NOR2_X1   g598(.A1(new_n732), .A2(new_n594), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n730), .A2(new_n704), .A3(new_n731), .A4(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801), .B2(new_n471), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n670), .B(new_n800), .C1(new_n595), .C2(new_n598), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n773), .A2(KEYINPUT51), .A3(new_n670), .A4(new_n800), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n707), .A2(new_n640), .A3(new_n704), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT110), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT111), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n802), .A2(new_n813), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1336gat));
  OAI21_X1  g614(.A(G92gat), .B1(new_n801), .B2(new_n495), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n414), .A2(new_n641), .A3(new_n704), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT112), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n819), .B1(new_n807), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n818), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n816), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n816), .B2(new_n822), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(G1337gat));
  OAI21_X1  g625(.A(G99gat), .B1(new_n801), .B2(new_n597), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n751), .A2(G99gat), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n807), .A2(new_n704), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1338gat));
  OAI21_X1  g629(.A(G106gat), .B1(new_n801), .B2(new_n280), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n280), .A2(G106gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n807), .A2(new_n704), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1339gat));
  INV_X1    g637(.A(new_n769), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n557), .A2(new_n567), .A3(new_n568), .ZN(new_n840));
  OAI22_X1  g639(.A1(new_n840), .A2(new_n571), .B1(new_n576), .B2(new_n577), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n586), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n590), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT114), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n688), .A2(new_n690), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n701), .A2(KEYINPUT54), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n676), .B1(new_n691), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(KEYINPUT55), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT55), .B1(new_n846), .B2(new_n848), .ZN(new_n851));
  INV_X1    g650(.A(new_n703), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n590), .A2(new_n854), .A3(new_n842), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n844), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n670), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n704), .A2(new_n590), .A3(new_n842), .ZN(new_n858));
  INV_X1    g657(.A(new_n851), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n703), .A3(new_n849), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n669), .B(new_n858), .C1(new_n591), .C2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n861), .A3(new_n637), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n671), .A2(new_n591), .A3(new_n774), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT115), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n862), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n839), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n471), .A2(new_n414), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n591), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n865), .A2(new_n867), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n462), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n331), .A3(new_n869), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n874), .B2(new_n591), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1340gat));
  OAI21_X1  g676(.A(G120gat), .B1(new_n870), .B2(new_n774), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n869), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n704), .A2(new_n329), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(G1341gat));
  NOR3_X1   g680(.A1(new_n870), .A2(new_n335), .A3(new_n637), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n873), .A2(new_n732), .A3(new_n869), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n335), .B2(new_n883), .ZN(G1342gat));
  NAND2_X1  g683(.A1(new_n495), .A2(new_n670), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT117), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n873), .A2(new_n338), .A3(new_n707), .A4(new_n886), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT56), .ZN(new_n888));
  OAI21_X1  g687(.A(G134gat), .B1(new_n870), .B2(new_n669), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(KEYINPUT56), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(G1343gat));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n872), .A2(new_n892), .A3(new_n477), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n597), .A2(new_n869), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n864), .A2(new_n477), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(KEYINPUT57), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n594), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G141gat), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n471), .B1(new_n865), .B2(new_n867), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n280), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n862), .A2(new_n863), .A3(new_n866), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n866), .B1(new_n862), .B2(new_n863), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n707), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n788), .B1(new_n904), .B2(KEYINPUT118), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n901), .A2(new_n905), .A3(new_n213), .A4(new_n495), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n898), .B1(new_n906), .B2(new_n591), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT58), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n909), .B(new_n898), .C1(new_n906), .C2(new_n591), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n896), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT59), .B(new_n210), .C1(new_n913), .C2(new_n704), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT57), .B(new_n477), .C1(new_n902), .C2(new_n903), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT119), .B1(new_n895), .B2(new_n892), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n872), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n477), .ZN(new_n919));
  INV_X1    g718(.A(new_n894), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n704), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n921), .B2(G148gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n901), .A2(new_n905), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n495), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n704), .A2(new_n210), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n914), .A2(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G1345gat));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n495), .A3(new_n732), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n732), .A2(G155gat), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT120), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n928), .A2(new_n230), .B1(new_n913), .B2(new_n930), .ZN(G1346gat));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n204), .A2(new_n205), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n913), .B2(new_n670), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n886), .A2(new_n933), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n923), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n912), .A2(new_n669), .ZN(new_n938));
  OAI221_X1 g737(.A(KEYINPUT121), .B1(new_n923), .B2(new_n935), .C1(new_n938), .C2(new_n933), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n707), .A2(new_n495), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n873), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n290), .A3(new_n594), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n872), .A2(new_n769), .A3(new_n941), .ZN(new_n945));
  OAI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n591), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1348gat));
  NOR3_X1   g746(.A1(new_n945), .A2(new_n291), .A3(new_n774), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n291), .B1(new_n942), .B2(new_n774), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g750(.A(KEYINPUT122), .B(new_n291), .C1(new_n942), .C2(new_n774), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G1349gat));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n954), .B1(new_n945), .B2(new_n637), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n868), .A2(KEYINPUT123), .A3(new_n732), .A4(new_n941), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(G183gat), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n873), .A2(new_n283), .A3(new_n732), .A4(new_n941), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT60), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n284), .A3(new_n670), .ZN(new_n964));
  INV_X1    g763(.A(new_n945), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n284), .B1(new_n965), .B2(new_n670), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n966), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  AND2_X1   g770(.A1(new_n918), .A2(new_n919), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n597), .A2(new_n941), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(G197gat), .B1(new_n975), .B2(new_n591), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n872), .A2(new_n477), .A3(new_n974), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  INV_X1    g777(.A(G197gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n280), .B1(new_n865), .B2(new_n867), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n980), .A2(new_n981), .A3(new_n974), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n978), .A2(new_n979), .A3(new_n594), .A4(new_n982), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n983), .A2(KEYINPUT125), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(KEYINPUT125), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n976), .B1(new_n984), .B2(new_n985), .ZN(G1352gat));
  NAND3_X1  g785(.A1(new_n972), .A2(new_n704), .A3(new_n974), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(G204gat), .ZN(new_n988));
  AOI21_X1  g787(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n980), .A2(new_n704), .A3(new_n974), .A4(new_n989), .ZN(new_n990));
  NOR2_X1   g789(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n988), .A2(new_n992), .ZN(G1353gat));
  AND2_X1   g792(.A1(new_n978), .A2(new_n982), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n994), .A2(new_n244), .A3(new_n732), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n918), .A2(new_n919), .A3(new_n732), .A4(new_n974), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n975), .B2(new_n669), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n994), .A2(new_n245), .A3(new_n670), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


