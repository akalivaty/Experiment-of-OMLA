//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT80), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G107), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n190), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n189), .A2(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n188), .B(G101), .C1(new_n194), .C2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n191), .B1(new_n193), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(new_n195), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .A4(new_n190), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n202), .A3(new_n190), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n188), .B1(new_n206), .B2(G101), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n187), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n204), .A2(KEYINPUT4), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n194), .B2(new_n198), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT80), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT81), .A4(new_n199), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT2), .A2(G113), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n216));
  INV_X1    g030(.A(G113), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n214), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G116), .ZN(new_n222));
  INV_X1    g036(.A(G116), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G119), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n220), .B(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n206), .A2(new_n227), .A3(G101), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n213), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G110), .B(G122), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT5), .ZN(new_n233));
  OAI21_X1  g047(.A(G113), .B1(new_n222), .B2(KEYINPUT5), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT86), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n220), .A2(new_n225), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n223), .A2(G119), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT5), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n217), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT86), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT5), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n236), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n193), .A2(new_n190), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n204), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT87), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n204), .A2(new_n245), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT87), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n239), .A2(new_n241), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n250), .A2(KEYINPUT86), .B1(new_n220), .B2(new_n225), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .A4(new_n242), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n231), .A2(new_n232), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n232), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n229), .B1(new_n208), .B2(new_n212), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n247), .A2(new_n252), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n258), .A3(KEYINPUT6), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(G146), .ZN(new_n263));
  INV_X1    g077(.A(G146), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT65), .A3(G143), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G143), .B(G146), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT0), .B(G128), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT64), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n263), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n268), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G125), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n261), .A2(G146), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n281));
  OAI21_X1  g095(.A(G128), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n274), .ZN(new_n283));
  INV_X1    g097(.A(G125), .ZN(new_n284));
  INV_X1    g098(.A(G128), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT1), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n262), .A2(new_n265), .A3(new_n286), .A4(new_n263), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G224), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(G953), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n289), .B(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n293), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n259), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT90), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n251), .A2(new_n246), .A3(new_n242), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n232), .B(KEYINPUT8), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n220), .A2(new_n225), .B1(new_n239), .B2(new_n241), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n204), .B(new_n245), .C1(new_n299), .C2(KEYINPUT88), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n299), .A2(KEYINPUT88), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n297), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT7), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n291), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT64), .B1(new_n269), .B2(new_n270), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n274), .A2(new_n276), .A3(new_n272), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n305), .A2(new_n306), .B1(new_n266), .B2(new_n267), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n288), .B(new_n304), .C1(new_n307), .C2(new_n284), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n279), .A2(KEYINPUT89), .A3(new_n288), .A4(new_n304), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n306), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n284), .B1(new_n312), .B2(new_n268), .ZN(new_n313));
  INV_X1    g127(.A(new_n288), .ZN(new_n314));
  OAI22_X1  g128(.A1(new_n313), .A2(new_n314), .B1(new_n303), .B2(new_n291), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n302), .A2(new_n310), .A3(new_n311), .A4(new_n315), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n213), .A2(new_n230), .B1(new_n252), .B2(new_n247), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n232), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n296), .B1(new_n318), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(G902), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n256), .A2(new_n257), .A3(new_n255), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT90), .B(new_n320), .C1(new_n321), .C2(new_n316), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n295), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G210), .B1(G237), .B2(G902), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT91), .Z(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n295), .A2(new_n319), .A3(new_n322), .A4(new_n324), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT20), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n331), .A2(KEYINPUT76), .A3(G125), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n284), .A2(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(G125), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT76), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n330), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n331), .A3(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT77), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n340), .A2(new_n330), .A3(new_n331), .A4(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n264), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n339), .A2(new_n341), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n332), .B1(new_n345), .B2(KEYINPUT76), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n344), .B(G146), .C1(new_n330), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n348));
  INV_X1    g162(.A(G237), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(G214), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n261), .ZN(new_n352));
  NOR2_X1   g166(.A1(G237), .A2(G953), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(G143), .A3(G214), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n348), .A2(new_n355), .A3(KEYINPUT17), .A4(G131), .ZN(new_n356));
  INV_X1    g170(.A(G131), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n352), .B2(new_n354), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n348), .B1(new_n358), .B2(KEYINPUT17), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n343), .B(new_n347), .C1(new_n356), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT94), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n355), .A2(KEYINPUT17), .A3(G131), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT93), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n348), .A3(KEYINPUT17), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n343), .A4(new_n347), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n355), .A2(G131), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n358), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n361), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G113), .B(G122), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n189), .ZN(new_n374));
  NAND2_X1  g188(.A1(KEYINPUT18), .A2(G131), .ZN(new_n375));
  OR3_X1    g189(.A1(new_n355), .A2(KEYINPUT92), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n355), .B2(KEYINPUT92), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n346), .A2(G146), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n345), .A2(new_n264), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n372), .A2(new_n374), .A3(new_n382), .ZN(new_n383));
  MUX2_X1   g197(.A(new_n345), .B(new_n346), .S(KEYINPUT19), .Z(new_n384));
  OAI221_X1 g198(.A(new_n347), .B1(new_n358), .B2(new_n368), .C1(new_n384), .C2(G146), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n374), .B1(new_n385), .B2(new_n382), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(G475), .A2(G902), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n329), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT20), .B(new_n391), .C1(new_n383), .C2(new_n387), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n372), .A2(new_n382), .ZN(new_n393));
  INV_X1    g207(.A(new_n374), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(G902), .B1(new_n395), .B2(new_n383), .ZN(new_n396));
  INV_X1    g210(.A(G475), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n390), .A2(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT9), .B(G234), .ZN(new_n399));
  INV_X1    g213(.A(G217), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n399), .A2(new_n400), .A3(G953), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT95), .ZN(new_n403));
  INV_X1    g217(.A(G122), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(G116), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n223), .A2(KEYINPUT95), .A3(G122), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n223), .A2(G122), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n192), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT97), .ZN(new_n411));
  XNOR2_X1  g225(.A(G128), .B(G143), .ZN(new_n412));
  INV_X1    g226(.A(G134), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n407), .A2(new_n415), .A3(new_n192), .A4(new_n409), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n223), .A2(KEYINPUT95), .A3(G122), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT95), .B1(new_n223), .B2(G122), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT98), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n421), .A3(new_n409), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n405), .B2(new_n406), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT98), .B1(new_n424), .B2(new_n408), .ZN(new_n425));
  INV_X1    g239(.A(new_n407), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n423), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n422), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n417), .B1(G107), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n285), .A2(G143), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(G134), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n261), .A2(G128), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n431), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n413), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n412), .A2(G134), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n430), .A2(G134), .A3(new_n433), .A4(new_n431), .ZN(new_n438));
  INV_X1    g252(.A(new_n410), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n192), .B1(new_n407), .B2(new_n409), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n402), .B1(new_n429), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n420), .A2(new_n409), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n444), .A2(KEYINPUT98), .B1(new_n423), .B2(new_n426), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n192), .B1(new_n445), .B2(new_n422), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n441), .B(new_n401), .C1(new_n446), .C2(new_n417), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT99), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT99), .B(new_n402), .C1(new_n429), .C2(new_n442), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n320), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT100), .ZN(new_n452));
  INV_X1    g266(.A(G478), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(KEYINPUT15), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT100), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n449), .A2(new_n455), .A3(new_n320), .A4(new_n450), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n451), .A2(new_n454), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n398), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G952), .ZN(new_n461));
  AOI211_X1 g275(.A(G953), .B(new_n461), .C1(G234), .C2(G237), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n320), .B(new_n350), .C1(G234), .C2(G237), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(G898), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT85), .Z(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n328), .A2(new_n460), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G469), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n413), .A2(G137), .ZN(new_n472));
  AND2_X1   g286(.A1(KEYINPUT67), .A2(G137), .ZN(new_n473));
  NOR2_X1   g287(.A1(KEYINPUT67), .A2(G137), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT11), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n413), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n472), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n413), .B2(G137), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(KEYINPUT66), .B(new_n476), .C1(new_n413), .C2(G137), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n478), .A2(new_n483), .A3(new_n357), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n357), .B1(new_n478), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n307), .A2(new_n228), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n208), .B2(new_n212), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n283), .A2(new_n287), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n248), .A2(KEYINPUT10), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n282), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n494), .A2(new_n287), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n492), .B1(new_n495), .B2(new_n246), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n487), .B1(new_n489), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G110), .B(G140), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n350), .A2(G227), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT83), .ZN(new_n503));
  INV_X1    g317(.A(new_n488), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n497), .B1(new_n213), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n503), .B1(new_n505), .B2(new_n486), .ZN(new_n506));
  NOR4_X1   g320(.A1(new_n489), .A2(KEYINPUT83), .A3(new_n497), .A4(new_n487), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n498), .B(new_n502), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n248), .A2(new_n490), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n495), .A2(new_n246), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n487), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT12), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n213), .A2(new_n504), .ZN(new_n513));
  INV_X1    g327(.A(new_n497), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n486), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT83), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n505), .A2(new_n503), .A3(new_n486), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n508), .B1(new_n518), .B2(new_n502), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n471), .B1(new_n519), .B2(new_n320), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n512), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT84), .B(new_n502), .C1(new_n506), .C2(new_n507), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n501), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n520), .B1(new_n529), .B2(new_n471), .ZN(new_n530));
  OAI21_X1  g344(.A(G221), .B1(new_n399), .B2(G902), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n470), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n347), .A2(new_n343), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT23), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n221), .B2(G128), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n285), .A2(KEYINPUT23), .A3(G119), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n537), .C1(G119), .C2(new_n285), .ZN(new_n538));
  XNOR2_X1  g352(.A(G119), .B(G128), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT24), .B(G110), .Z(new_n540));
  AOI22_X1  g354(.A1(new_n538), .A2(G110), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n538), .A2(G110), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n347), .A2(new_n380), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT22), .B(G137), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n545), .B(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n320), .C1(KEYINPUT78), .C2(KEYINPUT25), .ZN(new_n550));
  AND2_X1   g364(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G234), .ZN(new_n553));
  OAI21_X1  g367(.A(G217), .B1(new_n553), .B2(G902), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n550), .B2(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n320), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n549), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G472), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n307), .B1(new_n484), .B2(new_n485), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n478), .A2(new_n483), .A3(new_n357), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n475), .A2(G134), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n413), .A2(G137), .ZN(new_n565));
  OAI21_X1  g379(.A(G131), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n566), .A3(new_n490), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT74), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(new_n226), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(KEYINPUT74), .A3(new_n567), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT28), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n226), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n562), .B2(new_n567), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n562), .A2(new_n572), .A3(new_n567), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n571), .B1(KEYINPUT28), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n353), .A2(G210), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT27), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT26), .B(G101), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT29), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n577), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n562), .A2(new_n567), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT68), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT30), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n562), .A2(new_n587), .A3(new_n588), .A4(new_n567), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n572), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n575), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n582), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n596), .B2(new_n573), .ZN(new_n599));
  INV_X1    g413(.A(new_n570), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n600), .A2(new_n568), .A3(new_n226), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n601), .B2(KEYINPUT28), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n597), .B(new_n583), .C1(new_n602), .C2(new_n582), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n561), .B1(new_n585), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n575), .A2(new_n581), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT70), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n575), .A2(KEYINPUT70), .A3(new_n581), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n610));
  AOI211_X1 g424(.A(new_n589), .B(new_n591), .C1(new_n562), .C2(new_n567), .ZN(new_n611));
  INV_X1    g425(.A(new_n594), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n226), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT72), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n609), .A2(new_n613), .A3(KEYINPUT72), .A4(new_n610), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n609), .A2(new_n613), .ZN(new_n619));
  AOI22_X1  g433(.A1(KEYINPUT31), .A2(new_n619), .B1(new_n602), .B2(new_n582), .ZN(new_n620));
  AOI211_X1 g434(.A(G472), .B(G902), .C1(new_n618), .C2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n604), .B1(new_n621), .B2(KEYINPUT32), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n618), .A2(new_n620), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n561), .A3(new_n320), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT75), .B(KEYINPUT32), .Z(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n560), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n533), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT101), .B(G101), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G3));
  AND3_X1   g445(.A1(new_n575), .A2(KEYINPUT70), .A3(new_n581), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT70), .B1(new_n575), .B2(new_n581), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT31), .B1(new_n634), .B2(new_n595), .ZN(new_n635));
  INV_X1    g449(.A(new_n598), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n574), .B2(new_n575), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n582), .B1(new_n571), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n616), .B2(new_n617), .ZN(new_n640));
  OAI21_X1  g454(.A(G472), .B1(new_n640), .B2(G902), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n624), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n560), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n516), .A2(new_n517), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT84), .B1(new_n644), .B2(new_n502), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n525), .A2(new_n524), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n528), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n471), .A3(new_n320), .ZN(new_n648));
  INV_X1    g462(.A(new_n520), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n532), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n324), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n323), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n327), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n467), .ZN(new_n655));
  INV_X1    g469(.A(new_n382), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n360), .A2(KEYINPUT94), .B1(new_n370), .B2(new_n369), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(new_n367), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n386), .B1(new_n658), .B2(new_n374), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT20), .B1(new_n659), .B2(new_n391), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n388), .A2(new_n329), .A3(new_n389), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n383), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n374), .B1(new_n372), .B2(new_n382), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n320), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G475), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT102), .B(KEYINPUT33), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n449), .A2(new_n450), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n443), .A2(new_n447), .A3(KEYINPUT33), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n670), .A2(G478), .A3(new_n320), .A4(new_n671), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n662), .A2(new_n666), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n655), .A2(new_n465), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n651), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  AOI22_X1  g492(.A1(new_n660), .A2(new_n661), .B1(new_n665), .B2(G475), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n459), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n655), .A2(new_n465), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n651), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT35), .B(G107), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  INV_X1    g498(.A(KEYINPUT36), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n548), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n545), .B(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n556), .B1(new_n557), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n642), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n533), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  INV_X1    g507(.A(G900), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n463), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n462), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n679), .A2(new_n459), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT103), .B1(new_n655), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n698), .ZN(new_n700));
  INV_X1    g514(.A(new_n467), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n653), .B2(new_n327), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n689), .B1(new_n622), .B2(new_n627), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n650), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  XNOR2_X1  g522(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n697), .B(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n530), .A2(new_n532), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n328), .B(new_n715), .Z(new_n716));
  NAND4_X1  g530(.A1(new_n623), .A2(KEYINPUT32), .A3(new_n561), .A4(new_n320), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n609), .A2(new_n613), .B1(new_n582), .B2(new_n576), .ZN(new_n718));
  OAI21_X1  g532(.A(G472), .B1(new_n718), .B2(G902), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n627), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n398), .A2(new_n459), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n688), .A2(new_n701), .A3(new_n721), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n716), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n713), .A2(new_n714), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  NAND2_X1  g539(.A1(new_n667), .A2(new_n672), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n398), .A2(new_n726), .A3(new_n697), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n655), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n706), .A2(new_n650), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  INV_X1    g544(.A(new_n604), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n717), .B(new_n731), .C1(new_n621), .C2(new_n625), .ZN(new_n732));
  INV_X1    g546(.A(new_n560), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(KEYINPUT106), .A2(G469), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n502), .B1(new_n644), .B2(new_n498), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n501), .B1(new_n516), .B2(new_n517), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n512), .B1(new_n738), .B2(KEYINPUT84), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n737), .B1(new_n739), .B2(new_n523), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n736), .B1(new_n740), .B2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n647), .A2(new_n320), .A3(new_n735), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n531), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n734), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n675), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT107), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT41), .B(G113), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n681), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  NAND3_X1  g564(.A1(new_n679), .A2(new_n458), .A3(new_n457), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n465), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n717), .A2(new_n731), .ZN(new_n753));
  AOI21_X1  g567(.A(G902), .B1(new_n618), .B2(new_n620), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n625), .B1(new_n754), .B2(new_n561), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n752), .B(new_n688), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n741), .A2(new_n531), .A3(new_n702), .A4(new_n742), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n221), .ZN(G21));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n754), .B2(new_n561), .ZN(new_n761));
  OAI211_X1 g575(.A(KEYINPUT108), .B(G472), .C1(new_n640), .C2(G902), .ZN(new_n762));
  INV_X1    g576(.A(new_n618), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n635), .B1(new_n577), .B2(new_n581), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n561), .B(new_n320), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n733), .A2(new_n761), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n741), .A2(new_n531), .A3(new_n742), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n398), .A2(new_n459), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n702), .A2(new_n466), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT109), .B(G122), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G24));
  NAND4_X1  g587(.A1(new_n761), .A2(new_n762), .A3(new_n688), .A4(new_n765), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n727), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n673), .A2(KEYINPUT110), .A3(new_n697), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n757), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G125), .ZN(G27));
  NOR2_X1   g596(.A1(new_n778), .A2(KEYINPUT42), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n648), .A2(new_n649), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n328), .A2(new_n701), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n784), .A2(new_n785), .A3(new_n531), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n784), .B1(new_n650), .B2(new_n786), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n628), .B(new_n783), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT32), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n624), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n717), .A3(new_n731), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT110), .B1(new_n673), .B2(new_n697), .ZN(new_n793));
  AND4_X1   g607(.A1(KEYINPUT110), .A2(new_n398), .A3(new_n726), .A4(new_n697), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n795), .A3(new_n733), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n785), .A2(new_n531), .A3(new_n786), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n650), .A2(new_n784), .A3(new_n786), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT42), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n789), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n357), .ZN(G33));
  XNOR2_X1  g617(.A(new_n698), .B(KEYINPUT112), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n628), .B(new_n804), .C1(new_n787), .C2(new_n788), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT113), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n798), .A2(new_n799), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n628), .A4(new_n804), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G134), .ZN(G36));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n519), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT45), .B(new_n508), .C1(new_n518), .C2(new_n502), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(G469), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n471), .A2(new_n320), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(KEYINPUT46), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n648), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT46), .ZN(new_n820));
  INV_X1    g634(.A(new_n815), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n821), .B2(new_n816), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT114), .B1(new_n818), .B2(new_n648), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n531), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(new_n710), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n679), .A2(new_n726), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT43), .Z(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n642), .A3(new_n688), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT44), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n827), .A2(new_n786), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G137), .ZN(G39));
  INV_X1    g649(.A(KEYINPUT47), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT47), .B(new_n531), .C1(new_n823), .C2(new_n824), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n786), .A2(new_n560), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n840), .A2(new_n732), .A3(new_n727), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G140), .ZN(G42));
  NAND3_X1  g657(.A1(new_n733), .A2(new_n531), .A3(new_n469), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n716), .A2(new_n828), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n741), .A2(new_n742), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n720), .B(new_n845), .C1(KEYINPUT49), .C2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(KEYINPUT49), .B2(new_n846), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n829), .A2(new_n462), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n761), .A2(new_n733), .A3(new_n762), .A4(new_n765), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(new_n786), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n837), .A2(KEYINPUT117), .A3(new_n838), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n846), .A2(new_n531), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT117), .B1(new_n837), .B2(new_n838), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n852), .C1(new_n856), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n767), .A2(new_n786), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n849), .ZN(new_n863));
  INV_X1    g677(.A(new_n774), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n862), .ZN(new_n866));
  INV_X1    g680(.A(new_n720), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n733), .A3(new_n462), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n679), .A2(new_n667), .A3(new_n672), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n767), .A2(new_n701), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT119), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n849), .A2(new_n716), .A3(new_n850), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT50), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n872), .A2(KEYINPUT50), .A3(new_n873), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n859), .A2(new_n861), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n560), .B1(new_n622), .B2(new_n791), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n795), .B(new_n885), .C1(new_n787), .C2(new_n788), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n734), .B1(new_n798), .B2(new_n799), .ZN(new_n887));
  AOI22_X1  g701(.A1(KEYINPUT42), .A2(new_n886), .B1(new_n887), .B2(new_n783), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n533), .B1(new_n690), .B2(new_n628), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n628), .B(new_n767), .C1(new_n675), .C2(new_n681), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n780), .A2(new_n706), .A3(new_n752), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n674), .A2(new_n680), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n465), .B(new_n468), .C1(new_n326), .C2(new_n327), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n643), .A2(new_n650), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n771), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n650), .A2(new_n732), .A3(new_n688), .ZN(new_n899));
  INV_X1    g713(.A(new_n697), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT115), .B1(new_n751), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT115), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n460), .A2(new_n902), .A3(new_n697), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n786), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT116), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n901), .A2(new_n786), .A3(new_n903), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n899), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n810), .A2(new_n888), .A3(new_n897), .A4(new_n910), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n655), .A2(new_n688), .A3(new_n900), .A4(new_n721), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n650), .A3(new_n720), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n707), .A2(new_n781), .A3(new_n729), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT52), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n899), .A2(new_n705), .B1(new_n779), .B2(new_n780), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(KEYINPUT52), .A3(new_n729), .A4(new_n913), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n884), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n850), .A2(new_n743), .A3(new_n769), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n758), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n895), .A3(new_n889), .A4(new_n890), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n923), .A2(new_n802), .A3(new_n909), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n916), .A2(new_n918), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n884), .B1(new_n917), .B2(new_n915), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n924), .A2(new_n810), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT54), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n917), .A2(new_n915), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n884), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n924), .A2(new_n810), .A3(new_n925), .A4(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT54), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n920), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n863), .A2(new_n885), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT48), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n461), .B(G953), .C1(new_n851), .C2(new_n780), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n936), .B(new_n937), .C1(new_n674), .C2(new_n868), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n881), .B(new_n870), .C1(new_n876), .C2(new_n877), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n852), .B1(new_n839), .B2(new_n854), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n929), .A2(new_n934), .A3(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n882), .A2(new_n883), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(G952), .A2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n848), .B1(new_n943), .B2(new_n944), .ZN(G75));
  NOR2_X1   g759(.A1(new_n350), .A2(G952), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n320), .B1(new_n920), .B2(new_n932), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(new_n325), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n259), .A2(new_n294), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n292), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT56), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n947), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n948), .A2(G210), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n956), .B2(new_n953), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(G51));
  XNOR2_X1  g772(.A(new_n740), .B(KEYINPUT121), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n920), .A2(new_n932), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n933), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n816), .B(KEYINPUT57), .Z(new_n962));
  OAI21_X1  g776(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n948), .A2(new_n821), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n946), .B1(new_n963), .B2(new_n964), .ZN(G54));
  AND2_X1   g779(.A1(KEYINPUT58), .A2(G475), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n948), .A2(new_n388), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n388), .B1(new_n948), .B2(new_n966), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n967), .A2(new_n968), .A3(new_n946), .ZN(G60));
  XNOR2_X1  g783(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n453), .A2(new_n320), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n929), .B2(new_n934), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n670), .B2(new_n671), .ZN(new_n974));
  INV_X1    g788(.A(new_n972), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n670), .A2(new_n671), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n947), .B1(new_n961), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n974), .A2(new_n977), .ZN(G63));
  NAND2_X1  g792(.A1(G217), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT60), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n920), .B2(new_n932), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n947), .B1(new_n981), .B2(new_n549), .ZN(new_n982));
  AOI211_X1 g796(.A(new_n687), .B(new_n980), .C1(new_n920), .C2(new_n932), .ZN(new_n983));
  OAI211_X1 g797(.A(KEYINPUT123), .B(KEYINPUT61), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n687), .ZN(new_n986));
  INV_X1    g800(.A(new_n980), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n960), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n988), .B(new_n947), .C1(new_n549), .C2(new_n981), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT61), .B1(new_n989), .B2(KEYINPUT123), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n985), .A2(new_n990), .ZN(G66));
  OAI21_X1  g805(.A(G953), .B1(new_n464), .B2(new_n290), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT124), .Z(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n897), .B2(G953), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n950), .B1(G898), .B2(new_n350), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(G69));
  AOI21_X1  g810(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n885), .A2(new_n702), .A3(new_n768), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n826), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT126), .Z(new_n1000));
  AND2_X1   g814(.A1(new_n834), .A2(new_n842), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n917), .A2(new_n729), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n810), .A2(new_n888), .A3(new_n1003), .ZN(new_n1004));
  AND4_X1   g818(.A1(new_n350), .A2(new_n1000), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n593), .A2(new_n594), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT125), .Z(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(new_n384), .Z(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n694), .B2(new_n350), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n711), .A2(new_n628), .A3(new_n786), .A4(new_n893), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g827(.A(new_n724), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1013), .B1(new_n1014), .B2(new_n1002), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1003), .A2(KEYINPUT62), .A3(new_n724), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(G953), .B1(new_n1001), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1018), .A2(new_n1008), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n997), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n997), .ZN(new_n1021));
  OAI221_X1 g835(.A(new_n1021), .B1(new_n1018), .B2(new_n1008), .C1(new_n1005), .C2(new_n1009), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1020), .A2(new_n1022), .ZN(G72));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n619), .A2(new_n597), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n928), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1001), .A2(new_n1017), .A3(new_n897), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1028), .A2(new_n1025), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n581), .B1(new_n595), .B2(new_n596), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n947), .B(new_n1027), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1000), .A2(new_n897), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1032));
  AOI21_X1  g846(.A(KEYINPUT127), .B1(new_n1032), .B2(new_n1025), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n613), .A2(new_n575), .A3(new_n582), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1032), .A2(KEYINPUT127), .A3(new_n1025), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(G57));
endmodule


