//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND2_X1  g0042(.A1(KEYINPUT66), .A2(G1), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g0044(.A1(KEYINPUT66), .A2(G1), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g0046(.A1(new_n246), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT66), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .A4(new_n243), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n213), .A2(G33), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT68), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n212), .B1(new_n206), .B2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n255), .A2(new_n202), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n263), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n254), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n250), .A2(new_n243), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n213), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n264), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT9), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G41), .A2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(new_n249), .A4(G274), .ZN(new_n277));
  INV_X1    g0077(.A(new_n274), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(G77), .ZN(new_n280));
  MUX2_X1   g0080(.A(G222), .B(G223), .S(G1698), .Z(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n277), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n278), .B1(new_n246), .B2(new_n276), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT67), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n290), .B2(G226), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G190), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n272), .B(new_n292), .C1(new_n293), .C2(new_n291), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n291), .A2(G169), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(new_n271), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n260), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n269), .A2(KEYINPUT74), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT74), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n268), .B2(new_n260), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n305), .A2(new_n266), .B1(new_n254), .B2(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT16), .ZN(new_n307));
  INV_X1    g0107(.A(G58), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n217), .ZN(new_n309));
  OAI21_X1  g0109(.A(G20), .B1(new_n309), .B2(new_n201), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n256), .A2(G159), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n285), .A2(new_n213), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n213), .A2(KEYINPUT7), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT72), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT72), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n217), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT73), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n313), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n314), .A2(new_n315), .B1(new_n320), .B2(new_n321), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n326), .A2(KEYINPUT73), .A3(new_n217), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n307), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n217), .B1(new_n314), .B2(KEYINPUT7), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n315), .A2(new_n213), .A3(new_n285), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n312), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n265), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n306), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(G232), .B(new_n274), .C1(new_n267), .C2(new_n275), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n277), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n283), .A2(new_n284), .A3(G226), .A4(G1698), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT75), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n279), .A2(KEYINPUT75), .A3(G226), .A4(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G87), .ZN(new_n340));
  INV_X1    g0140(.A(G1698), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n279), .A2(G223), .A3(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n338), .A2(new_n339), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n335), .B1(new_n343), .B2(new_n278), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(G179), .B2(new_n344), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n333), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT18), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT76), .ZN(new_n350));
  AOI211_X1 g0150(.A(G190), .B(new_n335), .C1(new_n278), .C2(new_n343), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n343), .A2(new_n278), .ZN(new_n352));
  INV_X1    g0152(.A(new_n335), .ZN(new_n353));
  AOI21_X1  g0153(.A(G200), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(KEYINPUT76), .C1(G200), .C2(new_n344), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n333), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT77), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n362), .A3(new_n333), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n361), .A2(KEYINPUT78), .A3(KEYINPUT17), .A4(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n359), .A2(new_n362), .A3(new_n333), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n359), .B2(new_n333), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT17), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n360), .B2(KEYINPUT17), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n349), .B(new_n364), .C1(new_n368), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n255), .A2(new_n217), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT12), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n374));
  INV_X1    g0174(.A(G77), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n259), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n263), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT11), .ZN(new_n378));
  INV_X1    g0178(.A(new_n266), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(G68), .A3(new_n269), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n373), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n277), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n228), .A2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G226), .B2(G1698), .ZN(new_n384));
  INV_X1    g0184(.A(G97), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n384), .A2(new_n285), .B1(new_n262), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n386), .B2(new_n278), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n288), .B(KEYINPUT67), .ZN(new_n388));
  INV_X1    g0188(.A(G238), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  INV_X1    g0191(.A(new_n387), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n290), .B2(G238), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT14), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(G169), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n391), .A2(new_n395), .A3(G179), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n396), .B2(G169), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n381), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n396), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n381), .B1(new_n403), .B2(G190), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n396), .A2(G200), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT70), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n391), .A2(new_n395), .A3(G190), .ZN(new_n407));
  INV_X1    g0207(.A(new_n381), .ZN(new_n408));
  AND4_X1   g0208(.A1(KEYINPUT70), .A2(new_n405), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n402), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n379), .A2(G77), .A3(new_n269), .ZN(new_n411));
  XOR2_X1   g0211(.A(KEYINPUT15), .B(G87), .Z(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n258), .ZN(new_n414));
  INV_X1    g0214(.A(new_n256), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n260), .A2(new_n415), .B1(new_n213), .B2(new_n375), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n263), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n411), .B(new_n417), .C1(G77), .C2(new_n254), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n285), .A2(G1698), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(G232), .B1(G107), .B2(new_n285), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n279), .A2(G1698), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n216), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n382), .B1(new_n422), .B2(new_n278), .ZN(new_n423));
  INV_X1    g0223(.A(G244), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(new_n388), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n418), .B1(G200), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n356), .B2(new_n425), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n425), .A2(G179), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n345), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n418), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NOR4_X1   g0231(.A1(new_n300), .A2(new_n371), .A3(new_n410), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT81), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n274), .A2(G274), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT5), .B(G41), .Z(new_n435));
  NAND3_X1  g0235(.A1(new_n250), .A2(G45), .A3(new_n243), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n436), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT5), .B(G41), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n278), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(G270), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n279), .A2(G264), .A3(G1698), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n285), .A2(G303), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n279), .A2(G257), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(G1698), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n278), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n293), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT20), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n213), .ZN(new_n452));
  AND2_X1   g0252(.A1(KEYINPUT79), .A2(G97), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT79), .A2(G97), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n455), .B2(new_n262), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n263), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n450), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n459), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n453), .A2(new_n454), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G33), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n461), .B(KEYINPUT20), .C1(new_n463), .C2(new_n452), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n255), .A2(new_n457), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n246), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n254), .A2(G116), .A3(new_n265), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n433), .B1(new_n449), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n469), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(KEYINPUT81), .C1(new_n293), .C2(new_n448), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n470), .B(new_n472), .C1(new_n356), .C2(new_n447), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n345), .B1(new_n441), .B2(new_n446), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n448), .A2(new_n469), .A3(G179), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n469), .A2(new_n474), .A3(KEYINPUT21), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n419), .A2(KEYINPUT83), .A3(G250), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n279), .A2(G250), .A3(new_n341), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G294), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n444), .A2(new_n341), .B1(new_n262), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n278), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n437), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n440), .A2(G264), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n491), .A2(G190), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n487), .B2(new_n484), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n492), .B(new_n493), .C1(new_n495), .C2(new_n274), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n279), .A2(new_n213), .A3(G87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT22), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT22), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n279), .A2(new_n500), .A3(new_n213), .A4(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT24), .ZN(new_n503));
  INV_X1    g0303(.A(G107), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G20), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT23), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G116), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n505), .A2(KEYINPUT23), .B1(G20), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n505), .B2(KEYINPUT23), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n502), .A2(new_n503), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n503), .B1(new_n502), .B2(new_n512), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n263), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n254), .A2(new_n265), .A3(new_n467), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT25), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n254), .B2(G107), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n247), .A2(new_n253), .A3(KEYINPUT25), .A4(new_n504), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n517), .A2(G107), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n494), .A2(new_n497), .A3(new_n516), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n256), .A2(G77), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT6), .ZN(new_n524));
  AND2_X1   g0324(.A1(G97), .A2(G107), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G97), .A2(G107), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n462), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G20), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n523), .B(new_n530), .C1(new_n326), .C2(new_n504), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n263), .B1(new_n385), .B2(new_n255), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n517), .A2(G97), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n283), .A2(new_n284), .A3(G250), .A4(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n283), .A2(new_n284), .A3(G244), .A4(new_n341), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT4), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n451), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n278), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n440), .A2(G257), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n492), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n532), .A2(new_n533), .B1(new_n345), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n539), .A2(new_n540), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n297), .A3(new_n492), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(G190), .A3(new_n492), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(G200), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n546), .A2(new_n533), .A3(new_n532), .A4(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n522), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n491), .A2(new_n297), .A3(new_n492), .A4(new_n493), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n496), .A2(new_n345), .ZN(new_n551));
  INV_X1    g0351(.A(new_n515), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n265), .B1(new_n552), .B2(new_n513), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n517), .A2(G107), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n519), .A2(new_n520), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n550), .B(new_n551), .C1(new_n553), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G87), .A2(G107), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n462), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n213), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n279), .A2(new_n213), .A3(G68), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n462), .B2(new_n258), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n263), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n254), .A2(new_n265), .A3(new_n412), .A4(new_n467), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(new_n568), .C1(new_n254), .C2(new_n412), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n389), .A2(new_n341), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n424), .A2(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n279), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n274), .B1(new_n572), .B2(new_n509), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(G274), .ZN(new_n575));
  INV_X1    g0375(.A(new_n212), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(new_n273), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT80), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n438), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT80), .B1(new_n434), .B2(new_n436), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n436), .A2(G250), .A3(new_n274), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n574), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n345), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n574), .A2(new_n581), .A3(new_n297), .A4(new_n582), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n569), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(G200), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n255), .A2(new_n413), .B1(new_n566), .B2(new_n263), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n574), .A2(new_n581), .A3(G190), .A4(new_n582), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n254), .A2(G87), .A3(new_n265), .A4(new_n467), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n557), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n432), .A2(new_n483), .A3(new_n549), .A4(new_n592), .ZN(G372));
  INV_X1    g0393(.A(new_n299), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n430), .A2(KEYINPUT87), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT87), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n428), .A2(new_n596), .A3(new_n418), .A4(new_n429), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n595), .B(new_n597), .C1(new_n406), .C2(new_n409), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n402), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n599), .B(new_n364), .C1(new_n368), .C2(new_n370), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n349), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n594), .B1(new_n601), .B2(new_n295), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n569), .A2(new_n585), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n581), .A2(KEYINPUT84), .A3(new_n582), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT84), .B1(new_n581), .B2(new_n582), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n574), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n345), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(G200), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(KEYINPUT85), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT85), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n611), .A3(G200), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n607), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n542), .A2(new_n544), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n542), .A2(new_n544), .A3(new_n586), .A4(new_n591), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n607), .B1(new_n617), .B2(KEYINPUT26), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(KEYINPUT86), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n557), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(new_n480), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n549), .A2(new_n613), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT86), .B1(new_n616), .B2(new_n618), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n432), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n602), .A2(new_n626), .ZN(G369));
  INV_X1    g0427(.A(G13), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n628), .A2(G20), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n246), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n631), .A2(KEYINPUT88), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(KEYINPUT88), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(G213), .B1(new_n630), .B2(KEYINPUT27), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n471), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n480), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n482), .B2(new_n640), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G330), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n557), .A2(new_n638), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n638), .B1(new_n553), .B2(new_n556), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n522), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n647), .B2(new_n557), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n481), .A2(new_n638), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(G399));
  NOR2_X1   g0452(.A1(new_n559), .A2(G116), .ZN(new_n653));
  INV_X1    g0453(.A(new_n207), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n656), .A3(G1), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n210), .B2(new_n656), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT28), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT29), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n625), .A2(new_n660), .A3(new_n639), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n620), .B2(new_n480), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n478), .A2(new_n479), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(new_n557), .A3(KEYINPUT90), .A4(new_n477), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n664), .A2(new_n613), .A3(new_n549), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n581), .A2(new_n582), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT84), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n581), .A2(KEYINPUT84), .A3(new_n582), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n573), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n585), .B(new_n569), .C1(new_n672), .C2(G169), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n617), .B2(KEYINPUT26), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT85), .B1(new_n672), .B2(new_n293), .ZN(new_n675));
  INV_X1    g0475(.A(new_n608), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n612), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n615), .A3(new_n673), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n674), .B1(new_n678), .B2(KEYINPUT26), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n667), .B1(new_n679), .B2(KEYINPUT89), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT89), .ZN(new_n681));
  AOI211_X1 g0481(.A(new_n681), .B(new_n674), .C1(KEYINPUT26), .C2(new_n678), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n639), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n683), .A2(KEYINPUT29), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n662), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n483), .A2(new_n549), .A3(new_n592), .A4(new_n639), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n448), .A2(G179), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n491), .A2(new_n493), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n583), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n543), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n687), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(KEYINPUT30), .A3(new_n543), .A4(new_n691), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n448), .A2(G179), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n606), .A3(new_n541), .A4(new_n496), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n638), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n638), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n686), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n685), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n659), .B1(new_n706), .B2(G1), .ZN(G364));
  AOI21_X1  g0507(.A(new_n249), .B1(new_n629), .B2(G45), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n656), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n279), .A2(new_n207), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(KEYINPUT91), .B2(G355), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(KEYINPUT91), .B2(G355), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(G116), .B2(new_n207), .ZN(new_n714));
  INV_X1    g0514(.A(G45), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n238), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n654), .A2(new_n279), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n211), .B2(new_n715), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n714), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n212), .B1(G20), .B2(new_n345), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n710), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n213), .A2(new_n356), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n293), .A2(G179), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT94), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT94), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n297), .A2(G200), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n213), .A2(G190), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT93), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n737), .B1(new_n735), .B2(new_n736), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n734), .A2(G303), .B1(G311), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n736), .A2(new_n729), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n285), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n736), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(G329), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n213), .B1(new_n746), .B2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n356), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n751), .A2(G294), .B1(G326), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n742), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n728), .A2(new_n735), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n752), .A2(G190), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT33), .B(G317), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n757), .A2(G322), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT95), .Z(new_n761));
  NAND2_X1  g0561(.A1(new_n734), .A2(G87), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n756), .B(KEYINPUT92), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G58), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n741), .A2(G77), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n279), .B1(new_n743), .B2(new_n504), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G50), .B2(new_n753), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n762), .A2(new_n765), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n750), .A2(new_n385), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n748), .A2(G159), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(KEYINPUT32), .ZN(new_n772));
  INV_X1    g0572(.A(new_n758), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n772), .B1(KEYINPUT32), .B2(new_n771), .C1(new_n217), .C2(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n755), .A2(new_n761), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n727), .B1(new_n775), .B2(new_n724), .ZN(new_n776));
  INV_X1    g0576(.A(new_n723), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n642), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n643), .A2(new_n709), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n642), .A2(G330), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(G396));
  NAND2_X1  g0581(.A1(new_n625), .A2(new_n639), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n595), .A2(new_n418), .A3(new_n597), .A4(new_n638), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n638), .A2(new_n418), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n427), .A2(new_n430), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n785), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n639), .B(new_n788), .C1(new_n623), .C2(new_n624), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n710), .B1(new_n790), .B2(new_n704), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n704), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n724), .A2(new_n721), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n710), .B1(G77), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G150), .ZN(new_n796));
  INV_X1    g0596(.A(new_n753), .ZN(new_n797));
  INV_X1    g0597(.A(G137), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n773), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n740), .A2(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n799), .B(new_n801), .C1(G143), .C2(new_n764), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT34), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n279), .B1(new_n747), .B2(new_n804), .C1(new_n217), .C2(new_n743), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G58), .B2(new_n751), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n202), .B2(new_n733), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n770), .B1(new_n758), .B2(G283), .ZN(new_n808));
  INV_X1    g0608(.A(G303), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n797), .ZN(new_n810));
  INV_X1    g0610(.A(G87), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n743), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n285), .B1(new_n756), .B2(new_n489), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G311), .C2(new_n748), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n814), .B1(new_n504), .B2(new_n733), .C1(new_n457), .C2(new_n740), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n803), .A2(new_n807), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n795), .B1(new_n816), .B2(new_n724), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n788), .B2(new_n722), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n792), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G384));
  OAI21_X1  g0620(.A(G77), .B1(new_n308), .B2(new_n217), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n821), .A2(new_n210), .B1(G50), .B2(new_n217), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n822), .A2(new_n628), .A3(new_n267), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT96), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n825), .A2(G116), .A3(new_n214), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT36), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n381), .A2(new_n638), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n410), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n402), .B(new_n831), .C1(new_n406), .C2(new_n409), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n786), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT101), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n703), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n686), .A2(new_n701), .A3(KEYINPUT101), .A4(new_n702), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n361), .A2(new_n363), .ZN(new_n841));
  INV_X1    g0641(.A(new_n306), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n332), .B1(KEYINPUT16), .B2(new_n331), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n347), .A2(new_n636), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n365), .A2(new_n366), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n333), .A2(new_n636), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n348), .A2(new_n847), .A3(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n636), .B1(new_n842), .B2(new_n843), .ZN(new_n850));
  AOI221_X4 g0650(.A(new_n840), .B1(new_n845), .B2(new_n849), .C1(new_n371), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n371), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n845), .A2(new_n849), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT38), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT97), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n851), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n852), .A2(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n840), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT97), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n839), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT40), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n371), .A2(new_n847), .ZN(new_n865));
  INV_X1    g0665(.A(new_n360), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n333), .B1(new_n347), .B2(new_n636), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(KEYINPUT98), .A2(new_n868), .B1(new_n846), .B2(new_n848), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(KEYINPUT98), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n864), .B1(new_n851), .B2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n371), .A2(new_n847), .B1(new_n869), .B2(new_n870), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n859), .B(KEYINPUT102), .C1(new_n874), .C2(KEYINPUT38), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n873), .A2(new_n839), .A3(KEYINPUT40), .A4(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n863), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n837), .A2(new_n838), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(new_n432), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n879), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n880), .A2(G330), .A3(new_n881), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n402), .A2(new_n638), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT39), .B1(new_n851), .B2(new_n854), .ZN(new_n884));
  XNOR2_X1  g0684(.A(KEYINPUT99), .B(KEYINPUT39), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n859), .B(new_n885), .C1(new_n874), .C2(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT100), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n884), .A2(KEYINPUT100), .A3(new_n886), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n636), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n349), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n856), .A2(new_n860), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n833), .A2(new_n834), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n430), .A2(new_n638), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n789), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n894), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n891), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n432), .B1(new_n662), .B2(new_n684), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n903), .A2(new_n602), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n902), .B(new_n904), .Z(new_n905));
  OAI22_X1  g0705(.A1(new_n882), .A2(new_n905), .B1(new_n246), .B2(new_n629), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n882), .A2(new_n905), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n830), .B1(new_n906), .B2(new_n907), .ZN(G367));
  NAND2_X1  g0708(.A1(new_n588), .A2(new_n590), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n638), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n673), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT103), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n613), .A2(new_n910), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT104), .Z(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n723), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n740), .A2(new_n744), .B1(new_n504), .B2(new_n750), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT108), .Z(new_n918));
  NOR2_X1   g0718(.A1(new_n733), .A2(new_n457), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT46), .ZN(new_n920));
  INV_X1    g0720(.A(G317), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n285), .B1(new_n747), .B2(new_n921), .C1(new_n462), .C2(new_n743), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(KEYINPUT109), .B(G311), .Z(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(new_n753), .B1(G294), .B2(new_n758), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n925), .C1(new_n809), .C2(new_n763), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n918), .A2(new_n920), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT110), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n279), .B1(new_n747), .B2(new_n798), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n756), .A2(new_n796), .B1(new_n743), .B2(new_n375), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n930), .B(new_n931), .C1(new_n741), .C2(G50), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n750), .A2(new_n217), .ZN(new_n933));
  INV_X1    g0733(.A(G143), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n797), .A2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(G159), .C2(new_n758), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n932), .B(new_n936), .C1(new_n308), .C2(new_n733), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT111), .Z(new_n938));
  NAND2_X1  g0738(.A1(new_n928), .A2(KEYINPUT110), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n929), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT47), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n724), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n725), .B1(new_n207), .B2(new_n413), .C1(new_n234), .C2(new_n718), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n916), .A2(new_n710), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n915), .B(KEYINPUT43), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n532), .A2(new_n533), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n545), .B(new_n548), .C1(new_n946), .C2(new_n639), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n615), .A2(new_n638), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(new_n648), .A3(new_n650), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n545), .B1(new_n947), .B2(new_n557), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(new_n639), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n945), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT105), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n955), .A2(new_n960), .A3(new_n915), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n945), .A2(KEYINPUT105), .A3(new_n956), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n649), .A2(new_n949), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n959), .A2(new_n964), .A3(new_n961), .A4(new_n962), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n708), .B(KEYINPUT107), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n651), .A2(new_n950), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n651), .A2(new_n950), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n649), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n648), .B(new_n650), .Z(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n644), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n706), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n985));
  XNOR2_X1  g0785(.A(new_n655), .B(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n970), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n944), .B1(new_n968), .B2(new_n988), .ZN(G387));
  AOI22_X1  g0789(.A1(new_n924), .A2(new_n758), .B1(G322), .B2(new_n753), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n740), .B2(new_n809), .C1(new_n763), .C2(new_n921), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT48), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n734), .A2(G294), .B1(G283), .B2(new_n751), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT49), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n743), .A2(new_n457), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n279), .B(new_n999), .C1(G326), .C2(new_n748), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n997), .A2(KEYINPUT49), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n751), .A2(new_n412), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n773), .B2(new_n260), .C1(new_n800), .C2(new_n797), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n743), .A2(new_n385), .B1(new_n747), .B2(new_n796), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n285), .B(new_n1005), .C1(G50), .C2(new_n757), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n734), .A2(G77), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n741), .A2(G68), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1001), .A2(new_n1002), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1010), .A2(new_n724), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n653), .B(new_n715), .C1(new_n217), .C2(new_n375), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT113), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT113), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n260), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT50), .B1(new_n260), .B2(G50), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n717), .C1(new_n715), .C2(new_n231), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n653), .A2(new_n711), .B1(G107), .B2(new_n207), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT112), .Z(new_n1020));
  AND2_X1   g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n710), .B1(new_n1021), .B2(new_n726), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1011), .A2(KEYINPUT114), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT114), .B1(new_n1011), .B2(new_n1022), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n648), .C2(new_n777), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n705), .A2(new_n983), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n705), .A2(new_n983), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n655), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1025), .B1(new_n983), .B2(new_n969), .C1(new_n1029), .C2(new_n1030), .ZN(G393));
  INV_X1    g0831(.A(KEYINPUT116), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n980), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(new_n978), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n970), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n725), .B1(new_n207), .B2(new_n462), .C1(new_n241), .C2(new_n718), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n710), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n750), .A2(new_n375), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n279), .B1(new_n747), .B2(new_n934), .C1(new_n811), .C2(new_n743), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G50), .C2(new_n758), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n797), .A2(new_n796), .B1(new_n756), .B2(new_n800), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT51), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n734), .A2(G68), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n741), .A2(new_n301), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n285), .B1(new_n743), .B2(new_n504), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n773), .A2(new_n809), .B1(new_n750), .B2(new_n457), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(G322), .C2(new_n748), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n744), .B2(new_n733), .C1(new_n489), .C2(new_n740), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n757), .A2(G311), .B1(G317), .B2(new_n753), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1045), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1037), .B1(new_n1052), .B2(new_n724), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n950), .B2(new_n777), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1028), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1055), .A2(new_n1034), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n655), .B1(new_n1028), .B2(new_n981), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1035), .B(new_n1054), .C1(new_n1056), .C2(new_n1057), .ZN(G390));
  NAND2_X1  g0858(.A1(new_n900), .A2(new_n883), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n889), .A2(new_n890), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n883), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n639), .B(new_n788), .C1(new_n680), .C2(new_n682), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n898), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n833), .A2(new_n834), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n873), .A3(new_n875), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n835), .A2(new_n837), .A3(G330), .A4(new_n838), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n704), .A2(new_n786), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n1064), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1066), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1060), .A2(new_n1073), .A3(KEYINPUT117), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT117), .B1(new_n1060), .B2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n884), .A2(KEYINPUT100), .A3(new_n886), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT100), .B1(new_n884), .B2(new_n886), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n1078), .A3(new_n722), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n756), .A2(new_n457), .B1(new_n747), .B2(new_n489), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n743), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n279), .B(new_n1080), .C1(G68), .C2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n797), .A2(new_n744), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1038), .B(new_n1083), .C1(G107), .C2(new_n758), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n741), .A2(new_n455), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n762), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n733), .A2(new_n796), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G125), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n756), .A2(new_n804), .B1(new_n747), .B2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n773), .A2(new_n798), .B1(new_n750), .B2(new_n800), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G128), .C2(new_n753), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT54), .B(G143), .Z(new_n1094));
  OAI21_X1  g0894(.A(new_n279), .B1(new_n743), .B2(new_n202), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n741), .A2(new_n1094), .B1(KEYINPUT119), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1093), .B(new_n1096), .C1(KEYINPUT119), .C2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1086), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n724), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n710), .C1(new_n301), .C2(new_n794), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1076), .A2(new_n969), .B1(new_n1079), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1068), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT117), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n899), .A2(new_n1061), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1077), .A2(new_n1078), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1066), .A2(new_n1072), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1060), .A2(new_n1073), .A3(KEYINPUT117), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1103), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n878), .A2(G330), .A3(new_n788), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n896), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1063), .B1(new_n1071), .B2(new_n1064), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n789), .A2(new_n898), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1068), .B1(new_n1071), .B2(new_n1064), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1112), .A2(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n878), .A2(G330), .A3(new_n432), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n903), .A2(new_n602), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n655), .B1(new_n1110), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1070), .B(new_n1119), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1120), .A2(new_n1122), .A3(KEYINPUT118), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT118), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1119), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n656), .B1(new_n1076), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1124), .B1(new_n1126), .B2(new_n1121), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1102), .B1(new_n1123), .B2(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(G41), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n285), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G283), .B2(new_n748), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G107), .A2(new_n757), .B1(new_n1081), .B2(G58), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1007), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n797), .A2(new_n457), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n933), .B(new_n1134), .C1(G97), .C2(new_n758), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(new_n413), .C2(new_n740), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT58), .ZN(new_n1137));
  AOI21_X1  g0937(.A(G50), .B1(new_n262), .B2(new_n1129), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1136), .A2(new_n1137), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n734), .A2(new_n1094), .B1(G137), .B2(new_n741), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n757), .A2(G128), .B1(new_n751), .B2(G150), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n758), .A2(G132), .B1(new_n753), .B2(G125), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT59), .Z(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT121), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n262), .B(new_n1129), .C1(new_n743), .C2(new_n800), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G124), .B2(new_n748), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1144), .A2(KEYINPUT121), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1139), .B1(new_n1137), .B2(new_n1136), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n724), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT122), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n710), .B1(G50), .B2(new_n794), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT123), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n892), .A2(new_n271), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT124), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n300), .B(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1159));
  XNOR2_X1  g0959(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1152), .B(new_n1155), .C1(new_n1160), .C2(new_n721), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n863), .A2(G330), .A3(new_n876), .A4(new_n1160), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n858), .A2(KEYINPUT97), .A3(new_n859), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n855), .B1(new_n851), .B2(new_n854), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(G330), .B(new_n876), .C1(new_n1166), .C2(KEYINPUT40), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1160), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n902), .A2(new_n1162), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1061), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n901), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1162), .A2(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1161), .B1(new_n1174), .B2(new_n970), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1118), .B(KEYINPUT125), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1110), .B2(new_n1119), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n902), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n902), .A2(new_n1162), .A3(new_n1169), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n655), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1176), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1121), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1174), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1175), .B1(new_n1183), .B2(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1125), .A2(new_n987), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(G128), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n279), .B1(new_n747), .B2(new_n1190), .C1(new_n308), .C2(new_n743), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n764), .B2(G137), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n797), .A2(new_n804), .B1(new_n750), .B2(new_n202), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n758), .B2(new_n1094), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n734), .A2(G159), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n741), .A2(G150), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1192), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n756), .A2(new_n744), .B1(new_n747), .B2(new_n809), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n279), .B(new_n1198), .C1(G77), .C2(new_n1081), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n385), .B2(new_n733), .C1(new_n504), .C2(new_n740), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1003), .B1(new_n773), .B2(new_n457), .C1(new_n489), .C2(new_n797), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1197), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n724), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n709), .B1(new_n217), .B2(new_n793), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n1064), .C2(new_n722), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1116), .B2(new_n969), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1189), .A2(new_n1207), .ZN(G381));
  OR2_X1    g1008(.A1(G393), .A2(G396), .ZN(new_n1209));
  INV_X1    g1009(.A(G390), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n819), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1209), .A2(new_n1211), .A3(G387), .A4(G381), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1161), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n969), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT57), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1170), .A2(new_n1173), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n656), .B1(new_n1217), .B2(new_n1185), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1177), .B2(new_n1214), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1215), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1101), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1212), .A2(new_n1220), .A3(new_n1221), .ZN(G407));
  NAND2_X1  g1022(.A1(new_n637), .A2(G213), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(G407), .A2(G213), .A3(new_n1225), .ZN(G409));
  NAND2_X1  g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1209), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G387), .A2(new_n1210), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(G387), .A2(new_n1210), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n968), .A2(new_n988), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n944), .A3(G390), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1234), .A2(new_n1229), .A3(new_n1209), .A4(new_n1227), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(KEYINPUT60), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1237), .A2(new_n1188), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n655), .B1(new_n1237), .B2(new_n1188), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1240), .A2(new_n819), .A3(new_n1206), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n819), .B1(new_n1240), .B2(new_n1206), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1242), .A2(G2897), .A3(new_n1224), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1224), .A2(G2897), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1243), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n1241), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1185), .A2(new_n1174), .A3(new_n987), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1175), .A2(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G378), .A2(new_n1220), .B1(new_n1221), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1248), .B1(new_n1251), .B2(new_n1224), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1221), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT118), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1126), .A2(new_n1124), .A3(new_n1121), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1101), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1254), .B1(G375), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1246), .A2(new_n1241), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1223), .A4(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1252), .A2(new_n1253), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G378), .A2(new_n1220), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1224), .B1(new_n1263), .B2(new_n1254), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1259), .B1(new_n1264), .B2(new_n1260), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1236), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1223), .A4(new_n1260), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1232), .A2(new_n1253), .A3(new_n1235), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT126), .B1(new_n1251), .B2(new_n1224), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1258), .A2(new_n1271), .A3(new_n1223), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1248), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1258), .A2(new_n1223), .A3(new_n1260), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1269), .A2(new_n1273), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1266), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1266), .A2(new_n1277), .A3(KEYINPUT127), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(G405));
  INV_X1    g1082(.A(new_n1221), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1263), .B1(new_n1220), .B2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1260), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1236), .ZN(G402));
endmodule


