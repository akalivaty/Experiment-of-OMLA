

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U558 ( .A(n801), .ZN(n782) );
  AND2_X1 U559 ( .A1(n722), .A2(n956), .ZN(n719) );
  INV_X1 U560 ( .A(n956), .ZN(n724) );
  NAND2_X1 U561 ( .A1(n711), .A2(n710), .ZN(n757) );
  NAND2_X1 U562 ( .A1(G160), .A2(G40), .ZN(n709) );
  XOR2_X1 U563 ( .A(KEYINPUT0), .B(G543), .Z(n621) );
  NOR2_X2 U564 ( .A1(n530), .A2(n529), .ZN(G160) );
  INV_X1 U565 ( .A(G2104), .ZN(n525) );
  NOR2_X4 U566 ( .A1(G2105), .A2(n525), .ZN(n893) );
  NAND2_X1 U567 ( .A1(G101), .A2(n893), .ZN(n521) );
  XNOR2_X1 U568 ( .A(n521), .B(KEYINPUT23), .ZN(n522) );
  XNOR2_X1 U569 ( .A(n522), .B(KEYINPUT65), .ZN(n524) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U571 ( .A1(G113), .A2(n890), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n530) );
  AND2_X1 U573 ( .A1(n525), .A2(G2105), .ZN(n889) );
  NAND2_X1 U574 ( .A1(G125), .A2(n889), .ZN(n528) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n526), .Z(n894) );
  NAND2_X1 U577 ( .A1(G137), .A2(n894), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  INV_X1 U579 ( .A(G651), .ZN(n535) );
  NOR2_X1 U580 ( .A1(G543), .A2(n535), .ZN(n531) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n531), .Z(n649) );
  NAND2_X1 U582 ( .A1(G64), .A2(n649), .ZN(n534) );
  NOR2_X1 U583 ( .A1(G651), .A2(n621), .ZN(n532) );
  XNOR2_X2 U584 ( .A(KEYINPUT64), .B(n532), .ZN(n642) );
  NAND2_X1 U585 ( .A1(G52), .A2(n642), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n541) );
  NOR2_X1 U587 ( .A1(n621), .A2(n535), .ZN(n641) );
  NAND2_X1 U588 ( .A1(n641), .A2(G77), .ZN(n536) );
  XOR2_X1 U589 ( .A(KEYINPUT67), .B(n536), .Z(n538) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U591 ( .A1(n645), .A2(G90), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U594 ( .A1(n541), .A2(n540), .ZN(G171) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U596 ( .A1(G99), .A2(n893), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G111), .A2(n890), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U599 ( .A(n544), .B(KEYINPUT77), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G135), .A2(n894), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n889), .A2(G123), .ZN(n547) );
  XOR2_X1 U603 ( .A(KEYINPUT18), .B(n547), .Z(n548) );
  NOR2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U605 ( .A(KEYINPUT78), .B(n550), .Z(n932) );
  XNOR2_X1 U606 ( .A(n932), .B(G2096), .ZN(n551) );
  OR2_X1 U607 ( .A1(G2100), .A2(n551), .ZN(G156) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(n889), .A2(G126), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT84), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G138), .A2(n894), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G102), .A2(n893), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G114), .A2(n890), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U618 ( .A1(n558), .A2(n557), .ZN(G164) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U620 ( .A(n559), .B(KEYINPUT10), .ZN(n560) );
  XNOR2_X1 U621 ( .A(KEYINPUT68), .B(n560), .ZN(G223) );
  INV_X1 U622 ( .A(G223), .ZN(n838) );
  NAND2_X1 U623 ( .A1(n838), .A2(G567), .ZN(n561) );
  XNOR2_X1 U624 ( .A(n561), .B(KEYINPUT69), .ZN(n562) );
  XNOR2_X1 U625 ( .A(KEYINPUT11), .B(n562), .ZN(G234) );
  XOR2_X1 U626 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n564) );
  NAND2_X1 U627 ( .A1(G56), .A2(n649), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G81), .A2(n645), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT71), .B(n565), .Z(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT12), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G68), .A2(n641), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT13), .B(n569), .Z(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G43), .A2(n642), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n948) );
  INV_X1 U638 ( .A(G860), .ZN(n613) );
  OR2_X1 U639 ( .A1(n948), .A2(n613), .ZN(G153) );
  XOR2_X1 U640 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  INV_X1 U641 ( .A(G868), .ZN(n604) );
  NOR2_X1 U642 ( .A1(G301), .A2(n604), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G79), .A2(n641), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G92), .A2(n645), .ZN(n575) );
  NAND2_X1 U645 ( .A1(G66), .A2(n649), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G54), .A2(n642), .ZN(n576) );
  XNOR2_X1 U648 ( .A(KEYINPUT73), .B(n576), .ZN(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  AND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U651 ( .A(KEYINPUT15), .ZN(n581) );
  XNOR2_X2 U652 ( .A(n582), .B(n581), .ZN(n956) );
  AND2_X1 U653 ( .A1(n604), .A2(n956), .ZN(n583) );
  NOR2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U655 ( .A(KEYINPUT74), .B(n585), .ZN(G284) );
  XNOR2_X1 U656 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n597) );
  NAND2_X1 U657 ( .A1(n645), .A2(G89), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT4), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G76), .A2(n641), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U661 ( .A(KEYINPUT5), .B(n589), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n649), .A2(G63), .ZN(n590) );
  XOR2_X1 U663 ( .A(KEYINPUT75), .B(n590), .Z(n592) );
  NAND2_X1 U664 ( .A1(G51), .A2(n642), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT6), .B(n593), .Z(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n597), .B(n596), .ZN(G168) );
  XOR2_X1 U669 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U670 ( .A1(G65), .A2(n649), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G53), .A2(n642), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G91), .A2(n645), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G78), .A2(n641), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n959) );
  INV_X1 U677 ( .A(n959), .ZN(G299) );
  NAND2_X1 U678 ( .A1(G868), .A2(G286), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G299), .A2(n604), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U681 ( .A1(n613), .A2(G559), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n607), .A2(n956), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n948), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G868), .A2(n956), .ZN(n609) );
  NOR2_X1 U686 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G559), .A2(n956), .ZN(n612) );
  XOR2_X1 U689 ( .A(n948), .B(n612), .Z(n657) );
  NAND2_X1 U690 ( .A1(n613), .A2(n657), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G67), .A2(n649), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G55), .A2(n642), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G93), .A2(n645), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G80), .A2(n641), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n661) );
  XOR2_X1 U698 ( .A(n620), .B(n661), .Z(G145) );
  NAND2_X1 U699 ( .A1(n621), .A2(G87), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G49), .A2(n642), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U702 ( .A1(n649), .A2(n624), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G651), .A2(G74), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U705 ( .A1(G86), .A2(n645), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G61), .A2(n649), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n641), .A2(G73), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G48), .A2(n642), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G88), .A2(n645), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G75), .A2(n641), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n642), .A2(G50), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT79), .B(n636), .Z(n638) );
  NAND2_X1 U718 ( .A1(n649), .A2(G62), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U720 ( .A1(n640), .A2(n639), .ZN(G166) );
  NAND2_X1 U721 ( .A1(G72), .A2(n641), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G47), .A2(n642), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G85), .A2(n645), .ZN(n646) );
  XOR2_X1 U725 ( .A(KEYINPUT66), .B(n646), .Z(n647) );
  NOR2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n649), .A2(G60), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(G290) );
  XNOR2_X1 U729 ( .A(KEYINPUT19), .B(G288), .ZN(n656) );
  XOR2_X1 U730 ( .A(G166), .B(n661), .Z(n652) );
  XNOR2_X1 U731 ( .A(G305), .B(n652), .ZN(n653) );
  XNOR2_X1 U732 ( .A(n959), .B(n653), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n904) );
  XNOR2_X1 U735 ( .A(n904), .B(n657), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n658), .B(KEYINPUT80), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n659), .A2(G868), .ZN(n660) );
  XOR2_X1 U738 ( .A(KEYINPUT81), .B(n660), .Z(n663) );
  OR2_X1 U739 ( .A1(n661), .A2(G868), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n664) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n665), .ZN(n667) );
  XNOR2_X1 U744 ( .A(KEYINPUT82), .B(KEYINPUT21), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U746 ( .A1(G2072), .A2(n668), .ZN(G158) );
  XOR2_X1 U747 ( .A(KEYINPUT83), .B(G44), .Z(n669) );
  XNOR2_X1 U748 ( .A(KEYINPUT3), .B(n669), .ZN(G218) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U751 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U752 ( .A1(G96), .A2(n672), .ZN(n842) );
  NAND2_X1 U753 ( .A1(G2106), .A2(n842), .ZN(n676) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n673) );
  NOR2_X1 U755 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U756 ( .A1(G108), .A2(n674), .ZN(n843) );
  NAND2_X1 U757 ( .A1(G567), .A2(n843), .ZN(n675) );
  NAND2_X1 U758 ( .A1(n676), .A2(n675), .ZN(n844) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U760 ( .A1(n844), .A2(n677), .ZN(n841) );
  NAND2_X1 U761 ( .A1(n841), .A2(G36), .ZN(G176) );
  XNOR2_X1 U762 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n711), .A2(n709), .ZN(n823) );
  XNOR2_X1 U765 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n682) );
  NAND2_X1 U766 ( .A1(G128), .A2(n889), .ZN(n679) );
  NAND2_X1 U767 ( .A1(G116), .A2(n890), .ZN(n678) );
  NAND2_X1 U768 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U769 ( .A(n680), .B(KEYINPUT35), .ZN(n681) );
  XNOR2_X1 U770 ( .A(n682), .B(n681), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G104), .A2(n893), .ZN(n684) );
  NAND2_X1 U772 ( .A1(G140), .A2(n894), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n685), .ZN(n686) );
  NOR2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U776 ( .A(KEYINPUT36), .B(n688), .Z(n689) );
  XNOR2_X1 U777 ( .A(KEYINPUT89), .B(n689), .ZN(n879) );
  XNOR2_X1 U778 ( .A(KEYINPUT37), .B(G2067), .ZN(n821) );
  NOR2_X1 U779 ( .A1(n879), .A2(n821), .ZN(n924) );
  NAND2_X1 U780 ( .A1(n823), .A2(n924), .ZN(n818) );
  NAND2_X1 U781 ( .A1(G107), .A2(n890), .ZN(n690) );
  XNOR2_X1 U782 ( .A(n690), .B(KEYINPUT90), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n893), .A2(G95), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U785 ( .A1(G119), .A2(n889), .ZN(n694) );
  NAND2_X1 U786 ( .A1(G131), .A2(n894), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n882) );
  INV_X1 U789 ( .A(G1991), .ZN(n994) );
  NOR2_X1 U790 ( .A1(n882), .A2(n994), .ZN(n706) );
  NAND2_X1 U791 ( .A1(n889), .A2(G129), .ZN(n703) );
  NAND2_X1 U792 ( .A1(G141), .A2(n894), .ZN(n698) );
  NAND2_X1 U793 ( .A1(G117), .A2(n890), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n893), .A2(G105), .ZN(n699) );
  XOR2_X1 U796 ( .A(KEYINPUT38), .B(n699), .Z(n700) );
  NOR2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U799 ( .A(KEYINPUT91), .B(n704), .ZN(n878) );
  INV_X1 U800 ( .A(G1996), .ZN(n812) );
  NOR2_X1 U801 ( .A1(n878), .A2(n812), .ZN(n705) );
  NOR2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n927) );
  INV_X1 U803 ( .A(n823), .ZN(n707) );
  NOR2_X1 U804 ( .A1(n927), .A2(n707), .ZN(n815) );
  INV_X1 U805 ( .A(n815), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n818), .A2(n708), .ZN(n808) );
  INV_X1 U807 ( .A(n709), .ZN(n710) );
  NAND2_X1 U808 ( .A1(G1348), .A2(n757), .ZN(n712) );
  XOR2_X1 U809 ( .A(KEYINPUT97), .B(n712), .Z(n714) );
  INV_X1 U810 ( .A(n757), .ZN(n740) );
  NAND2_X1 U811 ( .A1(G2067), .A2(n740), .ZN(n713) );
  NAND2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U813 ( .A(n715), .B(KEYINPUT98), .ZN(n721) );
  NOR2_X1 U814 ( .A1(n757), .A2(n812), .ZN(n716) );
  XOR2_X1 U815 ( .A(n716), .B(KEYINPUT26), .Z(n718) );
  NAND2_X1 U816 ( .A1(n757), .A2(G1341), .ZN(n717) );
  AND2_X1 U817 ( .A1(n718), .A2(n717), .ZN(n723) );
  INV_X1 U818 ( .A(n948), .ZN(n722) );
  NAND2_X1 U819 ( .A1(n723), .A2(n719), .ZN(n720) );
  NAND2_X1 U820 ( .A1(n721), .A2(n720), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U822 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U823 ( .A1(n727), .A2(n726), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n740), .A2(G2072), .ZN(n728) );
  XNOR2_X1 U825 ( .A(n728), .B(KEYINPUT27), .ZN(n730) );
  AND2_X1 U826 ( .A1(G1956), .A2(n757), .ZN(n729) );
  NOR2_X1 U827 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U828 ( .A1(n733), .A2(n959), .ZN(n731) );
  NAND2_X1 U829 ( .A1(n732), .A2(n731), .ZN(n737) );
  NOR2_X1 U830 ( .A1(n733), .A2(n959), .ZN(n735) );
  XOR2_X1 U831 ( .A(KEYINPUT28), .B(KEYINPUT96), .Z(n734) );
  XNOR2_X1 U832 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U833 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U834 ( .A(KEYINPUT29), .B(n738), .ZN(n745) );
  XNOR2_X1 U835 ( .A(G2078), .B(KEYINPUT25), .ZN(n739) );
  XNOR2_X1 U836 ( .A(n739), .B(KEYINPUT94), .ZN(n997) );
  NOR2_X1 U837 ( .A1(n997), .A2(n757), .ZN(n742) );
  INV_X1 U838 ( .A(G1961), .ZN(n983) );
  NOR2_X1 U839 ( .A1(n740), .A2(n983), .ZN(n741) );
  NOR2_X1 U840 ( .A1(n742), .A2(n741), .ZN(n750) );
  NAND2_X1 U841 ( .A1(G171), .A2(n750), .ZN(n743) );
  XNOR2_X1 U842 ( .A(KEYINPUT95), .B(n743), .ZN(n744) );
  NOR2_X1 U843 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U844 ( .A(n746), .B(KEYINPUT99), .ZN(n755) );
  NOR2_X1 U845 ( .A1(G2084), .A2(n757), .ZN(n771) );
  NAND2_X1 U846 ( .A1(G8), .A2(n757), .ZN(n801) );
  NOR2_X1 U847 ( .A1(G1966), .A2(n801), .ZN(n769) );
  NOR2_X1 U848 ( .A1(n771), .A2(n769), .ZN(n747) );
  NAND2_X1 U849 ( .A1(G8), .A2(n747), .ZN(n748) );
  XNOR2_X1 U850 ( .A(KEYINPUT30), .B(n748), .ZN(n749) );
  NOR2_X1 U851 ( .A1(G168), .A2(n749), .ZN(n752) );
  NOR2_X1 U852 ( .A1(G171), .A2(n750), .ZN(n751) );
  NOR2_X1 U853 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U854 ( .A(KEYINPUT31), .B(n753), .Z(n754) );
  NAND2_X1 U855 ( .A1(n755), .A2(n754), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n767), .A2(G286), .ZN(n756) );
  XOR2_X1 U857 ( .A(KEYINPUT101), .B(n756), .Z(n763) );
  NOR2_X1 U858 ( .A1(G1971), .A2(n801), .ZN(n759) );
  NOR2_X1 U859 ( .A1(G2090), .A2(n757), .ZN(n758) );
  NOR2_X1 U860 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U861 ( .A1(n760), .A2(G303), .ZN(n761) );
  XNOR2_X1 U862 ( .A(KEYINPUT102), .B(n761), .ZN(n762) );
  NAND2_X1 U863 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U864 ( .A1(n764), .A2(G8), .ZN(n766) );
  XOR2_X1 U865 ( .A(KEYINPUT103), .B(KEYINPUT32), .Z(n765) );
  XNOR2_X1 U866 ( .A(n766), .B(n765), .ZN(n796) );
  INV_X1 U867 ( .A(n767), .ZN(n768) );
  NOR2_X1 U868 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U869 ( .A(n770), .B(KEYINPUT100), .ZN(n773) );
  NAND2_X1 U870 ( .A1(n771), .A2(G8), .ZN(n772) );
  NAND2_X1 U871 ( .A1(n773), .A2(n772), .ZN(n795) );
  NAND2_X1 U872 ( .A1(G288), .A2(G1976), .ZN(n774) );
  XOR2_X1 U873 ( .A(KEYINPUT105), .B(n774), .Z(n957) );
  AND2_X1 U874 ( .A1(n795), .A2(n957), .ZN(n775) );
  NAND2_X1 U875 ( .A1(n796), .A2(n775), .ZN(n781) );
  INV_X1 U876 ( .A(n957), .ZN(n779) );
  NOR2_X1 U877 ( .A1(G1976), .A2(G288), .ZN(n945) );
  NOR2_X1 U878 ( .A1(G1971), .A2(G303), .ZN(n776) );
  NOR2_X1 U879 ( .A1(n945), .A2(n776), .ZN(n777) );
  XNOR2_X1 U880 ( .A(n777), .B(KEYINPUT104), .ZN(n778) );
  OR2_X1 U881 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U882 ( .A1(n781), .A2(n780), .ZN(n783) );
  AND2_X1 U883 ( .A1(n783), .A2(n782), .ZN(n784) );
  OR2_X1 U884 ( .A1(KEYINPUT33), .A2(n784), .ZN(n790) );
  NAND2_X1 U885 ( .A1(n945), .A2(KEYINPUT33), .ZN(n785) );
  NOR2_X1 U886 ( .A1(n785), .A2(n801), .ZN(n788) );
  XOR2_X1 U887 ( .A(G1981), .B(KEYINPUT106), .Z(n786) );
  XNOR2_X1 U888 ( .A(G305), .B(n786), .ZN(n942) );
  INV_X1 U889 ( .A(n942), .ZN(n787) );
  NOR2_X1 U890 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U891 ( .A1(n790), .A2(n789), .ZN(n806) );
  XNOR2_X1 U892 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n791) );
  XNOR2_X1 U893 ( .A(n791), .B(KEYINPUT92), .ZN(n793) );
  NOR2_X1 U894 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XNOR2_X1 U895 ( .A(n793), .B(n792), .ZN(n794) );
  OR2_X1 U896 ( .A1(n801), .A2(n794), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n796), .A2(n795), .ZN(n800) );
  NOR2_X1 U898 ( .A1(G2090), .A2(G303), .ZN(n797) );
  NAND2_X1 U899 ( .A1(G8), .A2(n797), .ZN(n798) );
  XOR2_X1 U900 ( .A(KEYINPUT107), .B(n798), .Z(n799) );
  NAND2_X1 U901 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U902 ( .A1(n802), .A2(n801), .ZN(n803) );
  AND2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n805) );
  AND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n811) );
  XNOR2_X1 U906 ( .A(G1986), .B(KEYINPUT86), .ZN(n809) );
  XNOR2_X1 U907 ( .A(n809), .B(G290), .ZN(n966) );
  NAND2_X1 U908 ( .A1(n966), .A2(n823), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n826) );
  AND2_X1 U910 ( .A1(n812), .A2(n878), .ZN(n922) );
  AND2_X1 U911 ( .A1(n994), .A2(n882), .ZN(n930) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U913 ( .A1(n930), .A2(n813), .ZN(n814) );
  NOR2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n922), .A2(n816), .ZN(n817) );
  XNOR2_X1 U916 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n820), .B(KEYINPUT108), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n879), .A2(n821), .ZN(n926) );
  NAND2_X1 U920 ( .A1(n822), .A2(n926), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n827), .ZN(G329) );
  XOR2_X1 U924 ( .A(G2454), .B(G2430), .Z(n829) );
  XNOR2_X1 U925 ( .A(G2451), .B(G2446), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n836) );
  XOR2_X1 U927 ( .A(G2443), .B(G2427), .Z(n831) );
  XNOR2_X1 U928 ( .A(G2438), .B(KEYINPUT109), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U930 ( .A(n832), .B(G2435), .Z(n834) );
  XNOR2_X1 U931 ( .A(G1341), .B(G1348), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n837), .A2(G14), .ZN(n909) );
  XOR2_X1 U935 ( .A(KEYINPUT110), .B(n909), .Z(G401) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U938 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U947 ( .A(KEYINPUT111), .B(n844), .ZN(G319) );
  XOR2_X1 U948 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U950 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U951 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U953 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U954 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U955 ( .A(G2084), .B(G2078), .ZN(n851) );
  XNOR2_X1 U956 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U957 ( .A(G1976), .B(G1981), .Z(n854) );
  XNOR2_X1 U958 ( .A(G1966), .B(G1971), .ZN(n853) );
  XNOR2_X1 U959 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U960 ( .A(n855), .B(G2474), .Z(n857) );
  XNOR2_X1 U961 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U962 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT41), .B(G1956), .Z(n859) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1961), .ZN(n858) );
  XNOR2_X1 U965 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U967 ( .A1(n893), .A2(G100), .ZN(n862) );
  XNOR2_X1 U968 ( .A(n862), .B(KEYINPUT112), .ZN(n864) );
  NAND2_X1 U969 ( .A1(G112), .A2(n890), .ZN(n863) );
  NAND2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U971 ( .A(n865), .B(KEYINPUT113), .ZN(n867) );
  NAND2_X1 U972 ( .A1(G136), .A2(n894), .ZN(n866) );
  NAND2_X1 U973 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n889), .A2(G124), .ZN(n868) );
  XOR2_X1 U975 ( .A(KEYINPUT44), .B(n868), .Z(n869) );
  NOR2_X1 U976 ( .A1(n870), .A2(n869), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G103), .A2(n893), .ZN(n872) );
  NAND2_X1 U978 ( .A1(G139), .A2(n894), .ZN(n871) );
  NAND2_X1 U979 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G127), .A2(n889), .ZN(n874) );
  NAND2_X1 U981 ( .A1(G115), .A2(n890), .ZN(n873) );
  NAND2_X1 U982 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U984 ( .A1(n877), .A2(n876), .ZN(n916) );
  XNOR2_X1 U985 ( .A(n916), .B(G162), .ZN(n881) );
  XNOR2_X1 U986 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U987 ( .A(n881), .B(n880), .ZN(n886) );
  XOR2_X1 U988 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n884) );
  XNOR2_X1 U989 ( .A(n882), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U990 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U991 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U992 ( .A(G164), .B(G160), .ZN(n887) );
  XNOR2_X1 U993 ( .A(n888), .B(n887), .ZN(n902) );
  NAND2_X1 U994 ( .A1(G130), .A2(n889), .ZN(n892) );
  NAND2_X1 U995 ( .A1(G118), .A2(n890), .ZN(n891) );
  NAND2_X1 U996 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G106), .A2(n893), .ZN(n896) );
  NAND2_X1 U998 ( .A1(G142), .A2(n894), .ZN(n895) );
  NAND2_X1 U999 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U1000 ( .A(KEYINPUT45), .B(n897), .Z(n898) );
  NOR2_X1 U1001 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1002 ( .A(n932), .B(n900), .Z(n901) );
  XNOR2_X1 U1003 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U1005 ( .A(n948), .B(n904), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(G171), .B(n956), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n907), .B(G286), .ZN(n908) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n908), .ZN(G397) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n909), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n910) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  XNOR2_X1 U1013 ( .A(n911), .B(KEYINPUT115), .ZN(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1019 ( .A(G164), .B(G2078), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(G2072), .B(n916), .ZN(n917) );
  XNOR2_X1 U1021 ( .A(n917), .B(KEYINPUT116), .ZN(n918) );
  NAND2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(n920), .B(KEYINPUT50), .ZN(n938) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1025 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n923), .Z(n936) );
  INV_X1 U1027 ( .A(n924), .ZN(n925) );
  NAND2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G160), .B(G2084), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n1014) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n1014), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n941), .A2(G29), .ZN(n1024) );
  XOR2_X1 U1040 ( .A(KEYINPUT56), .B(G16), .Z(n968) );
  XNOR2_X1 U1041 ( .A(G168), .B(G1966), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(n944), .B(KEYINPUT57), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(n945), .B(KEYINPUT123), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(G171), .B(G1961), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G1341), .B(n948), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G303), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT124), .B(n953), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n964) );
  XNOR2_X1 U1053 ( .A(n956), .B(G1348), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n962) );
  XOR2_X1 U1055 ( .A(G1956), .B(n959), .Z(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT122), .B(n960), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n1021) );
  XOR2_X1 U1061 ( .A(G1986), .B(G24), .Z(n970) );
  XOR2_X1 U1062 ( .A(G1971), .B(G22), .Z(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1066 ( .A(KEYINPUT58), .B(n973), .Z(n990) );
  XNOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT59), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n974), .B(G4), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G20), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(G1981), .B(G6), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1073 ( .A(KEYINPUT125), .B(G1341), .Z(n979) );
  XNOR2_X1 U1074 ( .A(G19), .B(n979), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT60), .B(n982), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n983), .B(G5), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(G21), .B(G1966), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1081 ( .A(KEYINPUT126), .B(n988), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT61), .B(n991), .Z(n992) );
  NOR2_X1 U1084 ( .A1(G16), .A2(n992), .ZN(n1018) );
  XNOR2_X1 U1085 ( .A(G2084), .B(G34), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(KEYINPUT54), .ZN(n1013) );
  XOR2_X1 U1087 ( .A(G2090), .B(G35), .Z(n1010) );
  XNOR2_X1 U1088 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n1007) );
  XNOR2_X1 U1089 ( .A(n994), .B(G25), .ZN(n995) );
  NAND2_X1 U1090 ( .A1(n995), .A2(G28), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(n996), .B(KEYINPUT118), .ZN(n1005) );
  XOR2_X1 U1092 ( .A(n997), .B(G27), .Z(n999) );
  XNOR2_X1 U1093 ( .A(G32), .B(G1996), .ZN(n998) );
  NOR2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(G2067), .B(G26), .ZN(n1001) );
  XNOR2_X1 U1096 ( .A(G33), .B(G2072), .ZN(n1000) );
  NOR2_X1 U1097 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1098 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1100 ( .A(n1007), .B(n1006), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(n1008), .B(KEYINPUT53), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1103 ( .A(KEYINPUT121), .B(n1011), .Z(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1015), .B(n1014), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(G29), .A2(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(G11), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1022), .Z(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

