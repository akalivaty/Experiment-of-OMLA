//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n593, new_n595, new_n596,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n639, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(G137), .A3(new_n460), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n474));
  INV_X1    g049(.A(G124), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n463), .A2(KEYINPUT67), .A3(new_n464), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(G2105), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n477), .A2(new_n460), .A3(new_n478), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT68), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n477), .A2(new_n482), .A3(new_n460), .A4(new_n478), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n487));
  OAI221_X1 g062(.A(new_n474), .B1(new_n475), .B2(new_n479), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(KEYINPUT70), .A2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT70), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n464), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n460), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .A4(new_n460), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n493), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  AND3_X1   g077(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT5), .B1(KEYINPUT75), .B2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT76), .A3(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT76), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT71), .B(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n521), .B(G651), .C1(new_n516), .C2(new_n517), .ZN(new_n522));
  AND4_X1   g097(.A1(new_n506), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n519), .A2(G543), .A3(new_n520), .A4(new_n522), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT74), .B1(new_n526), .B2(G50), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  NOR3_X1   g104(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n515), .B(new_n524), .C1(new_n527), .C2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n535), .B1(new_n503), .B2(new_n504), .ZN(new_n536));
  NAND2_X1  g111(.A1(KEYINPUT75), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT5), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(KEYINPUT77), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n542), .A2(G63), .A3(G651), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n519), .A2(new_n506), .A3(new_n520), .A4(new_n522), .ZN(new_n547));
  INV_X1    g122(.A(G89), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT78), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n551), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n544), .B1(new_n550), .B2(new_n552), .ZN(G168));
  NAND2_X1  g128(.A1(new_n542), .A2(G64), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n513), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n557), .A2(new_n525), .B1(new_n547), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT79), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n561));
  OAI221_X1 g136(.A(new_n561), .B1(new_n525), .B2(new_n557), .C1(new_n558), .C2(new_n547), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n556), .B1(new_n560), .B2(new_n562), .ZN(G171));
  NAND2_X1  g138(.A1(new_n526), .A2(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n523), .A2(G81), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n536), .B2(new_n541), .ZN(new_n567));
  AND2_X1   g142(.A1(G68), .A2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n514), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n564), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  AND3_X1   g147(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G36), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(G188));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G65), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n505), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(G91), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n547), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  INV_X1    g160(.A(G53), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n525), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR4_X1   g164(.A1(new_n525), .A2(KEYINPUT80), .A3(KEYINPUT9), .A4(new_n586), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n584), .B1(new_n589), .B2(new_n590), .ZN(G299));
  NAND2_X1  g166(.A1(new_n560), .A2(new_n562), .ZN(new_n592));
  INV_X1    g167(.A(new_n556), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G301));
  NAND2_X1  g169(.A1(new_n550), .A2(new_n552), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n534), .A2(new_n543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G286));
  OAI21_X1  g172(.A(G651), .B1(new_n542), .B2(G74), .ZN(new_n598));
  INV_X1    g173(.A(G87), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n547), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G49), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n525), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G288));
  INV_X1    g179(.A(G61), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n505), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(G73), .A2(G543), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n514), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G86), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n547), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G48), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n525), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n613));
  OR3_X1    g188(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n610), .B2(new_n612), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(G305));
  XNOR2_X1  g191(.A(KEYINPUT82), .B(G47), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n525), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n523), .A2(G85), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n542), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n618), .B(new_n619), .C1(new_n513), .C2(new_n620), .ZN(G290));
  INV_X1    g196(.A(G54), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n525), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  AND2_X1   g199(.A1(G79), .A2(G543), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n506), .B2(G66), .ZN(new_n626));
  INV_X1    g201(.A(G651), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(KEYINPUT10), .B1(new_n523), .B2(G92), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n631));
  INV_X1    g206(.A(G92), .ZN(new_n632));
  NOR3_X1   g207(.A1(new_n547), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n624), .B(new_n629), .C1(new_n630), .C2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(G171), .ZN(G284));
  OAI21_X1  g212(.A(new_n636), .B1(new_n635), .B2(G171), .ZN(G321));
  NAND2_X1  g213(.A1(G299), .A2(new_n635), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n635), .B2(G168), .ZN(G297));
  OAI21_X1  g215(.A(new_n639), .B1(new_n635), .B2(G168), .ZN(G280));
  AND3_X1   g216(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n642), .A2(KEYINPUT10), .A3(G92), .A4(new_n506), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n631), .B1(new_n547), .B2(new_n632), .ZN(new_n644));
  AOI211_X1 g219(.A(new_n628), .B(new_n623), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G860), .ZN(G148));
  NAND2_X1  g222(.A1(new_n570), .A2(new_n635), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n634), .A2(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(new_n635), .ZN(G323));
  XNOR2_X1  g225(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g226(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT83), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT13), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  INV_X1    g232(.A(G123), .ZN(new_n658));
  NOR2_X1   g233(.A1(G99), .A2(G2105), .ZN(new_n659));
  OAI21_X1  g234(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n660));
  OAI22_X1  g235(.A1(new_n479), .A2(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n484), .B2(G135), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2096), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n657), .A2(new_n663), .ZN(G156));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2430), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2435), .ZN(new_n666));
  XOR2_X1   g241(.A(G2427), .B(G2438), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT14), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2443), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT85), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1341), .B(G1348), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n670), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT86), .B(G2446), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  AND2_X1   g253(.A1(new_n678), .A2(G14), .ZN(G401));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2067), .B(G2678), .Z(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n680), .B1(new_n684), .B2(KEYINPUT18), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n687), .A3(KEYINPUT17), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT18), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2096), .B(G2100), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n695), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n699), .A2(KEYINPUT20), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n701), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n703), .A2(new_n695), .A3(new_n698), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n702), .B(new_n704), .C1(KEYINPUT20), .C2(new_n699), .ZN(new_n705));
  XOR2_X1   g280(.A(G1991), .B(G1996), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT88), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(G229));
  INV_X1    g287(.A(G26), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(G29), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n484), .A2(G140), .ZN(new_n715));
  INV_X1    g290(.A(G128), .ZN(new_n716));
  NOR2_X1   g291(.A1(G104), .A2(G2105), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n718));
  OAI22_X1  g293(.A1(new_n479), .A2(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n714), .B1(new_n721), .B2(G29), .ZN(new_n722));
  MUX2_X1   g297(.A(new_n714), .B(new_n722), .S(KEYINPUT28), .Z(new_n723));
  INV_X1    g298(.A(G2067), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G5), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G171), .B2(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G1961), .ZN(new_n728));
  NOR2_X1   g303(.A1(G16), .A2(G21), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G168), .B2(G16), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n728), .B1(G1966), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G19), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n571), .B2(new_n732), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  INV_X1    g310(.A(G28), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(KEYINPUT30), .B2(new_n736), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT24), .B(G34), .ZN(new_n739));
  MUX2_X1   g314(.A(new_n739), .B(G160), .S(G29), .Z(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G29), .B2(new_n662), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT94), .ZN(new_n744));
  INV_X1    g319(.A(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G29), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(G29), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n501), .B2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n746), .B1(new_n748), .B2(new_n744), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT95), .B(G2078), .Z(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n743), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G32), .ZN(new_n754));
  INV_X1    g329(.A(G141), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n481), .B2(new_n483), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT26), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n759));
  INV_X1    g334(.A(G129), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n479), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n756), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n754), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT27), .B(G1996), .Z(new_n764));
  OAI211_X1 g339(.A(new_n735), .B(new_n753), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  OR3_X1    g340(.A1(new_n725), .A2(new_n731), .A3(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G35), .B(new_n488), .S(G29), .Z(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT29), .B(G2090), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n767), .B(new_n768), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n732), .A2(G20), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n642), .A2(new_n588), .A3(G53), .A4(G543), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(KEYINPUT9), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n587), .A2(new_n588), .A3(new_n585), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n583), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g349(.A(KEYINPUT23), .B(new_n770), .C1(new_n774), .C2(new_n732), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(KEYINPUT23), .B2(new_n770), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1956), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n769), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G33), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n465), .A2(G127), .ZN(new_n780));
  NAND2_X1  g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n460), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n484), .B2(G139), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT25), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n779), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G2072), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n732), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n645), .B2(new_n732), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n730), .A2(G1966), .B1(new_n793), .B2(G1348), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n791), .B(new_n794), .C1(G1348), .C2(new_n793), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n740), .A2(new_n741), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n763), .A2(new_n764), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n798), .B1(new_n796), .B2(new_n797), .C1(G1961), .C2(new_n727), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT93), .Z(new_n800));
  NOR4_X1   g375(.A1(new_n766), .A2(new_n778), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n732), .A2(G6), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G305), .B2(G16), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT32), .B(G1981), .Z(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n732), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n732), .ZN(new_n808));
  INV_X1    g383(.A(G1971), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n732), .A2(G23), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n603), .B2(new_n732), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1976), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  OR3_X1    g391(.A1(new_n806), .A2(new_n816), .A3(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(G290), .A2(G16), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n732), .A2(G24), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G1986), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(KEYINPUT34), .B1(new_n806), .B2(new_n816), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n484), .A2(G131), .ZN(new_n824));
  INV_X1    g399(.A(G119), .ZN(new_n825));
  NOR2_X1   g400(.A1(G95), .A2(G2105), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(new_n460), .B2(G107), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n479), .A2(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G25), .B(new_n830), .S(G29), .Z(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n820), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(G1986), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n817), .A2(new_n822), .A3(new_n823), .A4(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT90), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT31), .B(G11), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n837), .A2(KEYINPUT90), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n801), .A2(new_n839), .A3(new_n840), .A4(new_n842), .ZN(G150));
  INV_X1    g418(.A(G150), .ZN(G311));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n568), .B1(new_n542), .B2(G56), .ZN(new_n846));
  INV_X1    g421(.A(G43), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n846), .A2(new_n513), .B1(new_n525), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G81), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n547), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n845), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT98), .A4(new_n569), .ZN(new_n852));
  AND2_X1   g427(.A1(G80), .A2(G543), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n542), .B2(G67), .ZN(new_n854));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n854), .A2(new_n513), .B1(new_n525), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT97), .B(G93), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n547), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n851), .A2(new_n852), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G67), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n536), .B2(new_n541), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n514), .B1(new_n862), .B2(new_n853), .ZN(new_n863));
  OAI221_X1 g438(.A(new_n863), .B1(new_n855), .B2(new_n525), .C1(new_n547), .C2(new_n857), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n570), .A2(new_n864), .A3(new_n845), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n645), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT39), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n868), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT99), .B(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT100), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n859), .A2(new_n872), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G145));
  XNOR2_X1  g452(.A(new_n662), .B(G160), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n756), .A2(new_n758), .A3(new_n761), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT101), .ZN(new_n881));
  NOR4_X1   g456(.A1(new_n756), .A2(KEYINPUT101), .A3(new_n761), .A4(new_n758), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n721), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n762), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n720), .B1(new_n886), .B2(new_n882), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n884), .A2(new_n887), .A3(G164), .ZN(new_n888));
  AOI21_X1  g463(.A(G164), .B1(new_n884), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n787), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n721), .B1(new_n881), .B2(new_n883), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n886), .A2(new_n882), .A3(new_n720), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n501), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n884), .A2(new_n887), .A3(G164), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n789), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n890), .A2(new_n488), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n488), .B1(new_n890), .B2(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(G130), .ZN(new_n898));
  NOR2_X1   g473(.A1(G106), .A2(G2105), .ZN(new_n899));
  OAI21_X1  g474(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n900));
  OAI22_X1  g475(.A1(new_n479), .A2(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n484), .B2(G142), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n829), .B(new_n902), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n655), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n896), .A2(new_n897), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n789), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n888), .A2(new_n889), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n787), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n893), .B2(new_n894), .ZN(new_n910));
  OAI21_X1  g485(.A(G162), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n890), .A2(new_n488), .A3(new_n895), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n904), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n879), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n905), .B1(new_n896), .B2(new_n897), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n904), .A3(new_n912), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n878), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g495(.A(G85), .ZN(new_n921));
  OAI22_X1  g496(.A1(new_n620), .A2(new_n513), .B1(new_n547), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n525), .A2(new_n617), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(G288), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G290), .A2(new_n603), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT104), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G305), .A2(G166), .ZN(new_n928));
  NAND3_X1  g503(.A1(G303), .A2(new_n614), .A3(new_n615), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n932));
  NOR2_X1   g507(.A1(G288), .A2(new_n924), .ZN(new_n933));
  NOR2_X1   g508(.A1(G290), .A2(new_n603), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT104), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n930), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n866), .B1(G559), .B2(new_n634), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n649), .A2(new_n865), .A3(new_n860), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G299), .A2(new_n645), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n772), .A2(new_n773), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n634), .A2(new_n945), .A3(new_n584), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n944), .A2(new_n946), .A3(KEYINPUT41), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT41), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI211_X1 g525(.A(KEYINPUT103), .B(KEYINPUT41), .C1(new_n944), .C2(new_n946), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n943), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n944), .A2(new_n946), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT102), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n955));
  NOR2_X1   g530(.A1(G299), .A2(new_n645), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n774), .A2(new_n634), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n942), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n939), .B1(new_n952), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT41), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n956), .B2(new_n957), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n944), .A2(new_n946), .A3(KEYINPUT41), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(KEYINPUT103), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n948), .A2(new_n949), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n942), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n954), .A2(new_n958), .B1(new_n941), .B2(new_n940), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n967), .A2(KEYINPUT42), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n938), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n947), .A2(new_n948), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n951), .B1(new_n971), .B2(KEYINPUT103), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n939), .B(new_n960), .C1(new_n972), .C2(new_n942), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT42), .B1(new_n967), .B2(new_n968), .ZN(new_n974));
  INV_X1    g549(.A(new_n938), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(G868), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n864), .A2(new_n635), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT105), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(new_n977), .ZN(G295));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n983));
  INV_X1    g558(.A(new_n979), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n975), .B1(new_n973), .B2(new_n974), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n984), .B1(new_n987), .B2(G868), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n977), .A2(new_n981), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n983), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n980), .B(KEYINPUT106), .C1(new_n981), .C2(new_n977), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(G331));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n860), .A2(new_n865), .ZN(new_n994));
  NOR2_X1   g569(.A1(G301), .A2(G168), .ZN(new_n995));
  NOR2_X1   g570(.A1(G171), .A2(G286), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n998));
  NAND2_X1  g573(.A1(G301), .A2(G168), .ZN(new_n999));
  NAND2_X1  g574(.A1(G171), .A2(G286), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n866), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n994), .B(KEYINPUT107), .C1(new_n995), .C2(new_n996), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n953), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n997), .A2(new_n1001), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n972), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1008), .A3(new_n975), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n963), .A2(new_n964), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1002), .A2(new_n1010), .A3(new_n1003), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n954), .A2(new_n997), .A3(new_n958), .A4(new_n1001), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n938), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT108), .B(new_n930), .C1(new_n931), .C2(new_n937), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1009), .A2(new_n1018), .A3(new_n915), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1009), .A2(new_n1018), .A3(KEYINPUT110), .A4(new_n915), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n993), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1007), .A2(new_n966), .A3(new_n965), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n953), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(G37), .B1(new_n1026), .B2(new_n975), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1017), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT43), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT44), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT109), .B1(new_n1019), .B2(KEYINPUT43), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1009), .A3(new_n915), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT43), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1027), .A2(new_n1034), .A3(new_n993), .A4(new_n1018), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1030), .A2(new_n1038), .ZN(G397));
  INV_X1    g614(.A(G1384), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n501), .A2(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(KEYINPUT111), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(KEYINPUT111), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1042), .A2(new_n1043), .A3(KEYINPUT45), .ZN(new_n1044));
  INV_X1    g619(.A(G40), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n468), .A2(new_n471), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OR3_X1    g622(.A1(new_n1047), .A2(KEYINPUT113), .A3(G1996), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT113), .B1(new_n1047), .B2(G1996), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n762), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n720), .B(new_n724), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1047), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(G1996), .A3(new_n880), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1051), .A2(new_n1058), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n830), .A2(new_n832), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n830), .A2(new_n832), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1053), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G290), .A2(G1986), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n924), .A2(new_n821), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(KEYINPUT112), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1053), .B(new_n1065), .C1(KEYINPUT112), .C2(new_n1063), .ZN(new_n1066));
  AND4_X1   g641(.A1(new_n1057), .A2(new_n1059), .A3(new_n1062), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G299), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n945), .A2(KEYINPUT57), .A3(new_n584), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1040), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1046), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT45), .B1(new_n501), .B2(new_n1040), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n501), .A2(KEYINPUT50), .A3(new_n1040), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT50), .B1(new_n501), .B2(new_n1040), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1046), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT118), .B(G1956), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1076), .A2(new_n1077), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1072), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1072), .B2(new_n1083), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1072), .A2(new_n1083), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1068), .B1(new_n1088), .B2(KEYINPUT61), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT121), .B(G1341), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT58), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1046), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1041), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT122), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1075), .ZN(new_n1095));
  INV_X1    g670(.A(G1996), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1046), .A4(new_n1073), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(new_n1091), .C1(new_n1092), .C2(new_n1041), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1094), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n571), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1103), .A3(new_n571), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1092), .A2(new_n1041), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n724), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1079), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n501), .A2(KEYINPUT50), .A3(new_n1040), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1092), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1107), .B1(new_n1110), .B2(G1348), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n645), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1107), .B(new_n634), .C1(new_n1110), .C2(G1348), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT60), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1072), .A2(new_n1083), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1095), .A2(new_n1046), .A3(new_n1073), .A4(new_n1077), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1110), .B2(new_n1081), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1116), .A2(new_n1119), .A3(KEYINPUT61), .ZN(new_n1120));
  OR3_X1    g695(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n634), .ZN(new_n1121));
  AND4_X1   g696(.A1(new_n1105), .A2(new_n1115), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1086), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1072), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT123), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1089), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1119), .A2(new_n1112), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1123), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT120), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1128), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1129), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1076), .A2(G1966), .B1(new_n1080), .B2(G2084), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1135), .A2(G8), .A3(G286), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(G8), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n1138));
  INV_X1    g713(.A(G8), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1137), .B(new_n1138), .C1(new_n1139), .C2(G168), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT51), .B(G8), .C1(new_n1135), .C2(G286), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OR3_X1    g717(.A1(new_n1074), .A2(G2078), .A3(new_n1075), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n1144));
  INV_X1    g719(.A(G1961), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1143), .A2(new_n1144), .B1(new_n1145), .B2(new_n1080), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1144), .B2(new_n1143), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G301), .B(KEYINPUT54), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1142), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1148), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT125), .B(G2078), .Z(new_n1151));
  OR4_X1    g726(.A1(new_n1144), .A2(new_n1044), .A3(new_n1074), .A4(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n1154));
  NAND3_X1  g729(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT115), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT55), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(G166), .B2(new_n1139), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT115), .ZN(new_n1159));
  NAND4_X1  g734(.A1(G303), .A2(new_n1159), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT116), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT116), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1156), .A2(new_n1158), .A3(new_n1163), .A4(new_n1160), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1076), .A2(G1971), .B1(new_n1080), .B2(G2090), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(G8), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1167), .A2(new_n1158), .A3(new_n1156), .A4(new_n1160), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  OR3_X1    g746(.A1(new_n610), .A2(new_n612), .A3(G1981), .ZN(new_n1172));
  OAI21_X1  g747(.A(G1981), .B1(new_n610), .B2(new_n612), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT49), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1106), .A2(new_n1139), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(KEYINPUT49), .A3(new_n1173), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n603), .A2(G1976), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT52), .ZN(new_n1182));
  XOR2_X1   g757(.A(KEYINPUT117), .B(G1976), .Z(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT52), .B1(G288), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1179), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1171), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1154), .B1(new_n1169), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1167), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1170), .A2(new_n1179), .A3(new_n1182), .A4(new_n1185), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1189), .A2(new_n1190), .A3(KEYINPUT126), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1149), .B(new_n1153), .C1(new_n1188), .C2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1133), .A2(new_n1134), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1142), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(G171), .B1(new_n1142), .B2(new_n1194), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1197), .B(new_n1147), .C1(new_n1188), .C2(new_n1191), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1137), .A2(G286), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1169), .A2(new_n1187), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT63), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1186), .ZN(new_n1203));
  INV_X1    g778(.A(G1976), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1179), .A2(new_n1204), .A3(new_n603), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1172), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1189), .A2(new_n1203), .B1(new_n1177), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1198), .A2(new_n1202), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1067), .B1(new_n1193), .B2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1050), .B(KEYINPUT46), .Z(new_n1210));
  OAI21_X1  g785(.A(new_n1053), .B1(new_n1052), .B2(new_n880), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT127), .Z(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT47), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1213), .B(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n720), .A2(new_n724), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1047), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1047), .A2(new_n1064), .ZN(new_n1219));
  XOR2_X1   g794(.A(new_n1219), .B(KEYINPUT48), .Z(new_n1220));
  AND4_X1   g795(.A1(new_n1057), .A2(new_n1059), .A3(new_n1062), .A4(new_n1220), .ZN(new_n1221));
  NOR3_X1   g796(.A1(new_n1215), .A2(new_n1218), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1209), .A2(new_n1222), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g798(.A1(G227), .A2(new_n458), .ZN(new_n1225));
  NOR2_X1   g799(.A1(G401), .A2(G229), .ZN(new_n1226));
  AND4_X1   g800(.A1(new_n919), .A2(new_n1036), .A3(new_n1225), .A4(new_n1226), .ZN(G308));
  NAND4_X1  g801(.A1(new_n1036), .A2(new_n919), .A3(new_n1225), .A4(new_n1226), .ZN(G225));
endmodule


