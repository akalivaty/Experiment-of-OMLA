//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0007(.A(G97), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n215), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  OR3_X1    g0023(.A1(new_n215), .A2(KEYINPUT65), .A3(G13), .ZN(new_n224));
  OAI21_X1  g0024(.A(KEYINPUT65), .B1(new_n215), .B2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n213), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n206), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n223), .B(new_n228), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n237), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  OAI21_X1  g0050(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G150), .ZN(new_n253));
  XOR2_X1   g0053(.A(KEYINPUT8), .B(G58), .Z(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n213), .A2(G33), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n251), .B(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n229), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n213), .A2(G1), .ZN(new_n261));
  INV_X1    g0061(.A(G50), .ZN(new_n262));
  OR3_X1    g0062(.A1(new_n261), .A2(KEYINPUT69), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n259), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT69), .B1(new_n261), .B2(new_n262), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G50), .B2(new_n264), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n270), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n260), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n277), .A2(G274), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n229), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n277), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n280), .B1(G226), .B2(new_n283), .ZN(new_n284));
  XOR2_X1   g0084(.A(new_n284), .B(KEYINPUT67), .Z(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  INV_X1    g0088(.A(G77), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n286), .A2(G222), .A3(new_n292), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n291), .B1(new_n290), .B2(new_n293), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(new_n282), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n285), .A2(G190), .A3(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n260), .B(KEYINPUT9), .C1(new_n271), .C2(new_n272), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n275), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT10), .B1(new_n299), .B2(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n285), .A2(new_n296), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n299), .B(new_n302), .C1(KEYINPUT72), .C2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n273), .C1(G179), .C2(new_n301), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n252), .A2(G50), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT74), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n256), .A2(new_n289), .B1(new_n213), .B2(G68), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n259), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT11), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n317));
  OR3_X1    g0117(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n261), .A2(new_n202), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n317), .A2(new_n318), .B1(new_n266), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n315), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n280), .A2(KEYINPUT73), .B1(new_n283), .B2(G238), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n279), .A2(G274), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n276), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n286), .A2(G232), .A3(G1698), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n286), .A2(G226), .A3(new_n292), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n282), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n322), .A2(new_n325), .ZN(new_n334));
  INV_X1    g0134(.A(new_n332), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT13), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(G169), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(new_n336), .A3(G179), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n338), .B1(new_n337), .B2(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n321), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n337), .A2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(new_n321), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n333), .A2(new_n336), .A3(G190), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n259), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n254), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT15), .B(G87), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n350), .A2(new_n256), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n348), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n266), .ZN(new_n353));
  OAI21_X1  g0153(.A(G77), .B1(new_n213), .B2(G1), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n353), .A2(new_n354), .B1(G77), .B2(new_n264), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT71), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT71), .B1(new_n352), .B2(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G238), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n287), .A2(new_n361), .B1(new_n209), .B2(new_n286), .ZN(new_n362));
  INV_X1    g0162(.A(G33), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G33), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n367), .A2(new_n239), .A3(G1698), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n282), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n280), .B1(G244), .B2(new_n283), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n306), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n360), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n374), .A3(new_n370), .ZN(new_n375));
  INV_X1    g0175(.A(G200), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n369), .B2(new_n370), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n360), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n369), .A2(G190), .A3(new_n370), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n373), .A2(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n343), .A2(new_n347), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n309), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n255), .A2(new_n261), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n266), .B1(new_n255), .B2(new_n265), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G58), .A2(G68), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n203), .A2(new_n205), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(G20), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n252), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n388), .B2(G20), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n386), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(G20), .B1(new_n364), .B2(new_n366), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT75), .B1(new_n395), .B2(KEYINPUT7), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(KEYINPUT7), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(new_n286), .C2(G20), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G68), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n388), .A2(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT76), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n404), .A2(KEYINPUT77), .A3(new_n391), .A4(new_n390), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n394), .A2(new_n402), .A3(KEYINPUT16), .A4(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n406), .A2(new_n259), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT78), .B1(new_n395), .B2(KEYINPUT7), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT78), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n409), .B(new_n399), .C1(new_n286), .C2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n410), .A3(new_n397), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G68), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n394), .A2(new_n412), .A3(new_n405), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n385), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n286), .A2(G223), .A3(new_n292), .ZN(new_n417));
  INV_X1    g0217(.A(G87), .ZN(new_n418));
  INV_X1    g0218(.A(G226), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n417), .B1(new_n363), .B2(new_n418), .C1(new_n287), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n282), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n280), .B1(G232), .B2(new_n283), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n376), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g0223(.A1(KEYINPUT80), .A2(G190), .ZN(new_n424));
  NOR2_X1   g0224(.A1(KEYINPUT80), .A2(G190), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n421), .A2(new_n422), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n415), .A2(new_n259), .A3(new_n406), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(new_n384), .A3(new_n429), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n421), .A2(G179), .A3(new_n422), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n306), .B1(new_n421), .B2(new_n422), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI211_X1 g0238(.A(KEYINPUT18), .B(new_n438), .C1(new_n431), .C2(new_n384), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n413), .A2(new_n414), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n406), .A2(new_n259), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n384), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n438), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT79), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT18), .B1(new_n416), .B2(new_n438), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(new_n440), .A3(new_n444), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n435), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n382), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n364), .A2(new_n366), .A3(G244), .A4(new_n292), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT4), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT83), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(KEYINPUT83), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n460), .A2(KEYINPUT84), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n364), .A2(new_n366), .A3(G250), .A4(G1698), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n464), .C1(new_n453), .C2(new_n454), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n279), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G257), .A3(new_n279), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(G274), .A3(new_n279), .A4(new_n469), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT85), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT85), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n376), .B1(new_n467), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n453), .A2(KEYINPUT83), .A3(new_n454), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT83), .B1(new_n453), .B2(new_n454), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n282), .B1(new_n484), .B2(new_n465), .ZN(new_n485));
  INV_X1    g0285(.A(new_n479), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n478), .B1(new_n473), .B2(new_n475), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G190), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n264), .A2(new_n208), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n212), .A2(G33), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n264), .A2(new_n493), .A3(new_n229), .A4(new_n258), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n494), .B(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n492), .B1(new_n496), .B2(new_n208), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n252), .A2(G77), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n499), .A2(new_n208), .A3(G107), .ZN(new_n500));
  XNOR2_X1  g0300(.A(G97), .B(G107), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n502), .B2(new_n213), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n411), .B2(G107), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n497), .B1(new_n504), .B2(new_n348), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT82), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT82), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(new_n497), .C1(new_n504), .C2(new_n348), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n491), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT19), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n213), .B1(new_n330), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(G87), .B2(new_n210), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n364), .A2(new_n366), .A3(new_n213), .A4(G68), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n256), .B2(new_n208), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n259), .ZN(new_n516));
  XOR2_X1   g0316(.A(KEYINPUT15), .B(G87), .Z(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n264), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT86), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n516), .A2(KEYINPUT86), .A3(new_n519), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n523), .B1(G87), .B2(new_n496), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n279), .A2(G274), .A3(new_n469), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n212), .A2(G45), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(G250), .C1(new_n281), .C2(new_n229), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n364), .A2(new_n366), .A3(G244), .A4(G1698), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n364), .A2(new_n366), .A3(G238), .A4(new_n292), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n528), .B1(new_n532), .B2(new_n282), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n376), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(G190), .B2(new_n533), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n533), .A2(G169), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n374), .B2(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n496), .A2(new_n517), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT86), .B1(new_n516), .B2(new_n519), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n521), .B(new_n518), .C1(new_n515), .C2(new_n259), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n524), .A2(new_n535), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n467), .A2(new_n480), .A3(new_n374), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n306), .B1(new_n485), .B2(new_n488), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n505), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n509), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n364), .A2(new_n366), .A3(G257), .A4(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n364), .A2(new_n366), .A3(G250), .A4(new_n292), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n229), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n474), .A2(new_n469), .B1(new_n551), .B2(new_n278), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n550), .A2(new_n282), .B1(new_n552), .B2(G264), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n475), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n376), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G190), .B2(new_n554), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT90), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n364), .A2(new_n366), .A3(new_n213), .A4(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT22), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT22), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n286), .A2(new_n560), .A3(new_n213), .A4(G87), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n531), .A2(G20), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n213), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n209), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n562), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n563), .B1(new_n562), .B2(new_n568), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n259), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XOR2_X1   g0371(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n572));
  NOR2_X1   g0372(.A1(new_n264), .A2(G107), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT89), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n496), .A2(G107), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n556), .A2(new_n557), .A3(new_n571), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n571), .A2(new_n579), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n553), .A2(new_n489), .A3(new_n475), .ZN(new_n582));
  AOI21_X1  g0382(.A(G200), .B1(new_n553), .B2(new_n475), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT90), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n365), .A2(G33), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n588));
  OAI21_X1  g0388(.A(G303), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n364), .A2(new_n366), .A3(G264), .A4(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n364), .A2(new_n366), .A3(G257), .A4(new_n292), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n282), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(KEYINPUT87), .A3(new_n282), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  MUX2_X1   g0397(.A(new_n264), .B(new_n494), .S(G116), .Z(new_n598));
  OAI21_X1  g0398(.A(new_n213), .B1(new_n208), .B2(G33), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n463), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(G116), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n259), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT20), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n599), .B1(new_n461), .B2(new_n462), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n607), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n598), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n472), .A2(G270), .A3(new_n279), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n611), .A2(G179), .A3(new_n475), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n597), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(G169), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n475), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n595), .B2(new_n596), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT21), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n616), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n597), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n601), .A2(KEYINPUT20), .A3(new_n605), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n608), .B1(new_n607), .B2(new_n604), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n306), .B1(new_n624), .B2(new_n598), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n614), .B1(new_n618), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n597), .A2(new_n427), .A3(new_n619), .ZN(new_n628));
  INV_X1    g0428(.A(new_n610), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n628), .B(new_n629), .C1(new_n376), .C2(new_n617), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n554), .A2(new_n306), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n553), .A2(new_n374), .A3(new_n475), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n581), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n586), .A2(new_n627), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n452), .A2(new_n546), .A3(new_n634), .ZN(G372));
  NOR2_X1   g0435(.A1(new_n439), .A2(new_n445), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n435), .ZN(new_n638));
  INV_X1    g0438(.A(new_n347), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n373), .A2(new_n375), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n343), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n637), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n304), .A2(new_n305), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n308), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n543), .A2(new_n544), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n506), .A2(new_n508), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n536), .A2(KEYINPUT91), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n536), .A2(KEYINPUT91), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n533), .A2(new_n374), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n541), .B1(new_n524), .B2(new_n535), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT26), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n542), .A2(new_n646), .A3(new_n505), .ZN(new_n655));
  XOR2_X1   g0455(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n541), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n653), .A2(new_n586), .A3(new_n545), .A4(new_n509), .ZN(new_n660));
  INV_X1    g0460(.A(new_n627), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n581), .A2(new_n631), .A3(new_n632), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n659), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n645), .B1(new_n452), .B2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G213), .ZN(new_n667));
  INV_X1    g0467(.A(G13), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n668), .A2(G1), .A3(G20), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT27), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n669), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(KEYINPUT93), .A3(KEYINPUT27), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT93), .B1(new_n672), .B2(KEYINPUT27), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n581), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT95), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n662), .B1(new_n580), .B2(new_n585), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT96), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n662), .B2(new_n678), .ZN(new_n684));
  INV_X1    g0484(.A(new_n678), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n629), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n661), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n621), .B1(new_n620), .B2(new_n625), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n615), .A2(new_n617), .A3(KEYINPUT21), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n630), .B(new_n613), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n687), .B1(new_n690), .B2(new_n686), .ZN(new_n691));
  XNOR2_X1  g0491(.A(KEYINPUT94), .B(G330), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n684), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n662), .A2(new_n685), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n627), .A2(new_n678), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n683), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n226), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n418), .A2(new_n208), .A3(new_n209), .A4(new_n602), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n702), .A2(new_n212), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n232), .B2(new_n702), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  AND2_X1   g0506(.A1(new_n648), .A2(new_n653), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n707), .A2(KEYINPUT26), .B1(new_n655), .B2(new_n656), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n685), .B1(new_n708), .B2(new_n664), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n711), .B(new_n685), .C1(new_n658), .C2(new_n664), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n553), .A2(new_n612), .A3(new_n533), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n597), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n485), .A2(new_n488), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n467), .A2(new_n480), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(KEYINPUT30), .A3(new_n597), .A4(new_n715), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n533), .A2(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n620), .A2(new_n717), .A3(new_n554), .A4(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT31), .B1(new_n723), .B2(new_n678), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n509), .A2(new_n545), .A3(new_n542), .ZN(new_n727));
  INV_X1    g0527(.A(new_n690), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(new_n681), .A4(new_n685), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n693), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n713), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n706), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(new_n668), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n212), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n702), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n691), .B2(new_n693), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n693), .B2(new_n691), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n226), .A2(G355), .A3(new_n286), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G116), .B2(new_n226), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n226), .A2(new_n367), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n468), .B2(new_n232), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n246), .A2(new_n468), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n551), .B1(new_n213), .B2(G169), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n747), .A2(KEYINPUT97), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(KEYINPUT97), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n738), .B1(new_n746), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n376), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G20), .A3(G190), .ZN(new_n758));
  INV_X1    g0558(.A(G303), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n367), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n213), .A2(new_n374), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  INV_X1    g0565(.A(G294), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n213), .B1(new_n767), .B2(G190), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n213), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n757), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n760), .B(new_n769), .C1(G283), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n762), .A2(new_n426), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n213), .A2(new_n374), .A3(new_n376), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n427), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT98), .B(G326), .Z(new_n779));
  OAI22_X1  g0579(.A1(new_n775), .A2(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n777), .A2(new_n489), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G329), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n770), .A2(new_n767), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT99), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n773), .B(new_n784), .C1(new_n785), .C2(new_n787), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n764), .A2(new_n289), .B1(new_n202), .B2(new_n781), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G58), .B2(new_n774), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n286), .B1(new_n771), .B2(new_n209), .ZN(new_n791));
  INV_X1    g0591(.A(new_n758), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(G87), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  INV_X1    g0596(.A(new_n778), .ZN(new_n797));
  INV_X1    g0597(.A(new_n768), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n797), .A2(G50), .B1(G97), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n790), .A2(new_n793), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n788), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n756), .B1(new_n801), .B2(new_n750), .ZN(new_n802));
  INV_X1    g0602(.A(new_n753), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n691), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n740), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n665), .A2(new_n678), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n360), .A2(new_n678), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n360), .A2(new_n375), .A3(new_n372), .A4(new_n678), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n809), .A2(KEYINPUT102), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(KEYINPUT102), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n380), .A2(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n807), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n732), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT103), .ZN(new_n815));
  INV_X1    g0615(.A(new_n738), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n732), .C2(new_n813), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n750), .A2(new_n751), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(G77), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G143), .A2(new_n774), .B1(new_n782), .B2(G150), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n822), .B2(new_n778), .C1(new_n794), .C2(new_n764), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n758), .A2(new_n262), .B1(new_n771), .B2(new_n202), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G58), .B2(new_n798), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n286), .B1(new_n787), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT101), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n797), .A2(G303), .B1(G294), .B2(new_n774), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n781), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n764), .A2(new_n602), .B1(new_n208), .B2(new_n768), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n787), .A2(new_n765), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n367), .B1(new_n771), .B2(new_n418), .C1(new_n209), .C2(new_n758), .ZN(new_n838));
  OR3_X1    g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n829), .A2(new_n832), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n816), .B(new_n820), .C1(new_n840), .C2(new_n750), .ZN(new_n841));
  INV_X1    g0641(.A(new_n812), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n752), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n817), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  INV_X1    g0645(.A(new_n502), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT35), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT35), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(G116), .A3(new_n230), .A4(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT36), .Z(new_n850));
  NAND3_X1  g0650(.A1(new_n232), .A2(G77), .A3(new_n387), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(KEYINPUT104), .B1(new_n262), .B2(G68), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(KEYINPUT104), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n212), .A2(G13), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n735), .A2(new_n212), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n432), .B1(new_n416), .B2(new_n438), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n676), .B(KEYINPUT106), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n416), .A2(new_n860), .ZN(new_n861));
  OR3_X1    g0661(.A1(new_n858), .A2(new_n861), .A3(KEYINPUT37), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n394), .A2(new_n402), .A3(new_n405), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n414), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n385), .B1(new_n407), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n432), .B1(new_n865), .B2(new_n438), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n676), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n439), .A2(new_n445), .A3(KEYINPUT79), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n448), .B1(new_n447), .B2(new_n449), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n638), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT105), .B1(new_n872), .B2(new_n867), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  INV_X1    g0674(.A(new_n867), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n451), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT38), .B(new_n869), .C1(new_n873), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n416), .B(new_n860), .C1(new_n638), .C2(new_n636), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n858), .B2(new_n861), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n862), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT39), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n872), .A2(KEYINPUT105), .A3(new_n867), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n874), .B1(new_n451), .B2(new_n875), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n886), .B2(new_n869), .ZN(new_n887));
  INV_X1    g0687(.A(new_n869), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n878), .B(new_n888), .C1(new_n884), .C2(new_n885), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n883), .B1(new_n890), .B2(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n337), .A2(G169), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT14), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n340), .A3(new_n339), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n321), .A3(new_n685), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n869), .B1(new_n873), .B2(new_n876), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n878), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n877), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n321), .B(new_n678), .C1(new_n894), .C2(new_n639), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n321), .A2(new_n678), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n343), .A2(new_n347), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n685), .B(new_n842), .C1(new_n658), .C2(new_n664), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n373), .A2(new_n375), .A3(new_n685), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n900), .A2(new_n908), .B1(new_n637), .B2(new_n860), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n897), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n452), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT107), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n713), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n713), .B2(new_n911), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n645), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n910), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n726), .A2(new_n729), .A3(KEYINPUT108), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT108), .B1(new_n726), .B2(new_n729), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n812), .B1(new_n901), .B2(new_n903), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n918), .B1(new_n890), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n877), .A2(new_n882), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n923), .A2(new_n918), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n452), .A2(new_n920), .A3(new_n919), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n693), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n857), .B1(new_n917), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT109), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n932), .A2(new_n933), .B1(new_n917), .B2(new_n931), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n856), .B1(new_n934), .B2(new_n935), .ZN(G367));
  NOR2_X1   g0736(.A1(new_n524), .A2(new_n685), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n659), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n653), .B2(new_n937), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT110), .Z(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n648), .A2(new_n678), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n647), .A2(new_n678), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n545), .A3(new_n509), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n545), .B1(new_n947), .B2(new_n633), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n685), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n699), .A2(KEYINPUT111), .A3(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT111), .B1(new_n699), .B2(new_n947), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n950), .A2(KEYINPUT42), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT42), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n942), .B(new_n949), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT112), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n940), .B(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n696), .A2(new_n947), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n702), .B(KEYINPUT41), .Z(new_n966));
  XOR2_X1   g0766(.A(new_n694), .B(KEYINPUT113), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n694), .A2(KEYINPUT113), .ZN(new_n968));
  INV_X1    g0768(.A(new_n684), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n699), .B1(new_n969), .B2(new_n698), .ZN(new_n970));
  MUX2_X1   g0770(.A(new_n967), .B(new_n968), .S(new_n970), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n733), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n946), .B1(new_n699), .B2(new_n697), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT44), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n699), .A2(new_n697), .A3(new_n946), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n695), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n977), .A3(new_n696), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n972), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n966), .B1(new_n982), .B2(new_n733), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n964), .B(new_n965), .C1(new_n737), .C2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n237), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n754), .B1(new_n226), .B2(new_n350), .C1(new_n985), .C2(new_n743), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT114), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n816), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n987), .B2(new_n986), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n771), .A2(new_n289), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G58), .B2(new_n792), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n991), .B(new_n286), .C1(new_n822), .C2(new_n786), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n768), .A2(new_n202), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n774), .B2(G150), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n262), .B2(new_n764), .ZN(new_n995));
  INV_X1    g0795(.A(G143), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n778), .A2(new_n996), .B1(new_n794), .B2(new_n781), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n992), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT115), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n792), .A2(G116), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT46), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1000), .A2(new_n1001), .B1(new_n778), .B2(new_n765), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G283), .B2(new_n763), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1001), .A2(new_n1000), .B1(new_n774), .B2(G303), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n209), .B2(new_n768), .C1(new_n766), .C2(new_n781), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n772), .A2(G97), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n786), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(G317), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1008), .A3(new_n367), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n999), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT47), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1011), .A2(KEYINPUT47), .B1(new_n748), .B2(new_n749), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n989), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n941), .B2(new_n803), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n984), .A2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n684), .A2(new_n753), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G317), .A2(new_n774), .B1(new_n763), .B2(G303), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT116), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n778), .A2(new_n776), .B1(new_n765), .B2(new_n781), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT48), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT48), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n792), .A2(G294), .B1(new_n798), .B2(G283), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT49), .Z(new_n1027));
  OAI221_X1 g0827(.A(new_n367), .B1(new_n771), .B2(new_n602), .C1(new_n779), .C2(new_n786), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G50), .A2(new_n774), .B1(new_n782), .B2(new_n254), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n202), .B2(new_n764), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n792), .A2(G77), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1007), .A2(G150), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1032), .A2(new_n1006), .A3(new_n1033), .A4(new_n286), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n778), .A2(new_n794), .B1(new_n350), .B2(new_n768), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n750), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n242), .A2(new_n468), .A3(new_n286), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n255), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT50), .B1(new_n255), .B2(G50), .ZN(new_n1040));
  AOI21_X1  g0840(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n703), .B1(new_n1042), .B2(new_n367), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n226), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n755), .B1(G107), .B2(new_n701), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n816), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1037), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT117), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n971), .A2(new_n737), .B1(new_n1017), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n972), .A2(new_n702), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n971), .A2(new_n733), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n972), .A2(new_n981), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n982), .A2(new_n702), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n736), .B1(new_n981), .B2(KEYINPUT118), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(KEYINPUT118), .B2(new_n981), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n754), .B1(new_n208), .B2(new_n226), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n743), .A2(new_n249), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n738), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(G150), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n775), .A2(new_n794), .B1(new_n1060), .B2(new_n778), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT51), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n758), .A2(new_n202), .B1(new_n786), .B2(new_n996), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n367), .B(new_n1063), .C1(G87), .C2(new_n772), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n768), .A2(new_n289), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n781), .A2(new_n262), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n254), .C2(new_n763), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1062), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n797), .A2(G317), .B1(G311), .B2(new_n774), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT52), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n758), .A2(new_n834), .B1(new_n786), .B2(new_n776), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n286), .B(new_n1071), .C1(G107), .C2(new_n772), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n781), .A2(new_n759), .B1(new_n602), .B2(new_n768), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(KEYINPUT119), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(KEYINPUT119), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n763), .A2(G294), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1068), .B1(new_n1070), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1059), .B1(new_n1078), .B2(new_n750), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n946), .B2(new_n803), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1054), .A2(new_n1056), .A3(new_n1080), .ZN(G390));
  INV_X1    g0881(.A(KEYINPUT120), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n921), .A2(new_n1082), .A3(G330), .A4(new_n922), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT108), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n634), .A2(new_n546), .A3(new_n678), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n723), .A2(new_n678), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT31), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1084), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n726), .A2(new_n729), .A3(KEYINPUT108), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1091), .A2(new_n922), .A3(G330), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT120), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n908), .A2(new_n896), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT39), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n925), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n899), .A2(KEYINPUT39), .A3(new_n877), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n685), .B(new_n842), .C1(new_n708), .C2(new_n664), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n907), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n896), .B1(new_n1102), .B2(new_n904), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n925), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1095), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n732), .A2(new_n842), .A3(new_n904), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(new_n891), .C2(new_n1096), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n921), .A2(G330), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n911), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n645), .B(new_n1112), .C1(new_n914), .C2(new_n915), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n905), .B1(new_n731), .B2(new_n812), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1083), .A2(new_n1094), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n906), .A2(new_n907), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT121), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(KEYINPUT121), .A3(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n905), .B1(new_n1110), .B2(new_n812), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1122), .A2(new_n907), .A3(new_n1101), .A4(new_n1107), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1113), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1109), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1108), .A3(new_n1106), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n702), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1106), .A2(new_n1108), .A3(new_n737), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n738), .B1(new_n819), .B2(new_n254), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n763), .A2(new_n1132), .B1(G159), .B2(new_n798), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n822), .B2(new_n781), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n792), .A2(G150), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  INV_X1    g0936(.A(G128), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n775), .A2(new_n830), .B1(new_n1137), .B2(new_n778), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G125), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n286), .B1(new_n262), .B2(new_n771), .C1(new_n787), .C2(new_n1140), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT123), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n208), .A2(new_n764), .B1(new_n775), .B2(new_n602), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G283), .B2(new_n797), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n367), .B1(new_n771), .B2(new_n202), .C1(new_n418), .C2(new_n758), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1065), .B(new_n1150), .C1(G107), .C2(new_n782), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(new_n766), .C2(new_n787), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1146), .A2(new_n1147), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1130), .B1(new_n1153), .B2(new_n750), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n891), .B2(new_n752), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1128), .A2(new_n1129), .A3(new_n1155), .ZN(G378));
  INV_X1    g0956(.A(new_n676), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n273), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n309), .B(new_n1158), .Z(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n752), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n775), .A2(new_n209), .B1(new_n208), .B2(new_n781), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n764), .A2(new_n350), .ZN(new_n1165));
  INV_X1    g0965(.A(G41), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1032), .A2(new_n1166), .A3(new_n367), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n771), .A2(new_n201), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n993), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n834), .B2(new_n787), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1164), .B(new_n1170), .C1(G116), .C2(new_n797), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n797), .A2(G125), .B1(G132), .B2(new_n782), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G128), .A2(new_n774), .B1(new_n763), .B2(G137), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n792), .A2(new_n1132), .B1(new_n798), .B2(G150), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT124), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(G124), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(G124), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1007), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n363), .A3(new_n1166), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G159), .B2(new_n772), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1177), .A2(new_n1178), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G50), .B1(new_n363), .B2(new_n1166), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n286), .B2(G41), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1172), .A2(new_n1185), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n750), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n738), .C1(G50), .C2(new_n819), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1163), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n923), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT40), .B1(new_n900), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n927), .A2(G330), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT125), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(G330), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n925), .B2(new_n926), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT125), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n923), .B1(new_n899), .B2(new_n877), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1198), .B(new_n1199), .C1(new_n1200), .C2(KEYINPUT40), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1196), .A2(new_n1201), .A3(new_n1161), .ZN(new_n1202));
  OAI211_X1 g1002(.A(KEYINPUT125), .B(new_n1162), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1202), .A2(new_n910), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n910), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1192), .B1(new_n1206), .B2(new_n737), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1113), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1127), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n897), .A2(new_n909), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1201), .A2(new_n1161), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1199), .B1(new_n924), .B2(new_n1198), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1203), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1211), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1202), .A2(new_n910), .A3(new_n1203), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1216), .A2(new_n1209), .A3(KEYINPUT57), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n702), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1207), .B1(new_n1210), .B2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n905), .A2(new_n751), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n738), .B1(new_n819), .B2(G68), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n797), .A2(G294), .B1(G283), .B2(new_n774), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n602), .B2(new_n781), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n286), .B(new_n990), .C1(G97), .C2(new_n792), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n763), .A2(G107), .B1(new_n517), .B2(new_n798), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n759), .C2(new_n787), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n367), .B(new_n1168), .C1(G159), .C2(new_n792), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G137), .A2(new_n774), .B1(new_n782), .B2(new_n1132), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n1137), .C2(new_n787), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n763), .A2(G150), .B1(G50), .B2(new_n798), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n830), .B2(new_n778), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1225), .A2(new_n1228), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1223), .B1(new_n1234), .B2(new_n750), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1221), .A2(new_n737), .B1(new_n1222), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1121), .A2(new_n1113), .A3(new_n1123), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1124), .A2(new_n966), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G381));
  OR2_X1    g1041(.A1(G393), .A2(G396), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(G390), .A2(new_n1242), .A3(G384), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1243), .A2(new_n984), .A3(new_n1015), .A4(new_n1240), .ZN(new_n1244));
  OR3_X1    g1044(.A1(new_n1244), .A2(G378), .A3(G375), .ZN(G407));
  INV_X1    g1045(.A(G378), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n667), .A2(G343), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G407), .B(G213), .C1(G375), .C2(new_n1248), .ZN(G409));
  NAND2_X1  g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1242), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n984), .A2(new_n1015), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n984), .B2(new_n1015), .ZN(new_n1254));
  OAI21_X1  g1054(.A(G390), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1251), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(G390), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1252), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1207), .C1(new_n1210), .C2(new_n1219), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n966), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1216), .A2(new_n1209), .A3(new_n1262), .A4(new_n1217), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1216), .A2(new_n737), .A3(new_n1217), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n1163), .C2(new_n1191), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1246), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1247), .B1(new_n1261), .B2(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1238), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT60), .B1(new_n1238), .B2(KEYINPUT126), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n702), .B(new_n1125), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(G384), .A3(new_n1236), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G384), .B1(new_n1270), .B2(new_n1236), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT62), .B1(new_n1267), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1247), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI211_X1 g1079(.A(KEYINPUT127), .B(new_n1247), .C1(new_n1261), .C2(new_n1266), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1275), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1274), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1247), .A2(G2897), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1274), .A2(G2897), .A3(new_n1247), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1260), .B1(new_n1283), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1274), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1260), .A2(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1267), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1295), .B1(new_n1296), .B2(new_n1284), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1288), .A2(new_n1296), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1293), .A2(new_n1294), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1292), .A2(new_n1299), .ZN(G405));
  XNOR2_X1  g1100(.A(G375), .B(G378), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1284), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1260), .ZN(G402));
endmodule


