//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n652, new_n655, new_n657, new_n658, new_n659, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(KEYINPUT3), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n468), .A2(new_n469), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n462), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n471), .A2(new_n474), .A3(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n466), .A2(G2105), .A3(new_n470), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n484), .B1(new_n485), .B2(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n467), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n488), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(new_n467), .A3(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n478), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n467), .A2(G138), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n470), .A2(new_n464), .A3(new_n465), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n494), .A2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n508), .A2(G651), .B1(G50), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT68), .B1(new_n517), .B2(new_n507), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n513), .B1(new_n514), .B2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(new_n518), .A2(G89), .A3(new_n522), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(KEYINPUT70), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(G651), .B1(new_n505), .B2(new_n506), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G63), .B1(new_n512), .B2(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT70), .B1(new_n526), .B2(new_n528), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n507), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n512), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n523), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n541), .B1(new_n542), .B2(G90), .ZN(G171));
  NAND2_X1  g118(.A1(new_n512), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n523), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g123(.A(KEYINPUT72), .B(new_n544), .C1(new_n523), .C2(new_n545), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n507), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n552), .A2(new_n553), .A3(G651), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n553), .B1(new_n552), .B2(G651), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n548), .A2(new_n549), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g135(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n512), .A2(new_n565), .A3(G53), .ZN(new_n566));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n569), .B1(new_n566), .B2(new_n568), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  OAI21_X1  g149(.A(G65), .B1(new_n505), .B2(new_n506), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n574), .B1(new_n577), .B2(G651), .ZN(new_n578));
  INV_X1    g153(.A(G651), .ZN(new_n579));
  AOI211_X1 g154(.A(KEYINPUT75), .B(new_n579), .C1(new_n575), .C2(new_n576), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n542), .A2(G91), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n573), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G91), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n578), .A2(new_n580), .B1(new_n523), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n565), .B1(new_n512), .B2(G53), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT74), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(new_n570), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT76), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G299));
  INV_X1    g168(.A(G171), .ZN(G301));
  INV_X1    g169(.A(G168), .ZN(G286));
  NAND3_X1  g170(.A1(new_n518), .A2(G87), .A3(new_n522), .ZN(new_n596));
  OAI211_X1 g171(.A(G49), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT77), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n519), .A2(new_n599), .A3(G49), .A4(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n602), .B(G651), .C1(new_n520), .C2(G74), .ZN(new_n603));
  NAND2_X1  g178(.A1(G74), .A2(G651), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n530), .A2(KEYINPUT78), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n596), .A2(new_n601), .A3(new_n606), .ZN(G288));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  INV_X1    g183(.A(new_n506), .ZN(new_n609));
  NAND2_X1  g184(.A1(KEYINPUT5), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G73), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(KEYINPUT79), .A2(G73), .A3(G543), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(G651), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n518), .A2(G86), .A3(new_n522), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n512), .A2(G48), .ZN(new_n621));
  OAI211_X1 g196(.A(KEYINPUT80), .B(G651), .C1(new_n611), .C2(new_n616), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n622), .ZN(G305));
  XOR2_X1   g198(.A(KEYINPUT81), .B(G85), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n542), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(G72), .A2(G543), .ZN(new_n626));
  INV_X1    g201(.A(G60), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n507), .B2(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n628), .A2(G651), .B1(G47), .B2(new_n512), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n625), .A2(new_n629), .ZN(G290));
  NAND2_X1  g205(.A1(G301), .A2(G868), .ZN(new_n631));
  INV_X1    g206(.A(G79), .ZN(new_n632));
  OR3_X1    g207(.A1(new_n632), .A2(new_n509), .A3(KEYINPUT83), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT83), .B1(new_n632), .B2(new_n509), .ZN(new_n634));
  INV_X1    g209(.A(G66), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n507), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G651), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n512), .A2(G54), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G92), .ZN(new_n641));
  OAI21_X1  g216(.A(KEYINPUT82), .B1(new_n523), .B2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n518), .A2(new_n643), .A3(G92), .A4(new_n522), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT10), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(new_n647), .A3(new_n644), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n640), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n631), .B1(new_n649), .B2(G868), .ZN(G284));
  OAI21_X1  g225(.A(new_n631), .B1(new_n649), .B2(G868), .ZN(G321));
  NAND2_X1  g226(.A1(G286), .A2(G868), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(G868), .B2(new_n592), .ZN(G297));
  OAI21_X1  g228(.A(new_n652), .B1(G868), .B2(new_n592), .ZN(G280));
  INV_X1    g229(.A(G559), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n649), .B1(new_n655), .B2(G860), .ZN(G148));
  NOR2_X1   g231(.A1(new_n557), .A2(G868), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n649), .A2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT84), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n657), .B1(new_n659), .B2(G868), .ZN(G323));
  XNOR2_X1  g235(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g236(.A1(new_n472), .A2(new_n478), .A3(G2105), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT12), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT13), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  INV_X1    g240(.A(new_n485), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G135), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT85), .ZN(new_n668));
  AND4_X1   g243(.A1(G2105), .A2(new_n470), .A3(new_n464), .A4(new_n465), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G123), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n467), .A2(G111), .ZN(new_n671));
  OAI21_X1  g246(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n668), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n673), .A2(G2096), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(G2096), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n665), .A2(new_n674), .A3(new_n675), .ZN(G156));
  XNOR2_X1  g251(.A(KEYINPUT15), .B(G2435), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT86), .B(G2438), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2427), .B(G2430), .Z(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(KEYINPUT14), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2451), .B(G2454), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT16), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1341), .B(G1348), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n683), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2443), .B(G2446), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n691), .A3(G14), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g268(.A(G2072), .B(G2078), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT17), .ZN(new_n695));
  XNOR2_X1  g270(.A(G2067), .B(G2678), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G2084), .B(G2090), .Z(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n697), .B2(new_n694), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n698), .B1(KEYINPUT88), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(KEYINPUT88), .B2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(new_n694), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n703), .A2(new_n699), .A3(new_n696), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT18), .Z(new_n705));
  NAND3_X1  g280(.A1(new_n695), .A2(new_n699), .A3(new_n697), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G2096), .B(G2100), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(G227));
  XOR2_X1   g284(.A(G1971), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT19), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1956), .B(G2474), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1961), .B(G1966), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT20), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n712), .A2(new_n713), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n711), .A2(new_n714), .A3(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(G1991), .B(G1996), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(G1981), .B(G1986), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT89), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n722), .B(new_n726), .ZN(G229));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n728), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1971), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G23), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT92), .Z(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G288), .B2(new_n728), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT33), .B(G1976), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n728), .A2(G6), .ZN(new_n738));
  INV_X1    g313(.A(G305), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n728), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT32), .B(G1981), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n732), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(G290), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G16), .B2(G24), .ZN(new_n749));
  INV_X1    g324(.A(G1986), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT94), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G25), .ZN(new_n753));
  OR2_X1    g328(.A1(G95), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT90), .Z(new_n756));
  INV_X1    g331(.A(G119), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n488), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G131), .B2(new_n666), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(new_n752), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT35), .B(G1991), .Z(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n760), .B(new_n762), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n751), .B(new_n763), .C1(new_n750), .C2(new_n749), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n745), .A2(new_n746), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(KEYINPUT95), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n745), .A2(new_n767), .A3(new_n746), .A4(new_n764), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n766), .A2(KEYINPUT36), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n752), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  OR2_X1    g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n776));
  INV_X1    g351(.A(G128), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n488), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G140), .B2(new_n666), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(new_n752), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT96), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2067), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n728), .A2(G4), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n649), .B2(new_n728), .ZN(new_n784));
  INV_X1    g359(.A(G1348), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n728), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n558), .B2(new_n728), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1341), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n782), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT97), .ZN(new_n791));
  NOR2_X1   g366(.A1(G29), .A2(G33), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT98), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT25), .Z(new_n795));
  AND2_X1   g370(.A1(new_n462), .A2(new_n477), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n796), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n797));
  INV_X1    g372(.A(G139), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n795), .B1(new_n797), .B2(new_n467), .C1(new_n485), .C2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n793), .B1(new_n799), .B2(new_n752), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2072), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n752), .A2(G32), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n669), .A2(G129), .ZN(new_n803));
  NAND3_X1  g378(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT26), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n473), .A2(G105), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G141), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n803), .B(new_n808), .C1(new_n809), .C2(new_n485), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n802), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT27), .B(G1996), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G2084), .ZN(new_n814));
  INV_X1    g389(.A(G34), .ZN(new_n815));
  AOI21_X1  g390(.A(G29), .B1(new_n815), .B2(KEYINPUT24), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(KEYINPUT24), .B2(new_n815), .ZN(new_n817));
  INV_X1    g392(.A(G160), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n752), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n801), .B(new_n813), .C1(new_n814), .C2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT99), .Z(new_n821));
  NOR2_X1   g396(.A1(G168), .A2(new_n728), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n728), .B2(G21), .ZN(new_n823));
  INV_X1    g398(.A(G1966), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT100), .ZN(new_n826));
  NAND2_X1  g401(.A1(G171), .A2(G16), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G5), .B2(G16), .ZN(new_n828));
  INV_X1    g403(.A(G1961), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n673), .A2(new_n752), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n814), .B2(new_n819), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT30), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(G28), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n752), .B1(new_n832), .B2(G28), .ZN(new_n834));
  AND2_X1   g409(.A1(KEYINPUT31), .A2(G11), .ZN(new_n835));
  NOR2_X1   g410(.A1(KEYINPUT31), .A2(G11), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n833), .A2(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n811), .A2(new_n812), .ZN(new_n838));
  AOI211_X1 g413(.A(new_n837), .B(new_n838), .C1(new_n829), .C2(new_n828), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n752), .A2(G27), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G164), .B2(new_n752), .ZN(new_n841));
  INV_X1    g416(.A(G2078), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n831), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n752), .A2(G35), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G162), .B2(new_n752), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT29), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n847), .A2(G2090), .B1(new_n824), .B2(new_n823), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(G2090), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT101), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n728), .A2(G20), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT23), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n592), .B2(new_n728), .ZN(new_n854));
  INV_X1    g429(.A(G1956), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n849), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  NOR4_X1   g432(.A1(new_n791), .A2(new_n821), .A3(new_n826), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n771), .A2(new_n772), .A3(new_n858), .ZN(G150));
  INV_X1    g434(.A(G150), .ZN(G311));
  NAND2_X1  g435(.A1(G80), .A2(G543), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n507), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n863), .A2(G651), .B1(G55), .B2(new_n512), .ZN(new_n864));
  INV_X1    g439(.A(G93), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n523), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n864), .B(new_n868), .C1(new_n865), .C2(new_n523), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n557), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n556), .A2(new_n549), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n872), .A2(new_n548), .B1(new_n869), .B2(new_n867), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n649), .A2(G559), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n877), .A2(KEYINPUT39), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(KEYINPUT39), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n878), .A2(new_n879), .A3(G860), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n866), .A2(G860), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT37), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n880), .A2(new_n882), .ZN(G145));
  XNOR2_X1  g458(.A(new_n759), .B(new_n663), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n810), .B(new_n799), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n492), .A2(new_n493), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(new_n669), .B2(G126), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n890));
  INV_X1    g465(.A(new_n497), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g467(.A(KEYINPUT103), .B(new_n497), .C1(new_n499), .C2(KEYINPUT4), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n779), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n669), .A2(G130), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n467), .A2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(G142), .B2(new_n666), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n895), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n886), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n489), .B(new_n818), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n673), .B(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n902), .A2(new_n904), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n905), .A2(new_n906), .A3(G37), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g483(.A(new_n659), .B(new_n874), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n646), .A2(new_n648), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n910), .A2(new_n591), .A3(new_n584), .A4(new_n639), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n642), .A2(new_n647), .A3(new_n644), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n647), .B1(new_n642), .B2(new_n644), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n639), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n592), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n915), .A3(KEYINPUT104), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  NAND3_X1  g492(.A1(G299), .A2(new_n917), .A3(new_n649), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n911), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n909), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n916), .A2(new_n918), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n909), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n739), .B(G290), .ZN(new_n928));
  INV_X1    g503(.A(G288), .ZN(new_n929));
  XNOR2_X1  g504(.A(G303), .B(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n928), .B(new_n930), .Z(new_n931));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n923), .A2(new_n932), .A3(new_n925), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n927), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n927), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G868), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n866), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(G295));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n938), .ZN(G331));
  NAND4_X1  g515(.A1(new_n872), .A2(new_n548), .A3(new_n867), .A4(new_n869), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n557), .A2(new_n870), .ZN(new_n942));
  OAI21_X1  g517(.A(G301), .B1(new_n533), .B2(new_n534), .ZN(new_n943));
  INV_X1    g518(.A(new_n534), .ZN(new_n944));
  NAND4_X1  g519(.A1(G171), .A2(new_n944), .A3(new_n529), .A4(new_n532), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n941), .A2(new_n942), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n871), .B2(new_n873), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n916), .A2(new_n918), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n911), .A2(new_n915), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT41), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT41), .B1(new_n916), .B2(new_n918), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT105), .B(new_n949), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n924), .A2(new_n920), .ZN(new_n956));
  AOI22_X1  g531(.A1(KEYINPUT41), .A2(new_n950), .B1(new_n948), .B2(new_n946), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n955), .A2(new_n931), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n919), .A2(new_n921), .A3(new_n952), .ZN(new_n963));
  INV_X1    g538(.A(new_n931), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n949), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n960), .A2(new_n961), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n949), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n931), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n962), .A3(new_n965), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n966), .A2(KEYINPUT106), .B1(new_n969), .B2(KEYINPUT43), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n965), .A2(new_n962), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n961), .A4(new_n960), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT44), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(new_n961), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(KEYINPUT43), .A3(new_n960), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT107), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(KEYINPUT106), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n973), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n975), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n984));
  INV_X1    g559(.A(new_n978), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n979), .A2(new_n986), .ZN(G397));
  XNOR2_X1  g562(.A(KEYINPUT108), .B(G1384), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n894), .A2(KEYINPUT109), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT109), .B1(new_n894), .B2(new_n988), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT45), .ZN(new_n991));
  AND4_X1   g566(.A1(G40), .A2(new_n471), .A3(new_n474), .A4(new_n481), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n993), .A2(G1986), .A3(G290), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n993), .A2(new_n750), .A3(new_n747), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT110), .ZN(new_n997));
  INV_X1    g572(.A(G2067), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n779), .B(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n810), .B(G1996), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n759), .B(new_n762), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n997), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT120), .B(KEYINPUT51), .Z(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n500), .B(new_n889), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1007), .B2(new_n888), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT116), .B(new_n992), .C1(new_n1008), .C2(KEYINPUT45), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n894), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n992), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1011), .B1(new_n494), .B2(new_n500), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1009), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n824), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1013), .B1(KEYINPUT50), .B2(new_n1015), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n894), .A2(new_n1021), .A3(new_n1011), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(G2084), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1006), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G168), .A2(new_n1006), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT121), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1005), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(KEYINPUT51), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1024), .B1(new_n1018), .B2(new_n824), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1006), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT122), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT122), .B(new_n1030), .C1(new_n1031), .C2(new_n1006), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1029), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT62), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1031), .A2(new_n1006), .A3(G168), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n894), .A2(new_n1011), .A3(new_n992), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n596), .A2(G1976), .A3(new_n606), .A4(new_n601), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1044), .A3(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1041), .A2(new_n1044), .A3(KEYINPUT113), .A4(G8), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(KEYINPUT52), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G305), .A2(G1981), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n620), .A2(new_n621), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n620), .A2(new_n1053), .A3(new_n621), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n617), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1050), .B1(new_n1055), .B2(G1981), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT49), .B1(new_n1056), .B2(KEYINPUT115), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n894), .A2(new_n1011), .A3(new_n992), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n1006), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  INV_X1    g637(.A(new_n617), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1051), .B2(KEYINPUT114), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1064), .B2(new_n1054), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1060), .B(new_n1061), .C1(new_n1065), .C2(new_n1050), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1057), .A2(new_n1059), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n929), .B2(G1976), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1045), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1049), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G303), .A2(G8), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1072), .B(KEYINPUT55), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n894), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n992), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1971), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT111), .B(G2090), .Z(new_n1079));
  NAND3_X1  g654(.A1(new_n1020), .A2(new_n1022), .A3(new_n1079), .ZN(new_n1080));
  AOI211_X1 g655(.A(new_n1006), .B(new_n1073), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1071), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1074), .A2(new_n842), .A3(new_n992), .A4(new_n1075), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1023), .A2(new_n829), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n842), .A2(KEYINPUT53), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1085), .B(new_n1086), .C1(new_n1018), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1021), .B1(new_n894), .B2(new_n1011), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n992), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1091), .A2(new_n1079), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1073), .B1(new_n1092), .B2(new_n1006), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1082), .A2(G171), .A3(new_n1088), .A4(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1039), .A2(new_n1040), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1081), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G288), .A2(G1976), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1050), .B1(new_n1067), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1059), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1096), .A2(new_n1071), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1101), .B1(new_n1103), .B2(new_n1073), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1082), .A2(G168), .A3(new_n1104), .A4(new_n1026), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1082), .A2(G168), .A3(new_n1026), .A4(new_n1093), .ZN(new_n1106));
  AOI22_X1  g681(.A1(KEYINPUT117), .A2(new_n1105), .B1(new_n1106), .B2(new_n1101), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1100), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT124), .B(G2078), .Z(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(new_n1084), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1074), .A2(new_n992), .A3(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1086), .B(new_n1085), .C1(new_n991), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G171), .ZN(new_n1115));
  AOI21_X1  g690(.A(G171), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1086), .B(new_n1116), .C1(new_n1018), .C2(new_n1087), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1117), .A3(KEYINPUT54), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n1093), .A3(new_n1082), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1023), .A2(new_n785), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1058), .A2(new_n998), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1023), .A2(new_n785), .B1(new_n1058), .B2(new_n998), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n914), .B1(new_n1125), .B2(KEYINPUT60), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT58), .B(G1341), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1076), .A2(G1996), .B1(new_n1058), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1128), .A2(new_n558), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1124), .A2(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1128), .A2(new_n558), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1132), .A2(new_n914), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n581), .B(new_n583), .C1(new_n587), .C2(new_n588), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT118), .B1(new_n1139), .B2(KEYINPUT57), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n573), .A2(new_n581), .A3(KEYINPUT57), .A4(new_n583), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n855), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT56), .B(G2072), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1074), .A2(new_n992), .A3(new_n1075), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1145), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1137), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1153), .A2(new_n1140), .A3(new_n1141), .A4(new_n1144), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1131), .A2(new_n1136), .A3(new_n1152), .A4(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1125), .A2(new_n914), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1149), .B1(new_n1157), .B2(new_n1151), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1119), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1088), .A2(G171), .ZN(new_n1161));
  INV_X1    g736(.A(new_n991), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1113), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1162), .A2(new_n1163), .B1(new_n829), .B2(new_n1023), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1116), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1160), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1088), .A2(G171), .B1(new_n1164), .B2(new_n1116), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT125), .B1(new_n1169), .B2(new_n1160), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1110), .A2(new_n1159), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1109), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1004), .B1(new_n1095), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n759), .A2(new_n761), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT126), .Z(new_n1176));
  AOI22_X1  g751(.A1(new_n1176), .A2(new_n1001), .B1(new_n998), .B2(new_n779), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n993), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n994), .A2(KEYINPUT48), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1179), .A2(new_n1003), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n994), .A2(KEYINPUT48), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n993), .A2(G1996), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT46), .Z(new_n1184));
  INV_X1    g759(.A(KEYINPUT47), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n991), .B(new_n992), .C1(new_n810), .C2(new_n999), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1185), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1182), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1174), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g767(.A1(G227), .A2(new_n459), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1194), .A2(new_n692), .ZN(new_n1195));
  NOR3_X1   g769(.A1(new_n907), .A2(G229), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1196), .A2(new_n982), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


