//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT77), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT11), .B1(new_n198), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G134), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n201), .B2(G134), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(KEYINPUT66), .A3(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n199), .A2(new_n202), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n205), .A4(new_n206), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT64), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n215), .B1(new_n220), .B2(new_n214), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(G143), .A3(new_n219), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n217), .B2(G143), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT64), .A2(G146), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT64), .A2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n230), .B1(new_n233), .B2(G143), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n218), .A2(KEYINPUT65), .A3(G143), .A4(new_n219), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n228), .B(G128), .C1(new_n234), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n227), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT78), .B(G101), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT3), .B1(new_n240), .B2(G107), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n242));
  INV_X1    g056(.A(G107), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(G104), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(G107), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n239), .A2(new_n241), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n245), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n240), .A2(G107), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT10), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT0), .B(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n221), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  INV_X1    g069(.A(new_n230), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n223), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n255), .B1(new_n257), .B2(new_n235), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n254), .B1(new_n258), .B2(KEYINPUT0), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n241), .A2(new_n244), .A3(new_n245), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT78), .B(G101), .Z(new_n261));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(G101), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(KEYINPUT4), .A3(G101), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n238), .A2(new_n252), .B1(new_n259), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n250), .ZN(new_n268));
  AOI211_X1 g082(.A(KEYINPUT1), .B(new_n255), .C1(new_n257), .C2(new_n235), .ZN(new_n269));
  OAI21_X1  g083(.A(G128), .B1(new_n215), .B2(new_n228), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n257), .A2(new_n235), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n268), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT79), .B1(new_n273), .B2(new_n251), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n250), .B1(new_n237), .B2(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT79), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT10), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n213), .B(new_n267), .C1(new_n274), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n227), .A2(new_n250), .A3(new_n237), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n273), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n212), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT12), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT12), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n283), .A3(new_n212), .ZN(new_n284));
  AND4_X1   g098(.A1(KEYINPUT80), .A2(new_n278), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n280), .B2(new_n212), .ZN(new_n286));
  AOI211_X1 g100(.A(KEYINPUT12), .B(new_n213), .C1(new_n279), .C2(new_n273), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT80), .B1(new_n288), .B2(new_n278), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n197), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n267), .B1(new_n274), .B2(new_n277), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n212), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n197), .B1(new_n292), .B2(new_n278), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n190), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G469), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n278), .A2(new_n282), .A3(new_n196), .A4(new_n284), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT82), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT82), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n288), .A2(new_n299), .A3(new_n196), .A4(new_n278), .ZN(new_n300));
  INV_X1    g114(.A(new_n278), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n273), .A2(KEYINPUT79), .A3(new_n251), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n276), .B1(new_n275), .B2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n213), .B1(new_n304), .B2(new_n267), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n197), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n298), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT81), .B(G469), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n190), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n191), .B1(new_n296), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n198), .A2(G137), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n201), .A2(G134), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n211), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n227), .B2(new_n237), .ZN(new_n315));
  OAI211_X1 g129(.A(KEYINPUT0), .B(G128), .C1(new_n234), .C2(new_n236), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n221), .A2(new_n253), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n212), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT2), .B(G113), .Z(new_n319));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n320));
  INV_X1    g134(.A(G116), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(G119), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT68), .A3(G116), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(G119), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n319), .A2(new_n322), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT2), .B(G113), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n315), .A2(new_n318), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT30), .B1(new_n315), .B2(new_n318), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n212), .A2(new_n316), .A3(new_n317), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT67), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(G128), .A3(new_n224), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n338), .A2(new_n222), .B1(new_n228), .B2(new_n258), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n333), .B(new_n334), .C1(new_n339), .C2(new_n314), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n331), .B1(new_n341), .B2(new_n330), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G237), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n192), .A3(G210), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n345), .B(KEYINPUT27), .Z(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G101), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n350));
  INV_X1    g164(.A(new_n348), .ZN(new_n351));
  INV_X1    g165(.A(new_n314), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n238), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n330), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n334), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT69), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n330), .B1(new_n315), .B2(new_n318), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT28), .B1(new_n359), .B2(new_n358), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n351), .B(new_n357), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n349), .A2(new_n350), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n354), .B1(new_n353), .B2(new_n334), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n364), .B1(new_n331), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n355), .A2(KEYINPUT70), .A3(new_n359), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(KEYINPUT28), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n357), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n351), .A2(KEYINPUT29), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n190), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G472), .B1(new_n363), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT31), .B1(new_n342), .B2(new_n351), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n354), .B1(new_n332), .B2(new_n340), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT31), .ZN(new_n375));
  NOR4_X1   g189(.A1(new_n374), .A2(new_n375), .A3(new_n348), .A4(new_n331), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n356), .B1(new_n364), .B2(KEYINPUT69), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n377), .A2(new_n378), .B1(new_n356), .B2(new_n355), .ZN(new_n379));
  OAI22_X1  g193(.A1(new_n373), .A2(new_n376), .B1(new_n379), .B2(new_n351), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT32), .ZN(new_n381));
  NOR2_X1   g195(.A1(G472), .A2(G902), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n372), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G214), .B1(G237), .B2(G902), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT5), .A4(new_n325), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n321), .A2(KEYINPUT5), .A3(G119), .ZN(new_n388));
  INV_X1    g202(.A(G113), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT84), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  AND4_X1   g208(.A1(new_n268), .A2(new_n392), .A3(new_n326), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n266), .B2(new_n330), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n246), .A2(KEYINPUT4), .B1(G101), .B2(new_n260), .ZN(new_n399));
  INV_X1    g213(.A(new_n265), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n397), .B(new_n330), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n396), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G122), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n330), .B1(new_n399), .B2(new_n400), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT83), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n395), .B1(new_n408), .B2(new_n401), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n404), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G125), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n316), .B2(new_n317), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n339), .B2(new_n412), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n192), .A2(G224), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n415), .B(KEYINPUT86), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n414), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n401), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n404), .B1(new_n419), .B2(new_n396), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT85), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n423));
  NOR4_X1   g237(.A1(new_n409), .A2(new_n423), .A3(KEYINPUT6), .A4(new_n404), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n411), .B(new_n418), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n415), .A2(KEYINPUT7), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n392), .A2(new_n326), .A3(new_n394), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n326), .A2(new_n246), .A3(new_n249), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n427), .A2(new_n250), .B1(new_n428), .B2(new_n391), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n404), .B(KEYINPUT8), .Z(new_n430));
  OAI22_X1  g244(.A1(new_n414), .A2(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI211_X1 g245(.A(new_n405), .B(new_n395), .C1(new_n408), .C2(new_n401), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n413), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n434), .B(new_n426), .C1(new_n238), .C2(G125), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT87), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n414), .A2(new_n437), .A3(new_n426), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G210), .B1(G237), .B2(G902), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n425), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n425), .B2(new_n440), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n386), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G478), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(KEYINPUT15), .ZN(new_n446));
  INV_X1    g260(.A(G122), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G116), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n321), .A2(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(KEYINPUT94), .ZN(new_n451));
  XNOR2_X1  g265(.A(G116), .B(G122), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT94), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n243), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n450), .A2(KEYINPUT94), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n453), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(G107), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n214), .A2(G128), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT13), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n214), .A2(G128), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT95), .B1(new_n462), .B2(new_n461), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n462), .A2(KEYINPUT95), .A3(new_n461), .ZN(new_n466));
  OAI21_X1  g280(.A(G134), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n462), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(new_n460), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n198), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n459), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G134), .B1(new_n468), .B2(new_n460), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n449), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(new_n243), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n452), .A2(new_n473), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n470), .A2(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n455), .ZN(new_n478));
  INV_X1    g292(.A(G217), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n188), .A2(new_n479), .A3(G953), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n471), .A2(KEYINPUT96), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n455), .A2(new_n458), .B1(new_n198), .B2(new_n469), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n482), .A2(new_n467), .B1(new_n455), .B2(new_n477), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n483), .B2(new_n480), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT96), .B1(new_n483), .B2(new_n480), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n190), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT97), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n446), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n487), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n471), .A2(new_n478), .ZN(new_n491));
  INV_X1    g305(.A(new_n480), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n492), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n481), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT97), .A3(new_n190), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n488), .B1(new_n497), .B2(new_n446), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n344), .A2(new_n192), .A3(G214), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT90), .B1(new_n500), .B2(G143), .ZN(new_n501));
  OR2_X1    g315(.A1(KEYINPUT90), .A2(G143), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n501), .A2(new_n499), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT18), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(new_n210), .ZN(new_n507));
  INV_X1    g321(.A(G140), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G125), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n412), .A2(G140), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT72), .ZN(new_n512));
  XNOR2_X1  g326(.A(G125), .B(G140), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n515), .A3(new_n233), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n217), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g331(.A(G131), .B1(new_n503), .B2(new_n504), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n507), .B(new_n517), .C1(new_n506), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(KEYINPUT91), .B(G131), .C1(new_n503), .C2(new_n504), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(KEYINPUT17), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n513), .A2(KEYINPUT16), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n509), .A2(KEYINPUT16), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n217), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(G146), .A3(new_n525), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n530), .A3(KEYINPUT92), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n505), .A2(new_n210), .ZN(new_n533));
  INV_X1    g347(.A(new_n521), .ZN(new_n534));
  INV_X1    g348(.A(new_n522), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT92), .B1(new_n523), .B2(new_n530), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n519), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G113), .B(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G104), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n519), .A2(new_n541), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n545));
  INV_X1    g359(.A(new_n528), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n512), .A2(new_n515), .ZN(new_n547));
  MUX2_X1   g361(.A(new_n547), .B(new_n513), .S(KEYINPUT19), .Z(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n548), .B2(new_n233), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n544), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT20), .ZN(new_n552));
  NOR2_X1   g366(.A1(G475), .A2(G902), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n543), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n553), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n555), .B(new_n550), .C1(new_n539), .C2(new_n542), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n542), .A2(KEYINPUT93), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n539), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n190), .B1(new_n539), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g375(.A(G475), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT98), .B(G952), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G953), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n498), .A2(new_n558), .A3(new_n562), .A4(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n444), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n479), .B1(G234), .B2(new_n190), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT73), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT74), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n578), .A2(KEYINPUT73), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(KEYINPUT73), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G234), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n187), .A2(new_n585), .A3(G953), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n580), .B2(new_n584), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n577), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n580), .A2(new_n584), .ZN(new_n591));
  INV_X1    g405(.A(new_n586), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(KEYINPUT75), .A3(new_n587), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n255), .A2(KEYINPUT23), .A3(G119), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n323), .A2(G128), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n323), .A2(G128), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(KEYINPUT23), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT71), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G110), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n599), .A2(KEYINPUT71), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n255), .A2(G119), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT24), .B(G110), .ZN(new_n605));
  OAI221_X1 g419(.A(new_n529), .B1(new_n601), .B2(new_n602), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n599), .B2(G110), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n516), .A3(new_n528), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n595), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n606), .B(new_n609), .C1(new_n588), .C2(new_n589), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT25), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n613), .B2(KEYINPUT76), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(KEYINPUT76), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n576), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n616), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n611), .A2(new_n618), .A3(new_n612), .A4(new_n614), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n575), .A2(G902), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n611), .A2(new_n612), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n310), .A2(new_n385), .A3(new_n574), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(new_n261), .ZN(G3));
  OAI211_X1 g440(.A(new_n386), .B(new_n572), .C1(new_n442), .C2(new_n443), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n558), .A2(new_n562), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n492), .A2(KEYINPUT99), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n491), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n491), .A2(new_n630), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n495), .A2(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n445), .A2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n486), .A2(new_n445), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n628), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n380), .B2(new_n190), .ZN(new_n642));
  INV_X1    g456(.A(new_n382), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n341), .A2(new_n330), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n351), .A3(new_n355), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n375), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n342), .A2(KEYINPUT31), .A3(new_n351), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n348), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n643), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n642), .A2(new_n651), .A3(new_n623), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n310), .A2(new_n640), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  NOR2_X1   g469(.A1(new_n486), .A2(new_n487), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT97), .B1(new_n495), .B2(new_n190), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n446), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n488), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n556), .A2(new_n557), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n556), .A2(new_n557), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n660), .B(new_n562), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n627), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n310), .A3(new_n652), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  INV_X1    g481(.A(KEYINPUT36), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n590), .A2(new_n594), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n610), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n617), .A2(new_n619), .B1(new_n621), .B2(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n642), .A2(new_n651), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n310), .A2(new_n574), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  AOI22_X1  g490(.A1(new_n646), .A2(new_n647), .B1(new_n348), .B2(new_n649), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT32), .B1(new_n677), .B2(new_n643), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n672), .B1(new_n680), .B2(new_n372), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n567), .B1(new_n682), .B2(new_n570), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n562), .B(new_n684), .C1(new_n662), .C2(new_n661), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n498), .ZN(new_n686));
  INV_X1    g500(.A(new_n386), .ZN(new_n687));
  INV_X1    g501(.A(new_n443), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n425), .A2(new_n440), .A3(new_n441), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n681), .A2(new_n310), .A3(new_n686), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  XOR2_X1   g506(.A(new_n683), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n310), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT100), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n688), .A2(new_n689), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT38), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n343), .A2(new_n351), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n366), .A2(new_n367), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n700), .B(new_n190), .C1(new_n351), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G472), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n680), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n628), .A2(new_n660), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n672), .A2(new_n386), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n699), .A2(new_n705), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n696), .A2(new_n697), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  AOI22_X1  g524(.A1(new_n634), .A2(new_n635), .B1(new_n445), .B2(new_n486), .ZN(new_n711));
  AOI211_X1 g525(.A(new_n683), .B(new_n711), .C1(new_n558), .C2(new_n562), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n681), .A2(new_n310), .A3(new_n690), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  AND3_X1   g528(.A1(new_n307), .A2(new_n190), .A3(new_n308), .ZN(new_n715));
  INV_X1    g529(.A(G469), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n307), .B2(new_n190), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n715), .A2(new_n717), .A3(new_n191), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n640), .A2(new_n385), .A3(new_n624), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n664), .A2(new_n385), .A3(new_n624), .A4(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  INV_X1    g537(.A(new_n191), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n292), .A2(new_n278), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n197), .A2(new_n725), .B1(new_n297), .B2(KEYINPUT82), .ZN(new_n726));
  AOI21_X1  g540(.A(G902), .B1(new_n726), .B2(new_n300), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n724), .B(new_n309), .C1(new_n727), .C2(new_n716), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n444), .ZN(new_n729));
  INV_X1    g543(.A(new_n573), .ZN(new_n730));
  INV_X1    g544(.A(new_n672), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n729), .A2(new_n730), .A3(new_n385), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  NOR2_X1   g547(.A1(new_n706), .A2(new_n444), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n369), .A2(new_n348), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n643), .B1(new_n648), .B2(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n642), .A2(new_n736), .A3(new_n623), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n734), .A2(new_n737), .A3(new_n718), .A4(new_n572), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT101), .B(G122), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G24));
  NOR3_X1   g554(.A1(new_n642), .A2(new_n736), .A3(new_n672), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n729), .A2(new_n712), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NOR3_X1   g557(.A1(new_n442), .A2(new_n443), .A3(new_n687), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n310), .A2(new_n385), .A3(new_n624), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(KEYINPUT42), .A3(new_n712), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n310), .A2(new_n385), .A3(new_n624), .A4(new_n744), .ZN(new_n748));
  INV_X1    g562(.A(new_n712), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  INV_X1    g566(.A(new_n686), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n198), .ZN(G36));
  NOR2_X1   g569(.A1(new_n716), .A2(new_n190), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n290), .A2(new_n294), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n716), .B1(new_n757), .B2(KEYINPUT45), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(KEYINPUT45), .B2(new_n757), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT102), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n756), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n309), .B1(new_n763), .B2(KEYINPUT46), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n688), .A2(new_n386), .A3(new_n689), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT105), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n628), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n638), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT103), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT43), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n638), .A2(KEYINPUT104), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n638), .B1(KEYINPUT104), .B2(KEYINPUT43), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n770), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n772), .A2(KEYINPUT43), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n773), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n731), .B1(new_n642), .B2(new_n651), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT44), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n769), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n766), .A2(new_n724), .A3(new_n693), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  OAI21_X1  g598(.A(new_n724), .B1(new_n764), .B2(new_n765), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(KEYINPUT47), .B(new_n724), .C1(new_n764), .C2(new_n765), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n749), .A2(new_n385), .A3(new_n624), .A4(new_n767), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT106), .Z(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n704), .A2(new_n566), .A3(new_n623), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n718), .A3(new_n744), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n628), .A3(new_n638), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n773), .A2(new_n567), .A3(new_n776), .A4(new_n777), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n728), .A3(new_n767), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT116), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n797), .B1(new_n800), .B2(new_n741), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n802));
  INV_X1    g616(.A(new_n737), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n699), .A2(new_n687), .A3(new_n718), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n807));
  INV_X1    g621(.A(new_n699), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n386), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n798), .A2(new_n803), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n810), .A3(KEYINPUT112), .A4(new_n718), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n806), .A2(new_n811), .A3(new_n814), .A4(new_n807), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n809), .A2(new_n810), .A3(new_n718), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n817), .A2(KEYINPUT114), .A3(new_n807), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT114), .B1(new_n817), .B2(new_n807), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n816), .A2(KEYINPUT115), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT115), .B1(new_n816), .B2(new_n820), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n801), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n804), .A2(new_n769), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n715), .A2(new_n717), .A3(new_n724), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n789), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n787), .A2(KEYINPUT111), .A3(new_n788), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n794), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  AOI211_X1 g645(.A(G953), .B(new_n563), .C1(new_n810), .C2(new_n729), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n623), .B1(new_n680), .B2(new_n372), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n800), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n834), .A2(KEYINPUT48), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(KEYINPUT48), .ZN(new_n836));
  OAI221_X1 g650(.A(new_n832), .B1(new_n639), .B2(new_n796), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n801), .A2(KEYINPUT51), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n816), .B2(new_n820), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n824), .B1(new_n789), .B2(new_n826), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n831), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n731), .A2(new_n683), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n704), .A2(new_n310), .A3(new_n734), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n691), .A2(new_n713), .A3(new_n742), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT108), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n685), .A2(new_n660), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n385), .A2(new_n849), .A3(new_n731), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n278), .A2(new_n282), .A3(new_n284), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT80), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n288), .A2(KEYINPUT80), .A3(new_n278), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n293), .B1(new_n855), .B2(new_n197), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n716), .B1(new_n856), .B2(new_n190), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n744), .B(new_n724), .C1(new_n857), .C2(new_n715), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n848), .B1(new_n850), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n858), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n681), .A3(KEYINPUT108), .A4(new_n849), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n741), .A2(new_n712), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n745), .A2(new_n686), .B1(new_n863), .B2(new_n860), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n660), .A2(new_n558), .A3(new_n562), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n627), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n310), .A2(new_n867), .A3(new_n652), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n674), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT107), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT107), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n674), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n625), .A2(new_n653), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT110), .B1(new_n865), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n732), .A2(new_n722), .A3(new_n719), .A4(new_n738), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n751), .A2(new_n877), .A3(KEYINPUT53), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n868), .A2(new_n674), .A3(new_n871), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n871), .B1(new_n868), .B2(new_n674), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n625), .A2(new_n653), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n310), .A2(new_n741), .A3(new_n712), .A4(new_n744), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n748), .B2(new_n753), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n859), .B2(new_n861), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT110), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n847), .A2(new_n875), .A3(new_n878), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n876), .B1(new_n750), .B2(new_n746), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n882), .A3(new_n885), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n310), .A2(new_n385), .A3(new_n690), .A4(new_n731), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n892), .A2(new_n686), .B1(new_n729), .B2(new_n863), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n846), .A3(new_n713), .A4(new_n844), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n845), .A2(KEYINPUT52), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n889), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n888), .A2(new_n897), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n865), .A2(new_n874), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n847), .A2(KEYINPUT53), .A3(new_n900), .A4(new_n890), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n897), .A3(KEYINPUT109), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT109), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n903), .B(new_n889), .C1(new_n891), .C2(new_n896), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(KEYINPUT54), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  OAI22_X1  g720(.A1(new_n842), .A2(new_n906), .B1(G952), .B2(G953), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT49), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n715), .A2(new_n717), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n808), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n724), .A2(new_n386), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n704), .A2(new_n623), .A3(new_n771), .A4(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n910), .B(new_n912), .C1(new_n908), .C2(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n907), .A2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n192), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n190), .B1(new_n888), .B2(new_n897), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n411), .B1(new_n422), .B2(new_n424), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n418), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n921), .B2(new_n918), .ZN(G51));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n899), .A2(new_n924), .ZN(new_n925));
  OR3_X1    g739(.A1(new_n898), .A2(new_n924), .A3(KEYINPUT54), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n756), .B(KEYINPUT57), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n307), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n917), .A2(new_n762), .A3(new_n761), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n915), .B1(new_n931), .B2(new_n932), .ZN(G54));
  NAND3_X1  g747(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n543), .A2(new_n551), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n916), .B1(new_n934), .B2(new_n935), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G60));
  INV_X1    g755(.A(new_n634), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n928), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n916), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n899), .B2(new_n905), .ZN(new_n948));
  OR3_X1    g762(.A1(new_n948), .A2(KEYINPUT119), .A3(new_n634), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT119), .B1(new_n948), .B2(new_n634), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT60), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT120), .B1(new_n898), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT120), .ZN(new_n956));
  AOI211_X1 g770(.A(new_n956), .B(new_n953), .C1(new_n888), .C2(new_n897), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n611), .A2(new_n612), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n915), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n898), .A2(new_n954), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n956), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n898), .A2(KEYINPUT120), .A3(new_n954), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n961), .B1(new_n965), .B2(new_n671), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n961), .B(new_n671), .C1(new_n955), .C2(new_n957), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n960), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n960), .B(new_n970), .C1(new_n966), .C2(new_n968), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(G66));
  INV_X1    g788(.A(G224), .ZN(new_n975));
  OAI21_X1  g789(.A(G953), .B1(new_n568), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n874), .A2(new_n876), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(G953), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n919), .B1(G898), .B2(new_n192), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G69));
  INV_X1    g794(.A(G227), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n341), .B(new_n548), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI221_X1 g797(.A(G953), .B1(new_n981), .B2(new_n682), .C1(new_n983), .C2(KEYINPUT125), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n766), .A2(new_n724), .A3(new_n693), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT124), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n833), .A2(new_n734), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n987), .B1(new_n986), .B2(new_n988), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n754), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n893), .A2(new_n713), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  AND4_X1   g808(.A1(new_n751), .A2(new_n783), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n991), .A2(new_n192), .A3(new_n995), .A4(new_n792), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n983), .B1(G900), .B2(G953), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n767), .B1(new_n639), .B2(new_n866), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n833), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n695), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n783), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT123), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT123), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n783), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n709), .A2(new_n994), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT62), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1007), .A2(new_n792), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n982), .B1(new_n1010), .B2(new_n192), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n985), .B1(new_n999), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1010), .A2(new_n192), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n998), .B(new_n984), .C1(new_n1013), .C2(new_n982), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1014), .ZN(G72));
  NAND4_X1  g829(.A1(new_n1007), .A2(new_n792), .A3(new_n977), .A4(new_n1009), .ZN(new_n1016));
  XNOR2_X1  g830(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n700), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n342), .A2(new_n348), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n991), .A2(new_n792), .A3(new_n995), .A4(new_n977), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1021), .B1(new_n1022), .B2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n902), .A2(new_n904), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n349), .A2(new_n645), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n1019), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n916), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n1020), .A2(new_n1023), .A3(new_n1027), .ZN(G57));
endmodule


