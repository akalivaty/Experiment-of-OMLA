//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n211), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n219), .B1(new_n214), .B2(new_n213), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT65), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  OAI21_X1  g0051(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n209), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n215), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n221), .B1(new_n208), .B2(G20), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT69), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n263), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G50), .B2(new_n270), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT9), .ZN(new_n277));
  OR3_X1    g0077(.A1(new_n265), .A2(KEYINPUT9), .A3(new_n274), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT67), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n284), .B(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n286), .A2(G223), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G222), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n289), .A2(new_n290), .B1(new_n223), .B2(new_n283), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n282), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n282), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(new_n293), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n297), .B2(G226), .ZN(new_n298));
  AOI21_X1  g0098(.A(G200), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n292), .A2(new_n298), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT10), .B1(new_n281), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n299), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G190), .B2(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT70), .B1(new_n277), .B2(new_n278), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n301), .A2(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n300), .A2(G169), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n275), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n272), .B1(G1), .B2(new_n209), .ZN(new_n315));
  MUX2_X1   g0115(.A(new_n270), .B(new_n315), .S(G77), .Z(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT15), .B(G87), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n317), .A2(new_n259), .B1(new_n209), .B2(new_n223), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n257), .A2(new_n255), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n263), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n286), .A2(G238), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n283), .A2(G232), .A3(new_n288), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n205), .B2(new_n283), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n282), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n295), .B1(new_n297), .B2(G244), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(G190), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n321), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n321), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(G169), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n325), .A2(G179), .A3(new_n326), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n310), .A2(new_n314), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G68), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n269), .A2(G20), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT12), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n315), .B2(new_n339), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n260), .A2(G77), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n339), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n264), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n346));
  XNOR2_X1  g0146(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G97), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n289), .C2(new_n222), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n282), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n295), .B1(new_n297), .B2(G238), .ZN(new_n353));
  XOR2_X1   g0153(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n353), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  OAI211_X1 g0158(.A(G190), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n354), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n330), .B1(new_n361), .B2(new_n355), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT72), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n362), .A2(KEYINPUT72), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n348), .B(new_n359), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n355), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n354), .B1(new_n352), .B2(new_n353), .ZN(new_n368));
  OAI21_X1  g0168(.A(G169), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT14), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n371), .B(G169), .C1(new_n367), .C2(new_n368), .ZN(new_n372));
  OAI211_X1 g0172(.A(G179), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n348), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n366), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G58), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n339), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n379), .B2(new_n201), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n254), .A2(G159), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT3), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(G33), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(G33), .ZN(new_n386));
  INV_X1    g0186(.A(G33), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n209), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n339), .B1(new_n390), .B2(KEYINPUT7), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n392), .A3(new_n209), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n382), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT75), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT7), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n209), .B1(new_n396), .B2(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n283), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(G20), .B1(new_n392), .B2(KEYINPUT75), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n384), .A2(G33), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n401), .B(new_n397), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(G68), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(new_n380), .A3(new_n381), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n264), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n258), .A2(new_n271), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n315), .A2(new_n258), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n395), .A2(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n296), .A2(new_n293), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n412), .A2(new_n237), .B1(new_n294), .B2(new_n293), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n288), .A2(G223), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n222), .B2(new_n288), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n415), .A2(new_n385), .A3(new_n386), .A4(new_n388), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n296), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n302), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(G200), .B2(new_n419), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n411), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n419), .A2(G169), .ZN(new_n425));
  INV_X1    g0225(.A(G179), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n419), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n395), .A2(new_n408), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n410), .A2(new_n409), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n419), .A2(new_n426), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G169), .B2(new_n419), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT18), .B1(new_n411), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n411), .A2(KEYINPUT17), .A3(new_n421), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n424), .A2(new_n432), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n338), .A2(new_n377), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G238), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1698), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n385), .A2(new_n388), .A3(new_n441), .A4(new_n386), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G116), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT83), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT74), .B1(new_n387), .B2(KEYINPUT3), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n403), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(G244), .A3(G1698), .A4(new_n388), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n385), .A2(new_n388), .A3(G244), .A4(new_n386), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n442), .B(new_n443), .C1(new_n450), .C2(new_n288), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT83), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n452), .A3(new_n282), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n208), .A2(G45), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT82), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n455), .A3(G250), .ZN(new_n456));
  AOI21_X1  g0256(.A(G274), .B1(KEYINPUT82), .B2(G250), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n296), .B(new_n456), .C1(new_n454), .C2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n302), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n385), .A2(new_n388), .A3(new_n209), .A4(new_n386), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n339), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n350), .A2(KEYINPUT19), .A3(G20), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n350), .A2(new_n209), .ZN(new_n464));
  INV_X1    g0264(.A(G87), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n204), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n466), .B2(G107), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n463), .B1(new_n467), .B2(KEYINPUT19), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n263), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n208), .A2(G33), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n264), .A2(new_n270), .A3(new_n470), .ZN(new_n471));
  OR3_X1    g0271(.A1(new_n471), .A2(KEYINPUT84), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n271), .A2(new_n317), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT84), .B1(new_n471), .B2(new_n465), .ZN(new_n474));
  AND4_X1   g0274(.A1(new_n469), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n282), .B1(new_n451), .B2(KEYINPUT83), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n445), .B1(new_n444), .B2(new_n448), .ZN(new_n477));
  OAI211_X1 g0277(.A(G200), .B(new_n458), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G169), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n458), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n469), .B(new_n473), .C1(new_n471), .C2(new_n317), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(G179), .B1(new_n453), .B2(new_n458), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n460), .A2(new_n479), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n471), .A2(G97), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G97), .B2(new_n271), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n400), .A2(G107), .A3(new_n404), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G97), .A2(G107), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n206), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT77), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT6), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n206), .A2(new_n492), .A3(new_n493), .A4(new_n490), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n204), .A2(KEYINPUT6), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n495), .A2(G20), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n254), .A2(G77), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT76), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n489), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT78), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n501), .A2(new_n502), .A3(new_n263), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n501), .B2(new_n263), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n488), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT79), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(KEYINPUT79), .B(new_n488), .C1(new_n503), .C2(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n224), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n283), .A2(new_n288), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n510), .B1(new_n450), .B2(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n282), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT80), .ZN(new_n518));
  INV_X1    g0318(.A(G41), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n520), .B2(new_n454), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G41), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(KEYINPUT80), .A3(new_n208), .A4(G45), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G257), .A3(new_n296), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n296), .A2(G274), .A3(new_n525), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n521), .A2(KEYINPUT81), .A3(new_n524), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT81), .B1(new_n521), .B2(new_n524), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n517), .A2(new_n302), .A3(new_n527), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n527), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n296), .B1(new_n514), .B2(new_n515), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n535), .B2(G200), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n507), .A2(new_n508), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n517), .A2(new_n426), .A3(new_n527), .A4(new_n531), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n505), .B(new_n538), .C1(G169), .C2(new_n535), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n486), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n526), .A2(G264), .A3(new_n296), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT87), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT87), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n526), .A2(new_n543), .A3(G264), .A4(new_n296), .ZN(new_n544));
  INV_X1    g0344(.A(G250), .ZN(new_n545));
  INV_X1    g0345(.A(G257), .ZN(new_n546));
  MUX2_X1   g0346(.A(new_n545), .B(new_n546), .S(G1698), .Z(new_n547));
  INV_X1    g0347(.A(G294), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n389), .A2(new_n547), .B1(new_n387), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n282), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n542), .A2(new_n531), .A3(new_n544), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n330), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(G190), .B2(new_n551), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT86), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n386), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n209), .A3(G87), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n465), .A2(KEYINPUT22), .A3(G20), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n283), .A2(KEYINPUT86), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT22), .B1(new_n461), .B2(new_n465), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n209), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  INV_X1    g0367(.A(new_n443), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n566), .A2(new_n567), .B1(new_n568), .B2(new_n209), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n263), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT24), .B1(new_n564), .B2(new_n569), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n269), .A2(G20), .A3(new_n205), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT25), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n471), .A2(new_n205), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n553), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n526), .A2(G270), .A3(new_n296), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n546), .A2(G1698), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(G264), .B2(G1698), .ZN(new_n582));
  INV_X1    g0382(.A(G303), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n582), .A2(new_n389), .B1(new_n583), .B2(new_n283), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n282), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n531), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(KEYINPUT21), .A3(G169), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n531), .A2(G179), .A3(new_n580), .A4(new_n585), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n471), .A2(G116), .ZN(new_n590));
  INV_X1    g0390(.A(G116), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n270), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(G20), .B1(G33), .B2(G283), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n387), .A2(G97), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT85), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n262), .A2(new_n215), .B1(G20), .B2(new_n591), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT20), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n596), .A2(new_n597), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT85), .B1(new_n594), .B2(new_n595), .ZN(new_n602));
  OAI211_X1 g0402(.A(KEYINPUT20), .B(new_n599), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n593), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(G169), .A3(new_n586), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n589), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n551), .A2(G169), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n541), .A2(KEYINPUT87), .B1(new_n282), .B2(new_n549), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(G179), .A3(new_n531), .A4(new_n544), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n578), .B1(new_n572), .B2(new_n573), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n605), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n586), .A2(new_n330), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n586), .A2(G190), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n579), .A2(new_n608), .A3(new_n614), .A4(new_n618), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n439), .A2(new_n540), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT88), .ZN(G372));
  NAND2_X1  g0421(.A1(new_n589), .A2(new_n605), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n607), .A2(new_n606), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n614), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n579), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n540), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n481), .A2(new_n482), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n484), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n538), .B1(new_n535), .B2(G169), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n507), .B2(new_n508), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT26), .B1(new_n631), .B2(new_n486), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n475), .A2(new_n478), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n633), .A2(new_n459), .B1(new_n627), .B2(new_n484), .ZN(new_n634));
  XNOR2_X1  g0434(.A(KEYINPUT89), .B(KEYINPUT26), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n539), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n629), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n438), .B1(new_n626), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT90), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT90), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n432), .A2(new_n435), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n366), .A2(new_n336), .B1(new_n375), .B2(new_n374), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n424), .A2(new_n436), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n313), .B1(new_n644), .B2(new_n310), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n639), .A2(new_n640), .A3(new_n645), .ZN(G369));
  INV_X1    g0446(.A(new_n269), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .A3(G20), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT27), .B1(new_n647), .B2(G20), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n612), .A2(new_n613), .A3(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT91), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n613), .A2(new_n652), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n579), .A2(new_n614), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(KEYINPUT91), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n608), .A2(new_n652), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n614), .A2(new_n652), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n608), .A2(new_n618), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n605), .A2(new_n652), .ZN(new_n664));
  MUX2_X1   g0464(.A(new_n608), .B(new_n663), .S(new_n664), .Z(new_n665));
  INV_X1    g0465(.A(G330), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n658), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n662), .A2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n212), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n466), .A2(G107), .A3(G116), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n217), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n652), .A2(KEYINPUT31), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n517), .A2(new_n527), .A3(new_n531), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n610), .A2(new_n544), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n678), .A2(new_n679), .A3(new_n588), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n453), .A2(new_n458), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(KEYINPUT30), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n681), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n586), .A2(new_n426), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(new_n678), .A4(new_n551), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT30), .B1(new_n680), .B2(new_n681), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n677), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT92), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n678), .A2(new_n679), .ZN(new_n691));
  INV_X1    g0491(.A(new_n588), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n681), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n682), .A3(new_n685), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(KEYINPUT92), .A3(new_n677), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n652), .B1(new_n696), .B2(KEYINPUT31), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT31), .B1(new_n540), .B2(new_n619), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n666), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n624), .A2(new_n486), .A3(new_n579), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n537), .A2(new_n539), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n537), .A2(KEYINPUT93), .A3(new_n539), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n631), .A2(new_n486), .A3(KEYINPUT26), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n635), .B1(new_n539), .B2(new_n634), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n628), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n652), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  INV_X1    g0513(.A(new_n652), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n637), .B2(new_n626), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n702), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n676), .B1(new_n718), .B2(G1), .ZN(G364));
  NOR2_X1   g0519(.A1(new_n268), .A2(G20), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G45), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n672), .A2(G1), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n665), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n209), .A2(new_n302), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n426), .A3(G200), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT95), .Z(new_n729));
  AOI21_X1  g0529(.A(new_n283), .B1(new_n729), .B2(G303), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT96), .Z(new_n731));
  NOR2_X1   g0531(.A1(new_n426), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G322), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n426), .A2(new_n330), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n727), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G326), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n209), .A2(G190), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n732), .ZN(new_n740));
  INV_X1    g0540(.A(G311), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n737), .A2(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n739), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(G179), .A3(new_n330), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n735), .B(new_n742), .C1(G283), .C2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(new_n426), .A3(new_n330), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G329), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n302), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n209), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G294), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n736), .A2(new_n739), .ZN(new_n756));
  XNOR2_X1  g0556(.A(KEYINPUT33), .B(G317), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(KEYINPUT97), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(KEYINPUT97), .B2(new_n757), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n745), .A2(new_n751), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G159), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n749), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT32), .Z(new_n763));
  INV_X1    g0563(.A(new_n744), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n205), .ZN(new_n765));
  INV_X1    g0565(.A(new_n740), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n556), .B1(new_n766), .B2(G77), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n767), .B1(new_n221), .B2(new_n737), .C1(new_n339), .C2(new_n756), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n728), .A2(new_n465), .B1(new_n733), .B2(new_n378), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n753), .A2(new_n204), .ZN(new_n770));
  OR4_X1    g0570(.A1(new_n765), .A2(new_n768), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n731), .A2(new_n760), .B1(new_n763), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n215), .B1(G20), .B2(new_n480), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n725), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n670), .A2(new_n556), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n775), .A2(G355), .B1(new_n591), .B2(new_n670), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n218), .A2(G45), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n245), .B2(G45), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n212), .A2(new_n389), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n722), .B1(new_n726), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n665), .B(new_n666), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n722), .ZN(G396));
  OAI22_X1  g0584(.A1(new_n764), .A2(new_n465), .B1(new_n548), .B2(new_n733), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n737), .A2(new_n583), .B1(new_n740), .B2(new_n591), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n556), .B1(new_n756), .B2(new_n787), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n785), .A2(new_n786), .A3(new_n770), .A4(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n729), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n789), .B1(new_n205), .B2(new_n790), .C1(new_n741), .C2(new_n749), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n764), .A2(new_n339), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n389), .B(new_n792), .C1(G58), .C2(new_n754), .ZN(new_n793));
  INV_X1    g0593(.A(G132), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n221), .B2(new_n790), .C1(new_n794), .C2(new_n749), .ZN(new_n795));
  INV_X1    g0595(.A(new_n737), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(G137), .B1(new_n766), .B2(G159), .ZN(new_n797));
  INV_X1    g0597(.A(G143), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n797), .B1(new_n798), .B2(new_n733), .C1(new_n253), .C2(new_n756), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT34), .Z(new_n800));
  OAI21_X1  g0600(.A(new_n791), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n773), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n773), .A2(new_n723), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n722), .B1(new_n223), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n331), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n333), .B1(new_n805), .B2(new_n328), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n321), .A2(new_n652), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n336), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n336), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n652), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n802), .B(new_n804), .C1(new_n811), .C2(new_n724), .ZN(new_n812));
  INV_X1    g0612(.A(new_n808), .ZN(new_n813));
  INV_X1    g0613(.A(new_n810), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n715), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n811), .B(new_n714), .C1(new_n626), .C2(new_n637), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(new_n702), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n702), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n722), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n812), .B1(new_n820), .B2(new_n822), .ZN(G384));
  NAND3_X1  g0623(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT35), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n826), .A2(G116), .A3(new_n216), .A4(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT36), .Z(new_n829));
  OR3_X1    g0629(.A1(new_n217), .A2(new_n223), .A3(new_n379), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n221), .A2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n208), .B(G13), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n366), .B(new_n376), .C1(new_n348), .C2(new_n714), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n359), .A2(new_n348), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n362), .A2(KEYINPUT72), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n363), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n375), .B(new_n652), .C1(new_n837), .C2(new_n374), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n817), .B2(new_n814), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT99), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n427), .A2(new_n430), .ZN(new_n844));
  INV_X1    g0644(.A(new_n650), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n430), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g0646(.A1(new_n843), .A2(new_n844), .A3(new_n846), .A4(new_n422), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT98), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n848), .B(new_n263), .C1(new_n394), .C2(KEYINPUT16), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n395), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n389), .A2(new_n392), .A3(new_n209), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n392), .B1(new_n389), .B2(new_n209), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n851), .A2(new_n852), .A3(new_n339), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n407), .B1(new_n853), .B2(new_n382), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n848), .B1(new_n854), .B2(new_n263), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n429), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n427), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n845), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n422), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n847), .B1(new_n859), .B2(KEYINPUT37), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n437), .A2(new_n845), .A3(new_n856), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n842), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n437), .A2(new_n845), .A3(new_n856), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n856), .A2(new_n845), .B1(new_n411), .B2(new_n421), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n843), .B1(new_n864), .B2(new_n857), .ZN(new_n865));
  OAI211_X1 g0665(.A(KEYINPUT38), .B(new_n863), .C1(new_n865), .C2(new_n847), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n841), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n862), .A2(new_n841), .A3(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n840), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n376), .A2(new_n652), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n844), .A2(new_n846), .A3(new_n422), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n844), .A2(new_n846), .A3(new_n843), .A4(new_n422), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n411), .A2(new_n650), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n872), .A2(new_n873), .B1(new_n437), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n866), .B1(new_n875), .B2(KEYINPUT38), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n862), .B2(new_n866), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n870), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n641), .A2(new_n845), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n869), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n438), .A2(new_n713), .A3(new_n717), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n645), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n882), .B(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n699), .A2(new_n700), .B1(new_n696), .B2(new_n677), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n886), .A2(new_n839), .A3(new_n815), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n868), .B2(new_n867), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n876), .A2(KEYINPUT40), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n888), .A2(new_n889), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n439), .A2(new_n886), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n885), .B1(new_n893), .B2(new_n666), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n208), .B2(new_n720), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n885), .A2(new_n893), .A3(new_n666), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n833), .B1(new_n895), .B2(new_n896), .ZN(G367));
  INV_X1    g0697(.A(new_n722), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n774), .B1(new_n212), .B2(new_n317), .C1(new_n241), .C2(new_n779), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n729), .A2(KEYINPUT46), .A3(G116), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n750), .A2(G317), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n744), .A2(G97), .ZN(new_n903));
  INV_X1    g0703(.A(new_n756), .ZN(new_n904));
  AOI22_X1  g0704(.A1(G294), .A2(new_n904), .B1(new_n766), .B2(G283), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n901), .A2(new_n902), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n737), .A2(new_n741), .B1(new_n733), .B2(new_n583), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT105), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n728), .A2(new_n591), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n389), .B1(new_n205), .B2(new_n753), .C1(new_n909), .C2(KEYINPUT46), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n906), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n283), .B1(new_n764), .B2(new_n223), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n753), .A2(new_n339), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n733), .A2(new_n253), .B1(new_n740), .B2(new_n221), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n728), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n916), .A2(G58), .B1(new_n904), .B2(G159), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n798), .B2(new_n737), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(G137), .B2(new_n750), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n911), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT47), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n773), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(KEYINPUT47), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n475), .A2(new_n714), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n628), .A2(new_n924), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n486), .A2(new_n925), .B1(new_n926), .B2(KEYINPUT100), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(KEYINPUT100), .B2(new_n926), .ZN(new_n928));
  INV_X1    g0728(.A(new_n725), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n900), .B1(new_n922), .B2(new_n923), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n507), .A2(new_n508), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n706), .B(new_n707), .C1(new_n931), .C2(new_n714), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n631), .A2(new_n652), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n539), .B1(new_n935), .B2(new_n614), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n714), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n660), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n938), .A2(KEYINPUT103), .A3(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT103), .B1(new_n938), .B2(KEYINPUT42), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n928), .B(KEYINPUT101), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT43), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n945), .A2(KEYINPUT102), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(KEYINPUT102), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n942), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n948), .B1(new_n942), .B2(new_n949), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n935), .A2(new_n668), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT104), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n671), .B(KEYINPUT41), .Z(new_n958));
  OR3_X1    g0758(.A1(new_n662), .A2(KEYINPUT44), .A3(new_n934), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT44), .B1(new_n662), .B2(new_n934), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n662), .A2(new_n934), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT45), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(new_n667), .A3(new_n658), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n667), .B(new_n658), .ZN(new_n967));
  INV_X1    g0767(.A(new_n659), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n660), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n961), .A2(new_n964), .A3(new_n668), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n718), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n958), .B1(new_n971), .B2(new_n718), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n721), .A2(G1), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n957), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n954), .B1(new_n951), .B2(new_n952), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n955), .B2(new_n956), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n930), .B1(new_n974), .B2(new_n976), .ZN(G387));
  OR2_X1    g0777(.A1(new_n658), .A2(new_n929), .ZN(new_n978));
  INV_X1    g0778(.A(new_n673), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n775), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(G107), .B2(new_n212), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n238), .A2(G45), .ZN(new_n982));
  AOI211_X1 g0782(.A(G45), .B(new_n979), .C1(G68), .C2(G77), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n257), .A2(G50), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT50), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n779), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n981), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n774), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n898), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n903), .B1(new_n221), .B2(new_n733), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n753), .A2(new_n317), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n990), .A2(new_n991), .A3(new_n389), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n750), .A2(G150), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n737), .A2(new_n761), .B1(new_n740), .B2(new_n339), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n728), .A2(new_n223), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n258), .A2(new_n904), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n992), .A2(new_n993), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n389), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n744), .B2(G116), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n753), .A2(new_n787), .B1(new_n728), .B2(new_n548), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n796), .A2(G322), .B1(new_n766), .B2(G303), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n741), .B2(new_n756), .C1(new_n1003), .C2(new_n733), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT106), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1001), .B1(new_n1005), .B2(KEYINPUT48), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT48), .B2(new_n1005), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT49), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1000), .B1(new_n738), .B2(new_n749), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n998), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n989), .B1(new_n1011), .B2(new_n773), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n969), .A2(new_n973), .B1(new_n978), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n969), .A2(new_n718), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n671), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n969), .A2(new_n718), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(G393));
  INV_X1    g0817(.A(KEYINPUT107), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n970), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n970), .A2(new_n1018), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1019), .A2(new_n966), .A3(new_n973), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n250), .A2(new_n779), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n774), .B1(new_n204), .B2(new_n212), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n898), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n283), .B(new_n765), .C1(G116), .C2(new_n754), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n916), .A2(G283), .B1(new_n904), .B2(G303), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n548), .C2(new_n740), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n737), .A2(new_n1003), .B1(new_n733), .B2(new_n741), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n734), .B2(new_n749), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n737), .A2(new_n253), .B1(new_n733), .B2(new_n761), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n764), .A2(new_n465), .B1(new_n221), .B2(new_n756), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n728), .A2(new_n339), .B1(new_n740), .B2(new_n257), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n999), .B1(new_n223), .B2(new_n753), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n798), .B2(new_n749), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1027), .A2(new_n1031), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1024), .B1(new_n1040), .B2(new_n773), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n934), .B2(new_n929), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1021), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1019), .A2(new_n966), .A3(new_n1020), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1014), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n971), .A2(new_n671), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(G390));
  OR2_X1    g0848(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n879), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n840), .C2(new_n870), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n834), .A2(new_n838), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n702), .A2(new_n811), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n707), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n624), .A2(new_n486), .A3(new_n579), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT93), .B1(new_n537), .B2(new_n539), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n709), .A2(new_n710), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n629), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n714), .B(new_n813), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1060), .A2(KEYINPUT110), .A3(new_n814), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT110), .B1(new_n1060), .B2(new_n814), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1061), .A2(new_n1062), .A3(new_n839), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n870), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n876), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1051), .B(new_n1053), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1062), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1060), .A2(KEYINPUT110), .A3(new_n814), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n1052), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1065), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n715), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n810), .B1(new_n1071), .B2(new_n811), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1064), .B1(new_n1072), .B2(new_n839), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n877), .A2(new_n879), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1069), .A2(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n701), .A2(new_n688), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(G330), .A3(new_n811), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n839), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1066), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n438), .A2(G330), .A3(new_n1076), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n883), .A2(new_n1081), .A3(new_n645), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1072), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1052), .B1(new_n702), .B2(new_n811), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n839), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1086), .B(new_n1053), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1082), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1080), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1066), .B(new_n1088), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n671), .A3(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1066), .B(new_n973), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n803), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n898), .B1(new_n258), .B2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n283), .B1(new_n761), .B2(new_n753), .C1(new_n764), .C2(new_n221), .ZN(new_n1096));
  INV_X1    g0896(.A(G137), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n794), .A2(new_n733), .B1(new_n756), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n737), .A2(new_n1099), .B1(new_n740), .B2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1096), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n728), .A2(new_n253), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT53), .ZN(new_n1104));
  INV_X1    g0904(.A(G125), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1102), .B(new_n1104), .C1(new_n1105), .C2(new_n749), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G294), .A2(new_n750), .B1(new_n729), .B2(G87), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n792), .A2(new_n283), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n756), .A2(new_n205), .B1(new_n740), .B2(new_n204), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G283), .B2(new_n796), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n753), .A2(new_n223), .B1(new_n733), .B2(new_n591), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT111), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1106), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1095), .B1(new_n1114), .B2(new_n773), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1074), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n724), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1092), .A2(new_n1093), .A3(new_n1117), .ZN(G378));
  INV_X1    g0918(.A(KEYINPUT120), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1082), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1091), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT57), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n890), .A2(new_n887), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1076), .A2(new_n811), .A3(new_n1052), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n873), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT38), .B1(new_n1126), .B2(new_n863), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n866), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT99), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n862), .A2(new_n841), .A3(new_n866), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1124), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(G330), .B(new_n1123), .C1(new_n1131), .C2(KEYINPUT40), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT115), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n275), .A2(new_n650), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n310), .B2(new_n314), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n313), .B(new_n1136), .C1(new_n304), .C2(new_n309), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n281), .A2(new_n303), .A3(KEYINPUT10), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n314), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1136), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n310), .A2(new_n314), .A3(new_n1137), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n1145), .A3(new_n1134), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1132), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT116), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1140), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n891), .A2(G330), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n882), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1149), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1119), .B1(new_n1122), .B2(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1132), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1147), .B1(new_n891), .B2(G330), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n882), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1149), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1165), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n1121), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1159), .A2(new_n671), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(KEYINPUT118), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT118), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1157), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1164), .A2(KEYINPUT119), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT119), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1149), .A2(new_n1154), .A3(new_n1172), .A4(new_n1155), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT57), .B1(new_n1174), .B2(new_n1121), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1167), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n722), .B1(new_n221), .B2(new_n803), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT114), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n744), .A2(G58), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT112), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n756), .A2(new_n204), .B1(new_n740), .B2(new_n317), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n737), .A2(new_n591), .B1(new_n733), .B2(new_n205), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n913), .A2(new_n995), .A3(new_n999), .A4(G41), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n787), .C2(new_n749), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT113), .B(KEYINPUT58), .Z(new_n1187));
  OAI22_X1  g0987(.A1(new_n737), .A2(new_n1105), .B1(new_n756), .B2(new_n794), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1100), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n733), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n916), .A2(new_n1189), .B1(new_n1190), .B2(G128), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1097), .B2(new_n740), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1188), .B(new_n1192), .C1(G150), .C2(new_n754), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n750), .A2(G124), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n744), .C2(G159), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1186), .A2(new_n1187), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G41), .B1(new_n999), .B2(G33), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1200), .B1(G50), .B2(new_n1201), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1178), .B1(new_n1202), .B2(new_n773), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1153), .B2(new_n724), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT117), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1174), .B2(new_n973), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1176), .A2(new_n1206), .ZN(G375));
  NAND2_X1  g1007(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n839), .A2(new_n723), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n790), .A2(new_n761), .B1(new_n749), .B2(new_n1099), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G137), .A2(new_n1190), .B1(new_n904), .B2(new_n1189), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n389), .B1(new_n754), .B2(G50), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n253), .C2(new_n740), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n796), .A2(G132), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT121), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1210), .A2(new_n1181), .A3(new_n1213), .A4(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n790), .A2(new_n204), .B1(new_n749), .B2(new_n583), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n796), .A2(G294), .B1(new_n766), .B2(G107), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n591), .B2(new_n756), .C1(new_n787), .C2(new_n733), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n556), .B1(new_n764), .B2(new_n223), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1217), .A2(new_n991), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n773), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n898), .C1(G68), .C2(new_n1094), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT122), .Z(new_n1224));
  AOI22_X1  g1024(.A1(new_n1208), .A2(new_n973), .B1(new_n1209), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n958), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1089), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1208), .A2(new_n1120), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1225), .B1(new_n1227), .B2(new_n1228), .ZN(G381));
  INV_X1    g1029(.A(G375), .ZN(new_n1230));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1047), .B(new_n930), .C1(new_n976), .C2(new_n974), .ZN(new_n1232));
  OR2_X1    g1032(.A1(G393), .A2(G396), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1232), .A2(G384), .A3(G381), .A4(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1230), .A2(new_n1231), .A3(new_n1234), .ZN(G407));
  NAND2_X1  g1035(.A1(new_n651), .A2(G213), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1230), .A2(new_n1231), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(new_n1238), .A3(G213), .ZN(G409));
  NAND2_X1  g1039(.A1(G387), .A2(G390), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(G396), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1240), .A2(new_n1232), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1240), .B2(new_n1232), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G378), .B(new_n1206), .C1(new_n1167), .C2(new_n1175), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1174), .A2(new_n1226), .A3(new_n1121), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1205), .B1(new_n1165), .B2(new_n973), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1231), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1245), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1228), .B(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n671), .A3(new_n1089), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(G384), .A3(new_n1225), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G384), .B1(new_n1253), .B2(new_n1225), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1250), .A2(new_n1236), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT123), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1237), .B1(new_n1245), .B2(new_n1249), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT123), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1257), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT62), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1258), .A2(KEYINPUT62), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1250), .A2(new_n1236), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G2897), .B(new_n1237), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1256), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1237), .A2(G2897), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1254), .A3(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1264), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1244), .B1(new_n1263), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT124), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1259), .A2(new_n1275), .A3(new_n1276), .A4(new_n1262), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1242), .A2(new_n1243), .A3(KEYINPUT61), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1271), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1236), .A4(new_n1257), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1260), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1257), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1277), .A2(new_n1279), .A3(new_n1284), .ZN(new_n1285));
  AND4_X1   g1085(.A1(new_n1261), .A2(new_n1250), .A3(new_n1236), .A4(new_n1257), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1261), .B1(new_n1260), .B2(new_n1257), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1275), .B1(new_n1288), .B2(new_n1276), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1274), .B1(new_n1285), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1274), .B(KEYINPUT127), .C1(new_n1285), .C2(new_n1289), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(G405));
  XNOR2_X1  g1094(.A(new_n1244), .B(new_n1257), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(G375), .B(new_n1231), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1295), .B(new_n1296), .ZN(G402));
endmodule


