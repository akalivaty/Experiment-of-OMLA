//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n187), .B2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  INV_X1    g010(.A(G110), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n188), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(new_n199), .A2(KEYINPUT75), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(KEYINPUT75), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n204));
  XNOR2_X1  g018(.A(G125), .B(G140), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(KEYINPUT16), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n191), .A2(new_n192), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n195), .A2(new_n188), .A3(new_n196), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(G110), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n216));
  INV_X1    g030(.A(G140), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G125), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n203), .A2(G140), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n221), .B2(new_n216), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(new_n208), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n206), .A2(G146), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n215), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G137), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n226), .B(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n212), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n229), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n210), .B1(new_n200), .B2(new_n201), .ZN(new_n232));
  INV_X1    g046(.A(new_n225), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT73), .B(G902), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n230), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n230), .A2(new_n234), .A3(KEYINPUT25), .A4(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G217), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n235), .B2(G234), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n230), .A2(new_n234), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n245), .A2(G902), .A3(new_n242), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G472), .ZN(new_n249));
  NOR2_X1   g063(.A1(G237), .A2(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n187), .B2(G116), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT68), .A3(G119), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n258), .A2(G119), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT2), .B(G113), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n261), .B1(new_n257), .B2(new_n259), .ZN(new_n267));
  INV_X1    g081(.A(new_n264), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n263), .A2(new_n266), .A3(new_n264), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(G146), .C1(new_n189), .C2(KEYINPUT1), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n189), .A2(new_n208), .A3(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n274), .A2(new_n278), .A3(new_n275), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n280));
  XNOR2_X1  g094(.A(G143), .B(G146), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n208), .A2(G143), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n273), .A2(G146), .ZN(new_n285));
  AND4_X1   g099(.A1(new_n280), .A2(new_n282), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n277), .B(new_n279), .C1(new_n283), .C2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT11), .ZN(new_n288));
  INV_X1    g102(.A(G134), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(G137), .ZN(new_n290));
  INV_X1    g104(.A(G137), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT11), .A3(G134), .ZN(new_n292));
  INV_X1    g106(.A(G131), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n289), .A2(G137), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n290), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n289), .A2(G137), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n291), .A2(G134), .ZN(new_n297));
  OAI21_X1  g111(.A(G131), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n287), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(KEYINPUT0), .A2(G128), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n284), .A2(new_n285), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n281), .A2(KEYINPUT65), .A3(new_n302), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT64), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT0), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n189), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n302), .B1(new_n284), .B2(new_n285), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n305), .A2(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G131), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n295), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n272), .A2(new_n301), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n272), .A2(new_n301), .A3(KEYINPUT70), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n313), .A2(new_n316), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n274), .A2(new_n278), .A3(new_n275), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n278), .B1(new_n274), .B2(new_n275), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT66), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n281), .A2(new_n280), .A3(new_n282), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n299), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT30), .B1(new_n323), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n301), .A2(new_n333), .A3(new_n317), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n272), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n255), .B1(new_n322), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n318), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n254), .B(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n341));
  INV_X1    g155(.A(new_n272), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n323), .B2(new_n331), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n320), .A2(new_n343), .A3(new_n321), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n338), .B(new_n341), .C1(new_n344), .C2(new_n337), .ZN(new_n345));
  INV_X1    g159(.A(new_n338), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n320), .A2(new_n343), .A3(new_n321), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n255), .B(new_n346), .C1(new_n347), .C2(KEYINPUT28), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n336), .B(new_n345), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AOI211_X1 g164(.A(KEYINPUT74), .B(new_n249), .C1(new_n350), .C2(new_n235), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n336), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n346), .B1(new_n347), .B2(KEYINPUT28), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n349), .B1(new_n354), .B2(new_n254), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n235), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n352), .B1(new_n356), .B2(G472), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(G472), .A2(G902), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n323), .A2(new_n331), .A3(KEYINPUT30), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n333), .B1(new_n301), .B2(new_n317), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n342), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(new_n320), .A3(new_n321), .A4(new_n254), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT71), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n320), .A2(new_n321), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n366), .A2(KEYINPUT71), .A3(new_n362), .A4(new_n254), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n365), .A2(KEYINPUT31), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n340), .ZN(new_n369));
  OAI22_X1  g183(.A1(new_n354), .A2(new_n369), .B1(new_n363), .B2(KEYINPUT31), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n359), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT32), .ZN(new_n372));
  INV_X1    g186(.A(new_n359), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n338), .B1(new_n344), .B2(new_n337), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n322), .A2(new_n335), .A3(new_n255), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT31), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n374), .A2(new_n340), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n365), .A2(KEYINPUT31), .A3(new_n367), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n372), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n248), .B1(new_n358), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G475), .A2(G902), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n222), .A2(new_n208), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n227), .A3(G214), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(new_n273), .ZN(new_n388));
  AOI21_X1  g202(.A(G143), .B1(new_n250), .B2(G214), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT17), .B(G131), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n385), .A2(new_n207), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G131), .B1(new_n388), .B2(new_n389), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n273), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n250), .A2(G143), .A3(G214), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n293), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT91), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n399), .A3(new_n393), .A4(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT18), .B(G131), .C1(new_n388), .C2(new_n389), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n221), .A2(G146), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n209), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT18), .A2(G131), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n394), .A2(new_n395), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(G113), .B(G122), .Z(new_n408));
  XOR2_X1   g222(.A(KEYINPUT90), .B(G104), .Z(new_n409));
  XOR2_X1   g223(.A(new_n408), .B(new_n409), .Z(new_n410));
  NAND3_X1  g224(.A1(new_n401), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n392), .A2(new_n396), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT19), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n205), .B(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n412), .B(new_n207), .C1(G146), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n407), .ZN(new_n416));
  INV_X1    g230(.A(new_n410), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n411), .A2(KEYINPUT92), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT92), .B1(new_n411), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n384), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT20), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n411), .A2(new_n418), .ZN(new_n423));
  NOR3_X1   g237(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT93), .B(G475), .Z(new_n427));
  INV_X1    g241(.A(G902), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n401), .A2(new_n407), .A3(new_n410), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n410), .B1(new_n401), .B2(new_n407), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(new_n431), .B2(KEYINPUT94), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT94), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n433), .B(new_n428), .C1(new_n429), .C2(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  OR2_X1    g250(.A1(KEYINPUT77), .A2(G107), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT77), .A2(G107), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G122), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G116), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n258), .A2(G122), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n443), .A2(KEYINPUT14), .ZN(new_n445));
  INV_X1    g259(.A(G107), .ZN(new_n446));
  INV_X1    g260(.A(new_n442), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(KEYINPUT14), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n273), .A2(G128), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n189), .A2(G143), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT95), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G128), .B(G143), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT95), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n454), .A2(new_n456), .A3(new_n289), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n453), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(KEYINPUT95), .ZN(new_n459));
  AOI21_X1  g273(.A(G134), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n449), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n289), .B1(new_n454), .B2(new_n456), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n455), .A2(KEYINPUT13), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(G134), .C1(KEYINPUT13), .C2(new_n450), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n439), .A2(new_n443), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n462), .B(new_n464), .C1(new_n465), .C2(new_n444), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT9), .B(G234), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n467), .A2(new_n241), .A3(G953), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n461), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n461), .B2(new_n466), .ZN(new_n470));
  OAI211_X1 g284(.A(KEYINPUT96), .B(new_n235), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G478), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(KEYINPUT15), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n461), .A2(new_n466), .ZN(new_n475));
  INV_X1    g289(.A(new_n468), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n461), .A2(new_n466), .A3(new_n468), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n473), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(KEYINPUT96), .A3(new_n235), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n436), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G113), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(new_n261), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT5), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n263), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n267), .A2(new_n268), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT79), .ZN(new_n491));
  INV_X1    g305(.A(G104), .ZN(new_n492));
  AND2_X1   g306(.A1(KEYINPUT77), .A2(G107), .ZN(new_n493));
  NOR2_X1   g307(.A1(KEYINPUT77), .A2(G107), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G101), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n491), .B1(G104), .B2(new_n446), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n493), .A2(new_n494), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n492), .A2(KEYINPUT3), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n446), .A2(G104), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT3), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n446), .B2(G104), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n495), .A2(new_n499), .B1(new_n505), .B2(new_n496), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n490), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G122), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT83), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n509), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT8), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n514), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n485), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n267), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n518), .A2(new_n486), .B1(new_n267), .B2(new_n268), .ZN(new_n519));
  AOI21_X1  g333(.A(G104), .B1(new_n437), .B2(new_n438), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n502), .A2(KEYINPUT79), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n495), .B(G101), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n501), .A2(new_n437), .A3(new_n438), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n504), .A2(new_n502), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n496), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n507), .A2(new_n516), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT88), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n507), .A2(new_n516), .A3(new_n530), .A4(new_n527), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n312), .A2(new_n311), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT65), .B1(new_n281), .B2(new_n302), .ZN(new_n534));
  AND4_X1   g348(.A1(KEYINPUT65), .A2(new_n284), .A3(new_n285), .A4(new_n302), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n536), .A2(KEYINPUT85), .A3(G125), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT85), .B1(new_n536), .B2(G125), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT86), .B1(new_n287), .B2(G125), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT86), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n326), .A2(new_n541), .A3(new_n330), .A4(new_n203), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n227), .A2(G224), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT87), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT78), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n505), .B2(new_n496), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT4), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n551), .B1(new_n505), .B2(new_n496), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n496), .B1(new_n523), .B2(new_n524), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT78), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n551), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n271), .A3(new_n270), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n506), .A2(new_n519), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n512), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n539), .A2(new_n543), .A3(KEYINPUT7), .A4(new_n546), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n532), .A2(new_n548), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n428), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n564));
  INV_X1    g378(.A(new_n512), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT84), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n512), .B1(new_n557), .B2(new_n558), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT84), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n564), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n568), .A2(new_n564), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n567), .A2(new_n570), .B1(new_n571), .B2(new_n559), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n544), .A2(new_n546), .ZN(new_n573));
  INV_X1    g387(.A(new_n546), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n539), .B2(new_n543), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n562), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G210), .B1(G237), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT89), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n561), .A2(new_n428), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n563), .A2(new_n565), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT6), .A3(new_n559), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n568), .A2(new_n569), .A3(new_n564), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n569), .B1(new_n568), .B2(new_n564), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n576), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n580), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n581), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n227), .A2(G952), .ZN(new_n592));
  INV_X1    g406(.A(G234), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(new_n593), .B2(new_n386), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n227), .B(new_n235), .C1(G234), .C2(G237), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT21), .B(G898), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G214), .B1(G237), .B2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n483), .A2(new_n591), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G469), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n274), .B(new_n275), .C1(new_n283), .C2(new_n286), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n506), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n276), .B1(new_n328), .B2(new_n329), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n526), .A2(new_n608), .A3(KEYINPUT80), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  INV_X1    g425(.A(new_n316), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT81), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(new_n604), .C1(new_n607), .C2(new_n609), .ZN(new_n614));
  OAI211_X1 g428(.A(KEYINPUT4), .B(new_n525), .C1(new_n553), .C2(KEYINPUT78), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n505), .A2(new_n549), .A3(new_n496), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n313), .B(new_n556), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n506), .A2(KEYINPUT10), .A3(new_n287), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n611), .A2(new_n612), .A3(new_n614), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(G110), .B(G140), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n227), .A2(G227), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n506), .A2(new_n287), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n506), .A2(new_n605), .A3(new_n606), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT80), .B1(new_n526), .B2(new_n608), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT12), .B1(new_n628), .B2(new_n612), .ZN(new_n629));
  OR3_X1    g443(.A1(new_n628), .A2(KEYINPUT12), .A3(new_n612), .ZN(new_n630));
  AND4_X1   g444(.A1(new_n620), .A2(new_n624), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n619), .A2(new_n614), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n626), .A2(new_n627), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n613), .B1(new_n633), .B2(new_n604), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n316), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n624), .B1(new_n635), .B2(new_n620), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n603), .B(new_n235), .C1(new_n631), .C2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n603), .A2(new_n428), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n635), .A2(new_n620), .A3(new_n624), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n620), .A2(new_n629), .A3(new_n630), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n623), .B(KEYINPUT76), .ZN(new_n642));
  OAI211_X1 g456(.A(G469), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n637), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(G221), .B1(new_n467), .B2(G902), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n602), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n383), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT97), .B(G101), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G3));
  INV_X1    g464(.A(new_n235), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n377), .B2(new_n378), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n371), .B(new_n247), .C1(new_n652), .C2(new_n249), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n644), .A2(new_n645), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT98), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n646), .B2(new_n653), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n599), .B1(new_n577), .B2(new_n579), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n582), .A2(new_n587), .A3(new_n579), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n600), .B1(new_n588), .B2(new_n578), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n577), .A2(new_n579), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(KEYINPUT99), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n598), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n432), .A2(new_n434), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n421), .A2(KEYINPUT20), .B1(new_n423), .B2(new_n424), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT33), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n475), .B2(KEYINPUT100), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n479), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n469), .A2(new_n470), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n672), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n676), .A3(G478), .A4(new_n235), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n472), .B1(new_n675), .B2(new_n651), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n670), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n663), .A2(new_n666), .A3(new_n667), .A4(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n659), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT34), .B(G104), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G6));
  NAND2_X1  g498(.A1(new_n663), .A2(new_n666), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n598), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT20), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n687), .B(new_n384), .C1(new_n419), .C2(new_n420), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n422), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n689), .A2(new_n435), .A3(new_n482), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n659), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT35), .B(G107), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  OR2_X1    g508(.A1(new_n652), .A2(new_n249), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n371), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n212), .A2(new_n225), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n231), .A2(KEYINPUT36), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n242), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n428), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n243), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n696), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n647), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  NAND3_X1  g521(.A1(new_n644), .A2(new_n645), .A3(new_n702), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n579), .B1(new_n582), .B2(new_n587), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n662), .A2(new_n709), .A3(new_n660), .A4(new_n600), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT99), .B1(new_n664), .B2(new_n665), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n596), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(G900), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n594), .B(KEYINPUT101), .Z(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n690), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n358), .B2(new_n382), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G128), .ZN(G30));
  XOR2_X1   g535(.A(new_n716), .B(KEYINPUT39), .Z(new_n722));
  NAND2_X1  g536(.A1(new_n655), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT106), .Z(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT40), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n591), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(G472), .A2(G902), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT103), .B1(new_n344), .B2(new_n369), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n347), .A2(new_n730), .A3(new_n340), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(G472), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n365), .A2(new_n367), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n728), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT104), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(new_n728), .C1(new_n732), .C2(new_n733), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n377), .A2(new_n378), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n380), .B1(new_n738), .B2(new_n359), .ZN(new_n739));
  AOI211_X1 g553(.A(KEYINPUT32), .B(new_n373), .C1(new_n377), .C2(new_n378), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n735), .B(new_n737), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n436), .A2(new_n482), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n702), .A2(new_n600), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n727), .A2(new_n741), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(KEYINPUT105), .Z(new_n746));
  NAND2_X1  g560(.A1(new_n724), .A2(KEYINPUT40), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n725), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G143), .ZN(G45));
  NAND2_X1  g563(.A1(new_n677), .A2(new_n678), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n750), .B(new_n717), .C1(new_n668), .C2(new_n669), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n358), .B2(new_n382), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n712), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G146), .ZN(G48));
  OAI21_X1  g568(.A(KEYINPUT29), .B1(new_n374), .B2(new_n255), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n366), .A2(new_n362), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n354), .A2(new_n341), .B1(new_n756), .B2(new_n255), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n651), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT74), .B1(new_n758), .B2(new_n249), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n356), .A2(new_n352), .A3(G472), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n759), .B(new_n760), .C1(new_n739), .C2(new_n740), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n235), .B1(new_n631), .B2(new_n636), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(G469), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n763), .A2(new_n645), .A3(new_n637), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n247), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n765), .A2(new_n681), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT41), .B(G113), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G15));
  NAND4_X1  g582(.A1(new_n686), .A2(new_n383), .A3(new_n690), .A4(new_n764), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G116), .ZN(G18));
  NAND3_X1  g584(.A1(new_n764), .A2(new_n663), .A3(new_n666), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n483), .A2(new_n667), .A3(new_n702), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n382), .B2(new_n358), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G119), .ZN(G21));
  NOR3_X1   g590(.A1(new_n653), .A2(new_n598), .A3(new_n742), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  INV_X1    g593(.A(new_n751), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n695), .A2(new_n780), .A3(new_n371), .A4(new_n702), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT107), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n710), .A2(new_n711), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n652), .A2(new_n249), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n784), .A2(new_n751), .A3(new_n379), .A4(new_n703), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n783), .A2(new_n785), .A3(new_n786), .A4(new_n764), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G125), .ZN(G27));
  NAND4_X1  g603(.A1(new_n581), .A2(new_n590), .A3(new_n645), .A4(new_n599), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n637), .A2(new_n639), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT108), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n640), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n635), .A2(KEYINPUT108), .A3(new_n620), .A4(new_n624), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n641), .A2(new_n642), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(G469), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n761), .A2(new_n247), .A3(new_n791), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT109), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT42), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n751), .A2(KEYINPUT109), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT109), .B(KEYINPUT42), .C1(new_n800), .C2(new_n751), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT110), .B(G131), .Z(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G33));
  AOI21_X1  g622(.A(new_n790), .B1(new_n792), .B2(new_n798), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n383), .A2(new_n690), .A3(new_n717), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G134), .ZN(G36));
  NAND2_X1  g625(.A1(new_n670), .A2(new_n750), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT43), .Z(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n696), .A3(new_n702), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n581), .A2(new_n590), .A3(new_n599), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n813), .A2(KEYINPUT44), .A3(new_n696), .A4(new_n702), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n797), .A2(new_n640), .ZN(new_n821));
  OAI21_X1  g635(.A(G469), .B1(new_n821), .B2(KEYINPUT45), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT45), .ZN(new_n823));
  OAI211_X1 g637(.A(KEYINPUT46), .B(new_n639), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n637), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT111), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n822), .A2(new_n823), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n639), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT46), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n825), .A2(KEYINPUT111), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n722), .A2(new_n645), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n820), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G137), .ZN(G39));
  XNOR2_X1  g649(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n831), .A2(new_n830), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n825), .A2(KEYINPUT111), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n645), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n832), .A2(new_n645), .A3(new_n836), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n761), .A2(new_n247), .A3(new_n751), .A4(new_n817), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(G140), .ZN(G42));
  NAND2_X1  g660(.A1(new_n763), .A2(new_n637), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT49), .ZN(new_n848));
  INV_X1    g662(.A(new_n812), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n247), .A3(new_n645), .A4(new_n599), .ZN(new_n850));
  OR4_X1    g664(.A1(new_n727), .A2(new_n848), .A3(new_n741), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n813), .A2(new_n715), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n653), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n592), .B1(new_n854), .B2(new_n771), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n764), .A2(new_n818), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n856), .A2(new_n741), .A3(new_n248), .A4(new_n594), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n680), .B2(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n852), .A2(new_n856), .ZN(new_n859));
  INV_X1    g673(.A(new_n383), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT48), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(KEYINPUT117), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(KEYINPUT117), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n861), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n727), .A2(new_n599), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n853), .A2(new_n764), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT50), .Z(new_n869));
  NOR2_X1   g683(.A1(new_n436), .A2(new_n750), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n857), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n704), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n869), .B(new_n871), .C1(new_n872), .C2(new_n859), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n832), .A2(new_n645), .A3(new_n836), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n836), .B1(new_n832), .B2(new_n645), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n874), .A2(new_n875), .B1(new_n645), .B2(new_n847), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n854), .A2(new_n817), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n858), .B(new_n866), .C1(new_n878), .C2(KEYINPUT51), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(KEYINPUT51), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n702), .A2(new_n841), .A3(new_n716), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n741), .A2(new_n799), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n685), .A2(new_n742), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n883), .A2(new_n884), .B1(new_n712), .B2(new_n752), .ZN(new_n885));
  AND4_X1   g699(.A1(KEYINPUT52), .A2(new_n885), .A3(new_n788), .A4(new_n720), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n782), .A2(new_n787), .B1(new_n712), .B2(new_n719), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT52), .B1(new_n887), .B2(new_n885), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n804), .A2(new_n805), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n474), .A2(new_n481), .A3(new_n717), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n434), .B2(new_n432), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n702), .A2(new_n892), .A3(new_n689), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n581), .A3(new_n590), .A4(new_n599), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n382), .B2(new_n358), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n895), .A2(new_n655), .B1(new_n785), .B2(new_n809), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n647), .B1(new_n383), .B2(new_n704), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n591), .A2(new_n601), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n426), .A2(new_n435), .A3(new_n482), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT113), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n899), .A2(KEYINPUT113), .B1(new_n436), .B2(new_n750), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n656), .A2(new_n902), .A3(new_n658), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n896), .A2(new_n897), .A3(new_n810), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n772), .B1(new_n774), .B2(new_n777), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n766), .A2(new_n769), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n890), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n881), .B1(new_n889), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n885), .A2(new_n788), .A3(KEYINPUT52), .A4(new_n720), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(KEYINPUT114), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n889), .B2(KEYINPUT114), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n907), .A2(KEYINPUT53), .A3(new_n805), .A4(new_n804), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT116), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n904), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n904), .A2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI22_X1  g731(.A1(KEYINPUT115), .A2(new_n909), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n885), .A2(new_n788), .A3(new_n720), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT52), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n910), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n766), .A2(new_n769), .A3(new_n906), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n806), .A2(new_n904), .A3(new_n924), .ZN(new_n925));
  AOI211_X1 g739(.A(KEYINPUT115), .B(KEYINPUT53), .C1(new_n923), .C2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n918), .A2(new_n919), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n881), .B1(new_n923), .B2(new_n925), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n908), .A2(KEYINPUT53), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n912), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n879), .A2(new_n880), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(G952), .A2(G953), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n851), .B1(new_n934), .B2(new_n935), .ZN(G75));
  AOI21_X1  g750(.A(KEYINPUT53), .B1(new_n923), .B2(new_n925), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT115), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n922), .A2(KEYINPUT114), .A3(new_n910), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n910), .A2(KEYINPUT114), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n806), .A2(new_n924), .A3(new_n881), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n905), .A2(KEYINPUT116), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n904), .A2(new_n914), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  OAI22_X1  g759(.A1(new_n937), .A2(new_n938), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n651), .B(new_n579), .C1(new_n946), .C2(new_n926), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n572), .B(KEYINPUT118), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(new_n576), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n952), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n947), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n227), .A2(G952), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT119), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT119), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n953), .A2(new_n960), .A3(new_n955), .A4(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(G51));
  XNOR2_X1  g776(.A(new_n638), .B(KEYINPUT57), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n919), .B1(new_n918), .B2(new_n927), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n946), .A2(KEYINPUT54), .A3(new_n926), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n631), .A2(new_n636), .ZN(new_n969));
  OAI211_X1 g783(.A(KEYINPUT120), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n235), .B1(new_n918), .B2(new_n927), .ZN(new_n972));
  INV_X1    g786(.A(new_n827), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n956), .B1(new_n971), .B2(new_n974), .ZN(G54));
  NAND3_X1  g789(.A1(new_n972), .A2(KEYINPUT58), .A3(G475), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n419), .A2(new_n420), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(new_n956), .ZN(G60));
  AND2_X1   g794(.A1(new_n674), .A2(new_n676), .ZN(new_n981));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT59), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n933), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n964), .A2(new_n965), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n981), .A2(new_n983), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n956), .B(new_n984), .C1(new_n985), .C2(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(new_n918), .A2(new_n927), .ZN(new_n988));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT121), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT60), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n245), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n988), .A2(new_n699), .A3(new_n991), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n993), .A2(new_n957), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n993), .A2(KEYINPUT61), .A3(new_n957), .A4(new_n994), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(G66));
  INV_X1    g813(.A(G224), .ZN(new_n1000));
  OAI21_X1  g814(.A(G953), .B1(new_n597), .B2(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n907), .A2(new_n903), .A3(new_n897), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n950), .B1(G898), .B2(new_n227), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT122), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(new_n1005), .ZN(G69));
  AND2_X1   g820(.A1(new_n884), .A2(new_n383), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n832), .A2(new_n833), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1008), .A2(new_n890), .A3(new_n810), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n874), .A2(new_n875), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n844), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n820), .A2(new_n832), .A3(new_n833), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n887), .A2(new_n753), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n834), .A2(KEYINPUT124), .A3(new_n753), .A4(new_n887), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1011), .A2(KEYINPUT125), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n1008), .A2(new_n890), .A3(new_n810), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1015), .A2(new_n845), .A3(new_n1018), .A4(new_n1016), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT125), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1017), .A2(new_n1021), .A3(new_n227), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n360), .A2(new_n361), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(new_n414), .Z(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(G900), .B2(G953), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n383), .A2(new_n818), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n723), .B(new_n1027), .C1(new_n900), .C2(new_n901), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1013), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n748), .A2(new_n753), .A3(new_n887), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n1029), .B(new_n845), .C1(KEYINPUT62), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT123), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1030), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1024), .B1(new_n1036), .B2(G953), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1026), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT126), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1024), .A2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g854(.A(new_n227), .B(new_n1040), .C1(G227), .C2(G900), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1041), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1026), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1042), .A2(new_n1044), .ZN(G72));
  XNOR2_X1  g859(.A(new_n728), .B(KEYINPUT63), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g861(.A(new_n336), .ZN(new_n1048));
  OAI211_X1 g862(.A(new_n931), .B(new_n1047), .C1(new_n733), .C2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1046), .B1(new_n1036), .B2(new_n1002), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n756), .A2(new_n254), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n1049), .B(new_n957), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1017), .A2(new_n1021), .A3(new_n1002), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1053), .A2(KEYINPUT127), .A3(new_n1047), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n756), .A2(new_n254), .ZN(new_n1055));
  AND2_X1   g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1053), .A2(new_n1047), .ZN(new_n1057));
  INV_X1    g871(.A(KEYINPUT127), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1052), .B1(new_n1056), .B2(new_n1059), .ZN(G57));
endmodule


