//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  AOI211_X1 g0017(.A(new_n215), .B(new_n217), .C1(G68), .C2(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n204), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n210), .B(new_n227), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AOI21_X1  g0048(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT68), .B(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G226), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  OAI22_X1  g0052(.A1(new_n250), .A2(new_n251), .B1(new_n219), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n249), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT13), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G41), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n260), .B(G274), .C1(new_n265), .C2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(G45), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n267), .B(KEYINPUT67), .C1(G1), .C2(new_n261), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  OAI211_X1 g0069(.A(G1), .B(G13), .C1(new_n269), .C2(new_n261), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(new_n260), .C1(G41), .C2(G45), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G238), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n258), .A2(new_n259), .A3(new_n266), .A4(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n257), .B1(new_n253), .B2(new_n254), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n274), .B(new_n266), .C1(new_n276), .C2(new_n270), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT76), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OR3_X1    g0080(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(G169), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT14), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n280), .A2(new_n281), .A3(new_n284), .A4(G169), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n275), .A2(new_n278), .A3(G179), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n203), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(G50), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n229), .A2(new_n269), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n269), .A2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n288), .B1(new_n289), .B2(new_n290), .C1(new_n292), .C2(new_n211), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n228), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT11), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n260), .B2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n299), .A2(KEYINPUT12), .A3(G68), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT12), .B1(new_n299), .B2(G68), .ZN(new_n301));
  AOI22_X1  g0101(.A1(G68), .A2(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n287), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n280), .A2(new_n281), .A3(G200), .ZN(new_n306));
  INV_X1    g0106(.A(new_n303), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n275), .A2(new_n278), .A3(G190), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n299), .A2(G50), .ZN(new_n312));
  INV_X1    g0112(.A(new_n298), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n289), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT72), .ZN(new_n315));
  INV_X1    g0115(.A(G150), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n290), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT8), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT71), .B1(new_n319), .B2(G58), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(G58), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT71), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n315), .B(new_n318), .C1(new_n325), .C2(new_n292), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n292), .B1(new_n322), .B2(new_n324), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT72), .B1(new_n327), .B2(new_n317), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n201), .B2(new_n204), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n312), .B(new_n314), .C1(new_n330), .C2(new_n295), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT75), .B1(new_n331), .B2(KEYINPUT9), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n312), .B1(new_n330), .B2(new_n295), .ZN(new_n333));
  INV_X1    g0133(.A(new_n314), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT9), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(KEYINPUT74), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G33), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n345), .B1(new_n349), .B2(new_n252), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n254), .A2(KEYINPUT69), .A3(G1698), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(G223), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(G77), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT68), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(new_n254), .A3(G222), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n352), .A2(KEYINPUT70), .A3(new_n353), .A4(new_n358), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n249), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n273), .A2(G226), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n364), .A2(new_n266), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n344), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n363), .A2(G190), .A3(new_n365), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(new_n337), .C2(new_n335), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT10), .B1(new_n340), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n331), .A2(KEYINPUT9), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n339), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n350), .A2(G238), .A3(new_n351), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n213), .B2(new_n254), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n349), .A2(new_n250), .A3(new_n219), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n249), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n273), .A2(G244), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n379), .A2(new_n266), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G20), .A2(G77), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT8), .B(G58), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT15), .B(G87), .ZN(new_n386));
  OAI221_X1 g0186(.A(new_n384), .B1(new_n385), .B2(new_n290), .C1(new_n292), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n299), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n387), .A2(new_n295), .B1(new_n211), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n211), .B2(new_n313), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n383), .B(new_n390), .C1(G169), .C2(new_n381), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n381), .A2(G190), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n379), .A2(new_n266), .A3(new_n380), .ZN(new_n393));
  INV_X1    g0193(.A(new_n344), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n311), .A2(new_n375), .A3(new_n391), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n254), .B2(G20), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n349), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n203), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G159), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n290), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G58), .A2(G68), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n229), .B1(new_n204), .B2(new_n404), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT77), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT16), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n254), .A2(new_n398), .A3(G20), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n349), .B2(new_n229), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n405), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT77), .B(new_n409), .C1(new_n414), .C2(new_n403), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n408), .A2(new_n415), .A3(new_n295), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n325), .A2(new_n299), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n325), .B2(new_n298), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT78), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n357), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n421), .A2(new_n349), .B1(new_n269), .B2(new_n220), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n249), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n273), .A2(G232), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n266), .ZN(new_n425));
  INV_X1    g0225(.A(G169), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n425), .A2(G179), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n420), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n431), .A2(KEYINPUT79), .ZN(new_n432));
  INV_X1    g0232(.A(G190), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n425), .A2(G200), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n416), .A2(new_n434), .A3(new_n419), .A4(new_n435), .ZN(new_n436));
  XOR2_X1   g0236(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n437));
  OR3_X1    g0237(.A1(new_n436), .A2(KEYINPUT81), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT81), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n420), .A2(KEYINPUT18), .A3(new_n427), .A4(new_n428), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n431), .A2(KEYINPUT79), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n363), .A2(new_n365), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G179), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n445), .A2(KEYINPUT73), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n426), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(KEYINPUT73), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n335), .A4(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n432), .A2(new_n441), .A3(new_n443), .A4(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n397), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n221), .B1(new_n354), .B2(new_n356), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n224), .A2(new_n252), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n254), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G294), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n270), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n260), .B(G45), .C1(new_n457), .C2(G41), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n262), .A2(new_n264), .A3(new_n457), .ZN(new_n460));
  AOI211_X1 g0260(.A(new_n214), .B(new_n249), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n460), .A3(G274), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n433), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n463), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT88), .B1(new_n456), .B2(new_n461), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT88), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n249), .B1(new_n459), .B2(new_n460), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G264), .ZN(new_n469));
  INV_X1    g0269(.A(new_n455), .ZN(new_n470));
  INV_X1    g0270(.A(new_n453), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n250), .B2(new_n221), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(new_n254), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n467), .B(new_n469), .C1(new_n473), .C2(new_n270), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n465), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n464), .B1(new_n475), .B2(G200), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n346), .A2(new_n348), .A3(new_n229), .A4(G87), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT22), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT22), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n254), .A2(new_n479), .A3(new_n229), .A4(G87), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n291), .A2(G116), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n229), .A2(G107), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT23), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n481), .A2(KEYINPUT24), .A3(new_n482), .A4(new_n484), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n295), .A3(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n294), .A2(new_n228), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n260), .A2(G33), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(new_n299), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G107), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n299), .A2(G107), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n495), .B(KEYINPUT25), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n489), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n476), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n489), .A2(new_n494), .A3(new_n496), .ZN(new_n499));
  AOI211_X1 g0299(.A(new_n382), .B(new_n465), .C1(new_n466), .C2(new_n474), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n426), .B1(new_n462), .B2(new_n463), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n291), .A2(G97), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT19), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n229), .B1(new_n256), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G97), .A2(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n220), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n254), .A2(new_n229), .A3(G68), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n490), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n492), .A2(new_n386), .ZN(new_n511));
  INV_X1    g0311(.A(new_n386), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n299), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G274), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n267), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n270), .A2(G250), .A3(new_n267), .ZN(new_n518));
  INV_X1    g0318(.A(G238), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n250), .A2(new_n519), .B1(new_n212), .B2(new_n252), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(new_n254), .B1(G33), .B2(G116), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n517), .B(new_n518), .C1(new_n521), .C2(new_n270), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n514), .B1(new_n523), .B2(new_n382), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n426), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n508), .A2(new_n509), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n295), .ZN(new_n527));
  INV_X1    g0327(.A(new_n513), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n493), .A2(G87), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n394), .B2(new_n522), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n521), .A2(new_n270), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(G190), .A3(new_n517), .A4(new_n518), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n524), .A2(new_n525), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n498), .A2(new_n502), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G264), .A2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n254), .B(new_n536), .C1(new_n250), .C2(new_n224), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n249), .C1(G303), .C2(new_n254), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n468), .A2(G270), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n463), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n426), .ZN(new_n542));
  INV_X1    g0342(.A(G116), .ZN(new_n543));
  OR3_X1    g0343(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT86), .B1(new_n492), .B2(new_n543), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n299), .A2(G116), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(G20), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n295), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n549), .B1(new_n295), .B2(new_n550), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G283), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n554), .B(new_n229), .C1(G33), .C2(new_n223), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT20), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(KEYINPUT20), .B(new_n555), .C1(new_n551), .C2(new_n552), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n546), .B(new_n548), .C1(new_n556), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n542), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n540), .A2(G200), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n541), .A2(G190), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n540), .A2(new_n382), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n542), .A2(new_n559), .A3(KEYINPUT21), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n562), .A2(new_n566), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n535), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n468), .A2(G257), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n463), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n357), .A2(new_n254), .A3(G244), .ZN(new_n574));
  XOR2_X1   g0374(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n357), .A2(new_n254), .A3(KEYINPUT4), .A4(G244), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n346), .A2(new_n348), .A3(G250), .A4(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n576), .A2(new_n554), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n573), .B1(new_n579), .B2(new_n249), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n290), .A2(new_n211), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n223), .A2(new_n213), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n506), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n582), .B1(new_n587), .B2(G20), .ZN(new_n588));
  OAI21_X1  g0388(.A(G107), .B1(new_n410), .B2(new_n411), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n490), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n299), .A2(G97), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n492), .A2(new_n223), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n578), .A2(new_n554), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n574), .B2(new_n575), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n270), .B1(new_n595), .B2(new_n577), .ZN(new_n596));
  OAI21_X1  g0396(.A(G200), .B1(new_n596), .B2(new_n573), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n581), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n579), .A2(new_n249), .ZN(new_n601));
  INV_X1    g0401(.A(new_n573), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(G179), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n426), .B2(new_n580), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n588), .A2(new_n589), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n591), .B1(new_n605), .B2(new_n295), .ZN(new_n606));
  INV_X1    g0406(.A(new_n592), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT84), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT84), .ZN(new_n609));
  NOR4_X1   g0409(.A1(new_n590), .A2(new_n609), .A3(new_n591), .A4(new_n592), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n604), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n581), .A2(new_n593), .A3(KEYINPUT83), .A4(new_n597), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n600), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT85), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n600), .A2(new_n611), .A3(new_n615), .A4(new_n612), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n451), .A2(new_n571), .A3(new_n614), .A4(new_n616), .ZN(G372));
  INV_X1    g0417(.A(KEYINPUT91), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n340), .A2(new_n369), .A3(KEYINPUT10), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n373), .B1(new_n372), .B2(new_n339), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n370), .A2(new_n374), .A3(KEYINPUT91), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n391), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n309), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n304), .A2(new_n625), .A3(KEYINPUT90), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT90), .B1(new_n304), .B2(new_n625), .ZN(new_n627));
  INV_X1    g0427(.A(new_n441), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n431), .A2(new_n442), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n623), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n449), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n524), .A2(new_n525), .ZN(new_n634));
  INV_X1    g0434(.A(new_n593), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n604), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n534), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n634), .B1(new_n638), .B2(KEYINPUT26), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT89), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT89), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n562), .A2(new_n642), .A3(new_n568), .A4(new_n569), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n502), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n476), .A2(new_n497), .ZN(new_n645));
  INV_X1    g0445(.A(new_n534), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n613), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n639), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT26), .B1(new_n646), .B2(new_n611), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n451), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n633), .A2(new_n651), .ZN(G369));
  INV_X1    g0452(.A(G13), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G20), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n260), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n498), .B(new_n502), .C1(new_n497), .C2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n502), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT93), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n640), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n502), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n661), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n570), .B(KEYINPUT92), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n563), .A2(new_n661), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n641), .A2(new_n643), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n673), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n665), .A3(G330), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n671), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n208), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n265), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G1), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n506), .A2(new_n220), .A3(new_n543), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n683), .A2(new_n684), .B1(new_n231), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n660), .B1(new_n648), .B2(new_n649), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n646), .A2(new_n611), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n689), .A2(new_n690), .B1(new_n525), .B2(new_n524), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n692));
  INV_X1    g0492(.A(new_n613), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n531), .A2(new_n533), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n498), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n640), .A2(new_n668), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n691), .B(new_n692), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .A3(new_n661), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n688), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT94), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n355), .A2(G1698), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n703));
  OAI21_X1  g0503(.A(G250), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n349), .B1(new_n704), .B2(new_n471), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n249), .B1(new_n705), .B2(new_n470), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n467), .B1(new_n706), .B2(new_n469), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n456), .A2(KEYINPUT88), .A3(new_n461), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n523), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n567), .A2(new_n580), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n701), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n463), .B1(new_n707), .B2(new_n708), .ZN(new_n712));
  INV_X1    g0512(.A(new_n580), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n522), .A2(new_n382), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n712), .A2(new_n540), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n522), .B1(new_n466), .B2(new_n474), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(KEYINPUT30), .A3(new_n567), .A4(new_n580), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n711), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT31), .B1(new_n718), .B2(new_n660), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n700), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n660), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(KEYINPUT94), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n571), .A2(new_n614), .A3(new_n616), .A4(new_n661), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n721), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n699), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n686), .B1(new_n731), .B2(G1), .ZN(G364));
  NAND2_X1  g0532(.A1(new_n677), .A2(G330), .ZN(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n674), .A2(new_n734), .A3(new_n676), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n654), .A2(G45), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n682), .A2(G1), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n228), .B1(G20), .B2(new_n426), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n229), .A2(new_n382), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT95), .Z(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n433), .A3(new_n341), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n742), .A2(G190), .A3(new_n341), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G311), .A2(new_n744), .B1(new_n746), .B2(G322), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n741), .A2(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n433), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G326), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(new_n349), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n229), .A2(G179), .A3(G190), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n341), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n751), .B1(G329), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n433), .A2(G179), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n229), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n748), .A2(G190), .ZN(new_n760));
  AND2_X1   g0560(.A1(KEYINPUT33), .A2(G317), .ZN(new_n761));
  NOR2_X1   g0561(.A1(KEYINPUT33), .A2(G317), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n759), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n394), .A2(new_n752), .ZN(new_n766));
  INV_X1    g0566(.A(G303), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n229), .A2(new_n433), .A3(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n394), .A2(new_n768), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n764), .B1(new_n765), .B2(new_n766), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n754), .A2(G159), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n774));
  INV_X1    g0574(.A(new_n758), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n773), .A2(KEYINPUT96), .B1(G97), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n766), .A2(new_n213), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n774), .A2(new_n776), .A3(new_n254), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n745), .A2(new_n202), .ZN(new_n780));
  INV_X1    g0580(.A(new_n760), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n203), .ZN(new_n782));
  INV_X1    g0582(.A(new_n769), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G87), .ZN(new_n784));
  INV_X1    g0584(.A(new_n749), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n784), .B1(new_n289), .B2(new_n785), .C1(new_n743), .C2(new_n211), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n779), .A2(new_n780), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT97), .Z(new_n788));
  AOI21_X1  g0588(.A(new_n740), .B1(new_n770), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n739), .ZN(new_n793));
  INV_X1    g0593(.A(G45), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n232), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n680), .A2(new_n254), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(new_n247), .C2(new_n794), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n254), .A2(G355), .A3(new_n208), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n797), .B(new_n798), .C1(G116), .C2(new_n208), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n789), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n792), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n677), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n738), .B1(new_n802), .B2(new_n737), .ZN(G396));
  AOI22_X1  g0603(.A1(new_n392), .A2(new_n395), .B1(new_n390), .B2(new_n660), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n624), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n391), .A2(new_n660), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n687), .B(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(new_n729), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n737), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n781), .A2(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n781), .A2(KEYINPUT98), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n766), .A2(new_n220), .B1(new_n816), .B2(new_n753), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n815), .A2(new_n765), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n254), .B(new_n819), .C1(G303), .C2(new_n749), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n744), .A2(G116), .B1(G107), .B2(new_n783), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n756), .B2(new_n745), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n818), .B2(new_n817), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n820), .B(new_n823), .C1(new_n223), .C2(new_n758), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G143), .A2(new_n746), .B1(new_n744), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n825), .B1(new_n826), .B2(new_n785), .C1(new_n316), .C2(new_n781), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT34), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n758), .A2(new_n202), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n349), .B1(new_n754), .B2(G132), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT101), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n289), .A2(new_n769), .B1(new_n766), .B2(new_n203), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n829), .B(new_n832), .C1(new_n833), .C2(KEYINPUT100), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n828), .B(new_n834), .C1(KEYINPUT100), .C2(new_n833), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n830), .A2(new_n831), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n824), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n739), .ZN(new_n839));
  INV_X1    g0639(.A(new_n737), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n809), .A2(new_n790), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n739), .A2(new_n790), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n211), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n812), .A2(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n719), .A2(new_n720), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n727), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n451), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n658), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n420), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n628), .B2(new_n631), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n429), .A2(new_n436), .A3(new_n850), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n429), .A2(new_n850), .A3(KEYINPUT37), .A4(new_n436), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n855), .A2(KEYINPUT103), .A3(new_n856), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n432), .A2(new_n441), .A3(new_n443), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n851), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n867), .A3(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n809), .B1(new_n846), .B2(new_n727), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n307), .A2(new_n661), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n304), .A2(new_n309), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n287), .A2(new_n303), .A3(new_n660), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT40), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n865), .B2(new_n867), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n868), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n877), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n848), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g0685(.A(KEYINPUT40), .B(new_n876), .C1(new_n881), .C2(new_n868), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n883), .B1(new_n869), .B2(new_n877), .ZN(new_n887));
  OAI21_X1  g0687(.A(G330), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n451), .A2(G330), .A3(new_n847), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n805), .A2(new_n807), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n807), .B1(new_n687), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n882), .A2(new_n875), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n630), .B2(new_n849), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n305), .A2(new_n661), .ZN(new_n896));
  INV_X1    g0696(.A(new_n868), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT39), .B1(new_n897), .B2(new_n880), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n861), .A2(new_n899), .A3(new_n868), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n896), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n890), .B(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n688), .A2(new_n451), .A3(new_n698), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n633), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n904), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n260), .B2(new_n654), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n543), .B1(new_n587), .B2(KEYINPUT35), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n909), .B(new_n230), .C1(KEYINPUT35), .C2(new_n587), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT36), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n232), .A2(G77), .A3(new_n404), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT102), .Z(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n203), .B2(new_n201), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G1), .A3(new_n653), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n908), .A2(new_n911), .A3(new_n915), .ZN(G367));
  OAI21_X1  g0716(.A(new_n693), .B1(new_n593), .B2(new_n661), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n667), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n637), .A2(new_n660), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n611), .B1(new_n922), .B2(new_n502), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n661), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n918), .A2(KEYINPUT42), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n530), .A2(new_n660), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n634), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n534), .B2(new_n927), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n926), .A2(KEYINPUT43), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n926), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n678), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n921), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT104), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n939), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n931), .A2(new_n942), .A3(new_n935), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n681), .B(KEYINPUT41), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n671), .B2(new_n921), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n670), .A2(new_n922), .A3(new_n946), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n667), .A2(new_n669), .A3(new_n921), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT45), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n937), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT45), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n951), .B(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n955), .A2(new_n678), .A3(new_n949), .A4(new_n948), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n733), .A2(new_n664), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n957), .A2(new_n678), .A3(new_n666), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n666), .B1(new_n957), .B2(new_n678), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n953), .A2(new_n956), .A3(new_n731), .A4(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n945), .B1(new_n961), .B2(new_n731), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n736), .A2(G1), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n941), .B(new_n943), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n254), .B1(new_n815), .B2(new_n402), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G143), .B2(new_n749), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n202), .A2(new_n769), .B1(new_n766), .B2(new_n211), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n744), .B2(new_n201), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n775), .A2(G68), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n826), .B2(new_n753), .C1(new_n316), .C2(new_n745), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT46), .B1(new_n783), .B2(G116), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n785), .A2(new_n816), .B1(new_n213), .B2(new_n758), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT107), .B(G317), .Z(new_n974));
  OAI221_X1 g0774(.A(new_n349), .B1(new_n753), .B2(new_n974), .C1(new_n815), .C2(new_n756), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(G303), .C2(new_n746), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n783), .A2(KEYINPUT46), .A3(G116), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT106), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n744), .A2(G283), .ZN(new_n979));
  INV_X1    g0779(.A(new_n766), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(G97), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n976), .A2(new_n978), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n971), .B1(new_n972), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n739), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n929), .A2(new_n792), .ZN(new_n986));
  INV_X1    g0786(.A(new_n796), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n793), .B1(new_n208), .B2(new_n386), .C1(new_n240), .C2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n985), .A2(new_n840), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n964), .A2(new_n989), .ZN(G387));
  NAND2_X1  g0790(.A1(new_n960), .A2(new_n731), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n730), .B1(new_n958), .B2(new_n959), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n681), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n960), .A2(new_n963), .ZN(new_n994));
  INV_X1    g0794(.A(new_n815), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n995), .A2(G311), .B1(G322), .B2(new_n749), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n767), .B2(new_n743), .C1(new_n745), .C2(new_n974), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT48), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n775), .A2(G283), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n783), .A2(G294), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT49), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1001), .A2(new_n1002), .B1(new_n543), .B2(new_n766), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1001), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n349), .B1(new_n1004), .B2(KEYINPUT49), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(G326), .C2(new_n754), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n781), .A2(new_n325), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n289), .A2(new_n745), .B1(new_n743), .B2(new_n203), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(G150), .C2(new_n754), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n775), .A2(new_n512), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n749), .A2(G159), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1009), .A2(new_n981), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n349), .B(new_n1012), .C1(G77), .C2(new_n783), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n739), .B1(new_n1006), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n664), .A2(new_n792), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n796), .B1(new_n237), .B2(new_n794), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n254), .A2(new_n684), .A3(new_n208), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n684), .C1(G68), .C2(G77), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n385), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(new_n1017), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n208), .A2(G107), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n793), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1014), .A2(new_n840), .A3(new_n1015), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n993), .A2(new_n994), .A3(new_n1024), .ZN(G393));
  AOI21_X1  g0825(.A(new_n737), .B1(new_n922), .B2(new_n792), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n995), .A2(new_n201), .B1(G143), .B2(new_n754), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n203), .B2(new_n769), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n743), .A2(new_n385), .B1(new_n220), .B2(new_n766), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n758), .A2(new_n211), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n745), .A2(new_n402), .B1(new_n316), .B2(new_n785), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT51), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n254), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n746), .A2(G311), .B1(G317), .B2(new_n749), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n254), .B(new_n1037), .C1(G294), .C2(new_n744), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n758), .A2(new_n543), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1039), .B(new_n777), .C1(G322), .C2(new_n754), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(new_n767), .C2(new_n815), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n769), .A2(new_n765), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1035), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n739), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n793), .B1(new_n223), .B2(new_n208), .C1(new_n244), .C2(new_n987), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1026), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n953), .A2(new_n956), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n963), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n682), .B1(new_n1047), .B2(new_n991), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1049), .B1(new_n961), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(G390));
  AOI211_X1 g0852(.A(new_n871), .B(new_n310), .C1(new_n287), .C2(new_n303), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n874), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT108), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT108), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n873), .A2(new_n1056), .A3(new_n874), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n847), .A2(G330), .A3(new_n891), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n697), .A2(new_n661), .A3(new_n806), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1061), .A2(new_n808), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n728), .A2(new_n875), .A3(G330), .A4(new_n891), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n728), .A2(G330), .A3(new_n891), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n875), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT111), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n875), .A2(new_n847), .A3(G330), .A4(new_n891), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT109), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(KEYINPUT109), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT111), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1065), .A2(new_n1072), .A3(new_n1066), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1064), .B1(new_n1074), .B2(new_n893), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n633), .A2(new_n905), .A3(new_n889), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT112), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT112), .ZN(new_n1078));
  AND4_X1   g0878(.A1(new_n449), .A2(new_n905), .A3(new_n632), .A4(new_n889), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1065), .A2(new_n1072), .A3(new_n1066), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1072), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT109), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1069), .B(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n892), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1078), .B(new_n1079), .C1(new_n1085), .C2(new_n1064), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1077), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT113), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n896), .B1(new_n892), .B2(new_n1066), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n898), .A2(new_n900), .A3(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n869), .B(new_n896), .C1(new_n1062), .C2(new_n1058), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1063), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT110), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1084), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT110), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1091), .A2(new_n1098), .A3(new_n1063), .A4(new_n1092), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1094), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1077), .A2(new_n1086), .A3(KEYINPUT113), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1089), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1100), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1087), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n681), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n898), .A2(new_n790), .A3(new_n900), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n349), .B1(new_n980), .B2(new_n201), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G159), .A2(new_n775), .B1(new_n754), .B2(G125), .ZN(new_n1108));
  INV_X1    g0908(.A(G132), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1107), .B(new_n1108), .C1(new_n1109), .C2(new_n745), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n769), .A2(new_n316), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1112), .B1(new_n826), .B2(new_n815), .C1(new_n743), .C2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1110), .B(new_n1114), .C1(G128), .C2(new_n749), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n980), .A2(G68), .B1(G294), .B2(new_n754), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n995), .A2(G107), .B1(new_n1116), .B2(KEYINPUT114), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1117), .B(new_n349), .C1(new_n765), .C2(new_n785), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1116), .A2(KEYINPUT114), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n784), .B1(new_n745), .B2(new_n543), .C1(new_n223), .C2(new_n743), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1118), .A2(new_n1031), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n739), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n325), .A2(new_n842), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1106), .A2(new_n840), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1100), .B2(new_n1048), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(KEYINPUT115), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT115), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1105), .B1(new_n1127), .B2(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(new_n1087), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1079), .B1(new_n1131), .B2(new_n1100), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n331), .A2(new_n658), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT117), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n623), .B2(new_n449), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n449), .ZN(new_n1136));
  AOI211_X1 g0936(.A(KEYINPUT117), .B(new_n1136), .C1(new_n621), .C2(new_n622), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1133), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n619), .A2(new_n620), .A3(new_n618), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT91), .B1(new_n370), .B2(new_n374), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n449), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT117), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n623), .A2(new_n1134), .A3(new_n449), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1133), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1146));
  AND3_X1   g0946(.A1(new_n1138), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1138), .B2(new_n1145), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n888), .A2(new_n1149), .A3(KEYINPUT118), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n734), .B1(new_n879), .B2(new_n884), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1146), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1135), .A2(new_n1137), .A3(new_n1133), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1144), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1138), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(KEYINPUT118), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1150), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n903), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT119), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1150), .A2(new_n1158), .A3(new_n902), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1150), .A2(new_n902), .A3(new_n1158), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n902), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(KEYINPUT119), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1132), .A2(new_n1163), .A3(new_n1166), .A4(KEYINPUT57), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1076), .B1(new_n1103), .B2(new_n1087), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n1171), .A3(new_n681), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n963), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1149), .A2(new_n790), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n289), .B1(G33), .B2(G41), .C1(new_n265), .C2(new_n254), .ZN(new_n1176));
  INV_X1    g0976(.A(G128), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n745), .A2(new_n1177), .B1(new_n316), .B2(new_n758), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n760), .A2(G132), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n769), .B2(new_n1113), .C1(new_n743), .C2(new_n826), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G125), .C2(new_n749), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT59), .Z(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n402), .B2(new_n766), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT116), .Z(new_n1185));
  OAI21_X1  g0985(.A(new_n1176), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n254), .B(new_n265), .C1(new_n749), .C2(G116), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n223), .B2(new_n781), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n745), .A2(new_n213), .B1(new_n211), .B2(new_n769), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n512), .C2(new_n744), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n766), .A2(new_n202), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G68), .B2(new_n775), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n765), .C2(new_n753), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT58), .Z(new_n1194));
  OAI21_X1  g0994(.A(new_n739), .B1(new_n1186), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n842), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(new_n201), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1175), .A2(new_n840), .A3(new_n1195), .A4(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1172), .A2(new_n1174), .A3(new_n1198), .ZN(G375));
  AOI21_X1  g0999(.A(new_n791), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n745), .A2(new_n765), .B1(new_n211), .B2(new_n766), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G107), .B2(new_n744), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n223), .B2(new_n769), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n254), .B1(new_n995), .B2(G116), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n1010), .C1(new_n756), .C2(new_n785), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G303), .C2(new_n754), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT120), .Z(new_n1207));
  OAI22_X1  g1007(.A1(new_n815), .A2(new_n1113), .B1(new_n1177), .B2(new_n753), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n785), .A2(new_n1109), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1191), .B(new_n1208), .C1(KEYINPUT121), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n783), .A2(G159), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n746), .A2(G137), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n743), .A2(new_n316), .B1(new_n289), .B2(new_n758), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n254), .B1(new_n1209), .B2(KEYINPUT121), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n740), .B1(new_n1207), .B2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1196), .A2(G68), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1200), .A2(new_n1217), .A3(new_n737), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1075), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(new_n963), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1089), .A2(new_n1101), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1223), .B2(new_n945), .ZN(G381));
  INV_X1    g1024(.A(G375), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1105), .A2(new_n1126), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G381), .A2(G384), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n964), .A2(new_n989), .A3(new_n1051), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1229), .A2(G396), .A3(G393), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(G407));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1227), .B2(new_n659), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(G407), .ZN(G409));
  AOI21_X1  g1034(.A(new_n1051), .B1(new_n964), .B2(new_n989), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n1229), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n964), .A2(new_n989), .A3(new_n1051), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT125), .B1(new_n1239), .B2(new_n1235), .ZN(new_n1240));
  XOR2_X1   g1040(.A(G393), .B(G396), .Z(new_n1241));
  AND3_X1   g1041(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(G384), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1077), .A2(new_n1086), .A3(KEYINPUT60), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1246), .A2(KEYINPUT122), .A3(new_n1222), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT122), .B1(new_n1246), .B2(new_n1222), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1075), .A2(KEYINPUT60), .A3(new_n1076), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n681), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1221), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1246), .A2(new_n1222), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT122), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1246), .A2(KEYINPUT122), .A3(new_n1222), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n681), .A3(new_n1249), .A4(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(G384), .A3(new_n1221), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1253), .A2(KEYINPUT123), .A3(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1232), .A2(G343), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1260), .A2(G2897), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1253), .A2(new_n1259), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT123), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AOI211_X1 g1066(.A(KEYINPUT123), .B(KEYINPUT124), .C1(new_n1253), .C2(new_n1259), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1262), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1172), .A2(G378), .A3(new_n1174), .A4(new_n1198), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1163), .A2(new_n1166), .A3(new_n963), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1132), .A2(new_n1173), .A3(new_n944), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n1198), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1226), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1261), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1251), .A2(new_n1245), .A3(new_n1252), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1258), .B2(new_n1221), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT124), .B1(new_n1279), .B2(KEYINPUT123), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1260), .A2(G2897), .A3(new_n1261), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1264), .A2(new_n1265), .A3(new_n1263), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1268), .A2(new_n1276), .A3(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1274), .A2(new_n1279), .A3(new_n1275), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT62), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1274), .A2(new_n1288), .A3(new_n1279), .A4(new_n1275), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1244), .B1(new_n1284), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1285), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1268), .A2(new_n1276), .A3(new_n1283), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(KEYINPUT63), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1295), .B(new_n1287), .C1(new_n1296), .C2(new_n1285), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1291), .B1(new_n1294), .B2(new_n1297), .ZN(G405));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1226), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1269), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1264), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1279), .A2(KEYINPUT126), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1264), .A2(new_n1302), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(new_n1300), .A3(new_n1269), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1299), .B1(new_n1244), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1244), .A2(new_n1307), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1295), .A2(KEYINPUT127), .A3(new_n1303), .A4(new_n1306), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .ZN(G402));
endmodule


